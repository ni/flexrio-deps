`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTKvhqUA0VVZBaUbikje95EFLyuyWjuFQFq6LLrWmYUac
5oYcKqzZVgiga5GEpz7rQhNqokFxUzmuaIk7s6pHMc3Zr3fd604ieF40HaWD1Cwq
zJtIY8fP482h7yUl+daE7QM32IlbZY/ym913lk4/ZAtWYgl5I2oTtaGuVZ5s7onw
4Gab01URF7QFzC5AY5/z2I+RDBPIGjjMoGKZwWqZzWbxalxscFpedugfABwJTuwx
OtIxGvJfKzOWxD89iSNzfYgV99EaqHhXoV0LNzTeEGdrGOOVQNzI+979P2leoO9p
Y3xd88uriyuo+849WAlHk6oU0psg9/7nbwQssWyBJzJl9Rp3KRk0ct+JFl6T29ad
u3flZEl3NtU/H1k8EVaAdBjL8g/xS/QkopDuxtBy7oDK3AGQbHoA+nBNagi+NW8Q
8ieLCRE32+ms2nGu0AvbBgjMg0PBnhS0RKtQRS/g09y6sD/zvHKS3x3O+CaR++M9
gbLqW8031hTVvoj5Qc4n0Wb6HeJnegSzu0Hw/gYfZry+QLJoXPHvpWXIMyNx6TOC
jR17mmUmhd1ZgKVL9J7uYwRi6p6PEk+qFh6cBwGIL8PwSzsVjMRfhKM1+oaDPaHw
SPtA89ZbXEBsfpYuqKVxVug99kpDk5Fi4fZbU8ayCfx7ZnB9Ampt2ASzLorn1vsQ
lZTCl73mTHP6uHTno3A1SW31CZ7PNp/6zFZwZQiFjUG9YXNe3xvNt0z1/ahtMk4p
TMWUWaB64ip8xh8iFzaF49ufXjglvLAauUVx4m3sqkGRlkT+vlDtqtOutZOMt3+P
tUm2gesFDSkRsXlNJqhCXqam4Ue7Dy1ubQMN/00LXvAm9wM+T8aM36gOr4w50cZ4
lDSePHkAXEHwl5imeZIsI/6YyU1yKn843FVPKCegIoVjE87fJU2juuotvHZwF0Cn
k5J89ixbo2eV126edLak0mANGa+gBRLjbIOqz+F7s5OvhD6dC3GAZ6Dq2cdMbXdB
xICGaAaX2qWCljRimV+yj+hajzGZa64v/fdO+ti02FQfTOqWFQx5s8iPQaD2bR0+
BIpx8zvESFDB6qg0PXMFR0zFcJSAOPitB11vYlqx+vjTHn03+G3lUCwbX56KQL3/
Qp06gS8cO4sNwdlLW9/0NqzPQHYuCqvWpCNoDqhJ2BkuriC7MlvntYaWPRqMOVXr
QMyri752JA41Co9LtM3PtOnxhdIrHNbwu9VEPLhW0X5RM3Lxs7MmQ19Ehg+9EvmM
40yXozU548CUX5Qw6eKcsOa32j9JVZ82MI2hn+CEzel+Xvf26k7qf1dpzIKfp2Bj
0SwvqG8xUQmqZ59MuqHyDdcxYRLp2KfAQbR/upAEd5lix0IknsRgcpVZfNF8gmvD
gvU0fpLCR5kXnr2PEoK1mW+jcCQkPVrxX5Qv/c88UG0IaKONM7XF5DgXCsJnx0e+
RHJoUFGc7CnGso2DFwBdjuo5AFTSUoyClHqhSpWW281VZUwg7o003sZ0DyuutQZ+
AdGTBmu0ID7YMPxooQT/KSZUvAeqs3dF6+5E4rWV1IxnwDEj0hbrXH6/vH65EQAU
1I4mW5Yn/fWoG5zLMjhA6WBb5sYc2EqC7u820EcI8/GED9Kxz9Gx+GubwHPzhaUy
f23VFuG+mERmXgWNw3AM9r5N7y38ff5fANx9BOnk8tOJQAvGPMI5TslyLD8amLYf
mqdmSh45mBYbAL7PRAtKxQt9wuyiSiP3SxD9oDc0aTIJ6mLnsE7zQ6+phyNDbwjE
3tmwbg5q2oEWXsASpcNi6Mr8w/mDgaCo8g6ju+0BxEPc+l0gEVhQqbR2UHKMrpQk
eOva9EM+2DF/70P+/Xkl84JFtYSAsoiSOekzvVbS5/upCc4QIGIdvupman/re4c/
Z3PWng34hG4yVQr+1YEHEZSLWifRoednWCnOuv9EGITcR7jj4HYIAwnVr1hOUNNn
kw5D/YPhEDrrQPpAAXys/Ek58/BQATJWVspw8WvzH6goRQVVzeBarzgHV2fjPWAQ
6GuzbSw5D5N8aSyE3q4krG64xei7Ubzju2ioBMwRUT8rJ8AEazwdkQyO21aGWbOU
WZqU3AN3qDSGOL9oSodRqwvIfdMXGtyKo/qsz1U2G6QYs9hiwzvQX2nIBZRZDAyW
n6V6ef9b+0Y+9sSzj9rGi9zJJ/v5Aan5gAn8jyO8vYdDULs4E+WbdbqMB2y0F+a+
JhVtfxhf43PlO3UrDeBdgKzLo4aeE6WLpbUkSJs/78FT6/VCzjsyeKkPt1JvlP+6
GGjCh+OMlBsiwq0rc+M9YaTBAIAnksKDuVV7GtPoQM7AExknldV5Sx6ikG6aMQie
8WaQ+DUiMtSa03M90tc+AWq0XbXOhmg7r5RIXg2uu+ogzRPLLKVR3TqXHF/b5IPu
3FlL5Yo5IyftJB3KCGP6PVLptRRSjkqOMjC9l+6W59GAY0Xn1357N8CKnWlodcKt
/EaJtLw01uNbaZnSxaYdRXKcLhSPDemyo+zLAkE949gCA6ZKtv9b/Xf/9X7exSqk
VENAijC/vPb//nI7vRphZOuPO7ZgurzLgaFRl8QdMbJLKAARE8HzGwVjliY4oayw
+FeFeGhb7otU+1utRJsIMNuZ67cfFTxIgA0sr4d4IKc6OmNFgrFJ2jyNfOP9wPeb
k3f7wCMXWb8J3z5lyjXj6fKu4BHaCMzRvET8f4DCOlPXu/eOh7SO4mLPv0rvgLGM
adJTPcQXNV8VGAYZ9SHEYC69fJvsaSZJKCWTs/6s9uUzoZCkInTF3iTHMyH+GDji
C+Jyxb12rrajbdH7861yC+D0EbHU9ofUjIOkdTiV2AtduOraC/gfI4lOr7GLPfOQ
ykXGndLeLfLl2PMuPZGF8whRVFpLcfBHAhRDUlNIflzG5DubirGclXOn7p+CBZom
OcNZ2xq2y7fmARymmwBIWcEDvuIaBzDIVwi8QNr3kmFk8xBmUZMykVQyY8phkp2m
rmbBRtrcMNDKSYBCG6ZXfjudis0f0F2kHWV07wQyALrfeIeh1uNA+SkUs8GGZfz5
Vf+p74o3g+4WZdLTyo1ohuuGHjg6PvEn1a5GLUR1HsTxy+xA1Lr6URsg7ATnInYd
3Jncg6P6ZKUtwss8p8+qoFlrnjK3A5qIwNUIO2Y6PE9TXXjWUf8D/UALFQAL/G3C
Dbgfxo1xU+4J5r0UOMq3L7gDFo29sjH2w84CxtYW88EkfOvk7sqp0dBXazOel6vS
1SUj5zjpBv3D6TlLc9g2HZutnH/iXl46QGeXCwGdqDrDN9CJSCmQfsUPN/YO0SpE
h53v/1if6dUkMWTvHmQwEEAlmaVj5pN3Kkww2hcOsKz145jegUwSek8+3ym4WaZC
K8uYqRmwlTzA9i3EjdoF5Tt2nlq5SMQ+jH6dxID45mtTa2eFst7XNA5s/Q4k1opD
6/AiHY/0cP5B2FUjDVP3Cpk3dmbxV1Gxqg7/fXV+64s0Xdy3OWJsn8K8FaUM8xZZ
z6Qja+8Fu5wD8koL0oWzWk+QNQzgolCICEvImUdUFVAxftJKLh6hQMM1C8dEUonT
L1obt51tbJo6WlfFfp7U1XWjKOpdDe+MUDXaKdXZpu08OQF7tjvy6ip3LKCtM0hN
DvIO35uwTCgNzZm57/M9Y0bFD7B5ZOB96pI/PpbMexVxQ+bec3z4mmEnR6hf2ImR
SI8kAS5i/Obs0eP8LywWzwwUipcSimxV9hvosRsXUCXpjfeeAB1390NBwfqM7XAg
NJLgG1chYmE5/oOcUvQqqgYtMcL8mlLje8FfZIpK9dAeKIHpX/F5w0LsoUy92ZGl
pne8r2zkrb9M0/2Of+ieAj0GYrjcwvbZLMfvA1mEn/cI2NNsujc5KPYPjRzVXDPW
x778P1eWoY2XaSY7fWtKaBF6r6Bd5QBws5Q+MDsPRl9mvHeRoZ74HMauMXSI8+Uo
o7euM4wrhQYe0msOKO25s6E+j1VapCtQGPXQUccYxknmGpZ9DdkfYSa/njmVZnSD
QXroIgEB6xhLBlppOYR0YndmmxpbeAj/orlTOlCI8iP7j4KdcRI0Qh+E6wON9uFe
75jeqYWcUO37l2MhW/amDo6qfQIYYJl8iPqkJbYNpURk6LmQZ46TdlD0sok7igQG
T5F0s/PgaPNnQyP5TpGm/RsLZqKFkhB+D6RZs5b8bUnr9UrFAZ8P+rLfEBgX8Raj
l+YAMCIftHqBp5B86aYeRzL2aee8XC6yXF4VgXEkHc8cYuADe4T5C7JEA9TMi50b
YGNpFZCmofAfMPjAEgDb+Lb+gAVSODu43imz0PD2je7yPUFMAiMlwDibjd6SNOpp
C8e0GyZia6b6dRFvPrT8xpC2DJ79xJr+TYtwUSabCV+eTstn2cGTT8TLhkmI9I+T
iwba1bp81U8lnXhCJGbNbn+bSiwVqsJkVkIBbTs6r/Xnj2QVU/KRPZblJGXodcYg
WLrl2hzQ5911k8PjUYYQJDlPrkRapIIr8kEanFG3DOqU97UQI8le1SH57eBaVtdD
cw0Agdmu9FoqEKt9LMpl3bnEGMmFBBtobOoJjiCCjYH3YUrxm3dRqT+GXdpCoe8J
5bybmU/UR+2CgJ1Tmvclk4YSTZQ4062NbJIjPKL10iPFWCUixDV/ZoVw+xoqNYrq
Hf781laGKjsiIzs4SMi0KZvvUOpZ+9EihPWpTLy2vRci2Kg4WMddgTF36JJdIrSm
NmIP1e7GmetBf5p/37t5aG4bgLIKbhCyqoJFIEbTAXmwCXlo57YAe68UwAiHFkA/
zXqpf5fmezj7u/A5cwnIkOweXUb2wW9nRrml+pumor3NaWWiTK0iFFUwBR4jFaT6
XD2bPEIyAtviPE7n/zY5uiC0jRLvnv6yas+Cq1BUiySknJpA6Px39ztaX3Xz5IhC
/bKhcCAcrxgjj/S/p/sMWMHLXUlsjXHqxk8asQAhuqW3CYg5CdYXOWwVNbxz0A8g
Wng/df0053DOo4TDSzUFx0phH1JPMZLblZ899MWaFNU2J1vI5IlLiBvrhcUHYlFF
lGzTT+cB7iluP9SVXgSVj+YbuArw5QOOypE9gcdJ9uUUxlI+CmkKDtfyMpZb9dd1
1N7dYb1CSfmVkYArSBP9j3rL/UPn5SDjHmODubA1ezgtKj2VjePJq7KbuoizEJjK
i8V39L5UKFBlavS4yOIRQJZ17GrjnRSu1nnc5O9UHZuVx1JdgHo5h9dLeYBugAkd
yMZ6k9cGcocMA7M+ABY/SSbXFOxCN9FDpZ1sfanAvNE9os5+Mt5SRfP0AJ0j9SJT
5JECpJLn5PdOOwePH+r6712tmQR+7Bw34o9BHb64x1YT9JCad1bzSU8v+JVkol99
5TElCjZL2RyvFHu8ZrgrVJcs5jfRwLCOjaRAZ3sSnkIJRpPmdZI6/JVXGkxfcLId
mUyYY+ZIsMozIn6FD33xBS11ATwC17bfs1w9jpmrQMvlTT5bFGnzB2uFkEcSxx88
zkXXyaMA5Mjnivv6lATY/x83T+XmCqysoqkj/z0ePr1bVkIH0GpGOnghQEk9Px4Q
ZuWMDxWznLjSPedPSXweGrpz9vgOUGvaW02MrKSXWS41knoOnPAQJHrDh7Y2Iqdw
zs7UbDsdEjSRbGA3HStqF4De8BE3rh3GRQZcQ6xAwywussVdr7FRYL6Od+GBDklh
zTzUeZthdjD/VzkAemasqinsRI1FsfaP2X+BmZ4+En+nkrREL5X50o6XRK/dxowl
UKpMPnxo91CtfS5FdMmSdztMOEOQ/KWy/3cz1hAfZBcPr7/H+T7rfwg+LioLG/TJ
dBzmMEbhHI4aXjbsDCFKV9C3DLxJ0YJu5wB3W9yCOq+Q20Kh72MnvVuhc/hnIkCY
73BvU3EbtKWH45BGO1IIB60ZoHWW6NGCPPhuZ+x2v/ub/BggF+k1vVdypVx9hjBT
MM6ku6so/qvm+PIEogw9KlWuZHcQ1h5niqDU2zg1ZfkNRS8gKEwtH0LrQInHe1Uj
3QHWhhbL0e3qq31QdH1e1U4T9jwnQPmMEsVxswAz8S00Cdge7jKj8bkxNDr3kZSi
CCPQ2fsdE1EjsGqJWG9NIPhQOeD1+iovlWjn9IFNJgx+IxsscO8zh6G7fbrN8/OI
Be6tWFZgWwpuXyT2Vcnaq4/yEjWRWEezDBUvqeyuNzhRTr8S5sbZArRScdvThEY5
wRJdNK8hm92ol35xIES4tH7t5TuQ4AjKxRR2eiyFegN0+KhBZOfEu3BEJoSIMr7w
g+wBGcuaHDd4d7bp+PAvg53+Xq3EjtsIhWtEh0TeEUXvAjwsOC+/cQOtgsr29UJ1
FrfQzzxg6pIhFujuRJB1iVk8rOlT+aIMNLkAMCZYcc0YAC+tCLhE8Q7UzMWHZs/e
8B56duJjsUrESNBRVJjMA0xmTFJL+1lQ5xNemR8cvP0LtYdh8kveU/ebQp39Q2UN
p3qHRCIRdqiD6neUTS3NMuR/HPv41EvfMhO9orc0xgcFimebPi3WTeBm1xxApmNW
TVYvyU0o1icsRV4wH0ngYtAt88LRQhui/slRsLFcd+bL2vQQAN2Ut6dM3/49sPBN
cCKfb1YnmZk7flNe6n39ELF6f5ljQm0m/hf5JtxXO/tZwfeDu8pQr69RcsOswuuz
1n10sx5Ym6kv2GbYAcUBz8zkEi5bWgNYEY6RaMvtrjzSpea1lR68J4bgNH6fyg0M
drLVblPycXM0mVrqh9JX8Yn7ug5vKhkAvrU35nib54mhUB09seHNdj6zK6P5MAZM
ZmyGhBs9WwLSL3msf8ArZmdAxN/uuttRmSC3o9PBWIXEKCLJh71tY8yhV/VE2urt
q2cx2M+HL9cgEbrwvBe5jA6g6hjm72rfGCY/yWxum6xFg6DAeNYFJV/oZJ2Uuf9n
JYUFaQROydHwww8sPyBweF2YcL9pX4pCDtbzrj1LSvC4F69nHg6yTOWg8EAuVCi4
Tr1dLwd9+uU5t5ry9kG1XYOn+7ErhEid+ss3vsvVsn4lhPEPcQeL4LSuffHVqrOm
RBQYiA8GJFNgVi+jVkgmQ2WQolZgtH8oo6sjUSbJTcU4EV1XpFn0DSfha6Qp4Q9V
HwQVOMwNiqokTgRHN9CyCHXkjV1jdqLaN2zF94g3YZAcCK+Nd7EzJkwtl6EVfaOd
mwzleUTXAg9PiGSRii8tst/7Hl7l586osNleZcC776J985D/KWmB3U30rzpz/J/L
iAcaKwedsl1bO5w6ieLgNf7ezhIQg3/ACrFYfdAaT8r8n9RdrudHM+hoqA5z/ANV
vhrR74vF9jkyWBBK4W6RSl7l0WcKkgrve2mekJPRRH1AX0l2VoCTc1vnsphOQaLM
AOsI2zi1R4cmG/u0DD0bjr6r/HchZYNfby9Ln98kylKkrlwLycZf6nOQbEQyCezM
nfCcNT4F5WshefiCKinPNnuR3F6x1pVc4b3Cs8CKVmitkJVVpszMcAPyYP+bLkBq
z2msuL7tFlry5XQCXHzr5NwswY/iTD87hQyQ6bA7vWOR5PgmPpZN1sdQWRWdf50u
rXT8fv671RM1u93vwl296BN5mpnCG8kFfore33Hdlom44UL6M/YYZknw9iATzVQU
G6NBem9wcqxGjW+VCVMXx9rjBsBLvyXum/cn9luKsO29MLdmEoU6OlOM2QLlIUUC
5YY9wY8McbW6Qs+s/kNyU9EWpv2uFCUKoj5v6yXGZUxvcRLxRuVH+G5H1GOSIgXx
EyGXwvDGSKQH1Q4I98alXSfNPwBxLl/+SGORyqoD30JZMd90ULjXsVF8Y/EehTFW
RfooWnbC377Jx22SSbuH8/emewNz+9Z79siU2KDGm77aNRbKE+AKEFc4MEFMjgJn
PD0zed9Pw0KA8qFOsQO6nWtQiTIF60/Gw+X91JdD52eDXsX1fEln8ZI0ZXfmGgL7
29+cwrWXI2igSWdjhEuPMD/PWnGlNv1YOC72mRybhFHCzxPFEof9Wr7obcWGjiyc
3eY/OGkmpgyQiPOBGDo+doeE1Vi/+gUESy2r5axohyxGaAiaqvjEnYlp65h7tD2S
XdbP3tk+z/QeBs+HLx5UqCeDfe92F36LTI2xQYFWkMkMNy2p5c/xWZ+Hs67mKaGz
ldIKMJ6NjWT7QGReuzP3bNcL0HF433JD6Ehin6R+ruZIPfsy9bKPvmvPwRNSmf7a
wp+1PEXdRVcumAdQL9Sw3gxs2PlyVxKuzzmsvH774dt6RBNgHB0qvw03hfjzjRgd
t7GBWQx7Rz1gnFXZEb49Dp0W7Xy2RcxQSOinE/vyzSXIm/UlAEKwYDB+LjLrqQsR
X76H4CQJ+1Jp8RDZZsnJGCqlmxOm0tVXQsQUzMebmFPL9T8dOKg/M/Q3aamxAELy
pBwaqeeg1Tir0TDZUqy7KAEd7hgrJOgGJJlpuKocaAl7kdqDClrIJDAExWr6qUuO
oCq+BCLwwwTT0fn/bXx7CkUp6JVku640zv7wzQGxtf8R2l0oUP9KniJEq7ELcTVQ
n86PegVsZxr1LHyPFs8LZ5Nk3hSMgMsfP95tWEVZgg5Gs43vsjmM3lXcW3ikbMfr
1M+AiMSnUqJuT6QRDB05IUDkDYujX4Fp8ixvbjQ65/I7MCx57lq0HlkSah3dEakr
SFJsW3H4CI70kQvxiGUg17gPnEYh0gBCd/OVLG2cioZHuniilEGCa6gqCmNpt3ns
YiPSy8gBxM+zR9ha9tUF/kpMacAn4Fg0g2jqQrsJYlnOsA0SluByu2noogB/jqiV
qumUgpMILQQX3ySYpe2/y7hjiShfGQoJTsR1oTHw36IICbe2msihr+NYbj/fqdAM
eBn5zRNVcDnRPAbsjRpMe8d7KQipVpWk2H95xeEvGLGkVojrXld/5iprRGkRgndN
E2QkaEbDRjaRAsLotPpaSIpFI4yFhgLZ8sZCdPixbMQ9yBSkwJSOEKF8RyC4a5lD
EzxhPL9JzJS1+Zibs7ZaOfEN9PB6PmYTrGPy+QZ+hGuQ0ZDOcKwUMNUIQNDe9jgf
vRd1xOxysJUTB7YPLkzvBDGYiOz0s/WdGxmesm/dJoypAnul0grKiPHMAFAvvtZY
JXSkNVLTSIuB8Df5D8dLdAU5GgmW7ahbAkVCPWehnlE0PiJFlHthjaidNqR1yBOL
8jtOxF/lioBE5HPT9TSIy9a/tMme4sTzWekvGCL29zEDwrH4yaIyf8AbswHbomM1
nEnS3+1Kp/15LE3+wGBXqWgqG47smB5sJ9iNpliCbGDUZigVyS6jslhTKBCkkqX1
+EcOMI3CE20VwR/G8f44PhCQvlR6F37uv7BoIS/atIQo7SqvuIPrrCcwtQampEjo
Ti0vPNtOzc3uL9JrEOK1jy9N429w1+1Y5zFAEIQVslh8cSV7/6Knrr9HcTSDoalk
3XtVAJuGrex8HPAD1i+0zuAhiw4HgAgB6VdEAhVQNLH34hIzFekaWr8eLiqZ4GAx
3pSKStrKIBtsYwCE04qvWK/CQFOoH0BQaG93cS7GUgi3JsdKXavBhyoRXp0xZUeI
WnNzbtKEpIeS7dHhYOcIg/fzsZmvKWohUy8pFbSQDskDtHE7ApqghuwV1MQxEoqm
NFlnL7xtj9zuAx7QXCndW371VzGN8kmR+LKGMxBKtVnYCPOoIo97oMsHKIOm6M3P
h5M1f3bKK8CU6+G8ddsA4bino1mOlSvb6s2lRciFttt/CSdYRRq+7RgKff5SrqTF
+cS3xWaWgorH2ZJ7Y13uSuYhkaHp4wf3C/x4nTftTQ4a6yxXZgty6kUhixplvlI6
f4Hg42Aku7u91GVkvkzQZejYpdZmurnQ69SCkHEqAr3uKXlv/bz/9ypaBT5rz9YK
LAuRCCX8yxXSyfAZH8YUjtnaBWY/3S76G5/+4OulOxaccWb9o6bSQaLQzNTeqZFq
V75AmfCY0aE7mAbOfpDyM2eztZbNZ0x3c4hEdj0NETDmDnMs+nD4t1JqYNi3D+dV
pcwCrYlChq90QrMSC4vK50//ykysQe1AuRyu+ar4kaQHBOnCzE8yazZmxHHPcmDS
x/PqL6jmC6GYRraONGdQ8OIhVHFcfyrL4k8L9E6sytjA/ebvtsP8bnE/J8aaF5RF
mixzKniMCPhRp+v8C7YRk3hsmBGb2cJhft2jX23cqN/0aeWeLrgrbEICLDh8pNIc
Za88IyOoL275sUWQOvOwv2jyKedIf8oEo/RDAE3iovi6ihucw3/fH++cP0duzXR2
W5ub1HYW2Dl+dyv94/m6HlG6nuia5BGffg+RAGDvjXf5pbgxev8qCeKru6AZNYlk
bT0puiSfP8cz93URm8DrgS2hjfM3hJqVXWMd4Qe/QDdWjWZ1EBdjKU9THp+T3yoa
6Knm3E3kC3Xp0kKqm2PXXkrs/hgxpW6eqNx0GJdGIYlhoruO0J6DQDpprFUh0yOx
O9xl7mUX8mVGdeJKdRlL95wwjgZcGC9UCEEGRzFZuUPj0GaSKn6DSpwtfxmUk/5S
sJHN+gZxKDRrVA1bsvDkTXvFlNWfG/0Gnu8pVt5h5T7FHw5lfiiNeT9sHTNA1mAo
DbS1h+BauAoZXuV5bnsk3iH/0CgW+Ks7zWgUiOi604AZn3N7xQJTL3CeGK7AzyDn
dQ3Pi3LO/W/75O3b+a2cUM3wNDsuPWEoAdjhpkjJyOz1nmrxCxB/P05qcrq9gSbE
JVzUyCE7p5O2TOKYL7XGZzx+xLh8ybj32i6oCEmUqxQGYHpVatjGSOzX18zoWud7
7lRTJgOzjdZmEaXQpEIq6X7Q/Ab9QVWDLS6TzE/4RBb+KWfTRKQiBWE9Dn5gEcq/
+oO/kLZVOSRHYoGRbbCB4is7j7qh/LFiqGoeMny8FiO73fO53YlQ/H4DP41VmRqY
95/dlP7tQLLhJt6SvRSOneK6UvjMT9XwMCQoxAEy1mLdFyrHTQrfQ8JqIYFGh5gj
uy0VtrSxOrnNLlaWbuW3G1D1UY5cq0MRW9tp4H+MwpbIULfN4V1+xcFFzpumvb2r
udacKgPh0mDceYvdxC7vjhOH3+wVHr2AabjjiJwMZ2FkvRX0Dw6urEBeyl/SpkRx
96VycIOe3KbUuuR/Cn2Qq+XTL5Yij1OqYuEWar7e9j3B+RTzsVEBGPdAF+02sDOL
/r+4YQOhplBcneCnTgmt/jdXlNejyWdgbZZgp0Xaiu7NO8W/f+DsQqlvDgGkBMqr
lMYzUYUHOJYZACuRoxwL+VMsWJHHozOHqQpODOQOzQL/W5udjZziKjZZ+dVP+GP1
nhUt44+euSVJg30xc3KbY4QbjSmhy/O1wIT8FU278ie2XEgShiOSRM8Sj6AFiuVN
piVehMYgQV4xL529bDkeVnjT8qpErRfRRxcMoPy/AeqVl2PQcMDIQswkcBEMCS44
C6SlqveKyTDBbBX/nhDmAK5Q2lXPmRuctdyw8Dxewerx7sym7BmzHdHQbcsyxscm
3qShIcyOh309LsJ/IkvGc8LL3FhhavBtAPRofcjSUVbf8SbmWkWRUyH8VjpRfjHz
lLXxPyFBSGv7BVCiqFozuERhBmzzPBstOxG+Qp7Z3qTPWTTiFSNgHblnGAkiHLHI
76TRw19qiUKxV+J5Y9tjA1lg74rgft2BpD1+8cIvt9f0ed8K8tnOwqsfrBCkjvF1
kqcrGx3GH2bs0yDs/ZgNFnQLKhiaTAM6oAhIIhAOoZGPWfE0KG0SaNj+8Ye4UiN5
ORwVLNVktmejNUzUXMnNluxjd/WVChd/rCDKx5VYO0x9WpZ2IaBtOJ92pGRt4l3t
ZwrN98Qao1amc4eO8LisMaLf6bW6cn9RlxNWftMNfGNaUXHOTcNNWLR5nvZLA3SI
/pK9oXWZafjWK3n4nu11El2tXZbiyvwha9abvlZE6wlRVKnXO4td94nQhJuHrjMV
FUUD7tDW/Jyj55k8uU2zYGIWNctcTOjpc3RhxxV8kGQpT0p1FL9/41z8WtqcxGzU
EuU962vGzDwYTQC4CekqVBwLIUZ4FOCAgBB7W6WGF2yyIpmCn+K82+GA9y+BE9sY
fLU0vkzs40deau54Y5IMs5tZGpiq8vOT7kor7vaet0JXsHOW4R64gLIcY5PLS3sO
ywjOv++EDhVbVCbcpQryDWX9dJFNAdU5gTumJCHx6UFJudgEz2vmsogF3Qqfhzzf
KqQ9epbu1Lm6hww8KueLSpbHv0fMvKwdNUv2P1MpalLNjPG9L0p/hQ2b/ggaASYM
d400gVcF2EK0v1QFXQQDglVCgCL77tV19jK8GfpDXMNlhnZKquVF9X/okuaA3gsL
sYat10mxboK77VZHXZ2LkujlC2BdS8AtIUD6u2Ykn5z8kxPPKfIxO7UuajTT0UX7
bmxwoxX0jrGSerGwQP1S1HPAqTHA0RPs7ulznHJnRW1lXGBZd8fbDUGhHOxhxiH8
D28LoZ+s9FBXjUwTJyQhLF4rA3jbZJL9ik/daZWCTsyXyqnsaDNT7p9l37XLTUY5
DTlUq5JAiNFH+e+dfORzsHkwalvhLN3mGn7NXIQAb3Mxi3kB52IW45hPXlgf1LPy
6T6pAqohxqODx5RYWgeueo/EtfNSiurtkszi2nBfO1sVDd3ArB3h4v9iRyQBsVqr
+IzcHFYHtBH6lFwVuez9izr1IbwMutKYKCAsyzwVM5Akl7gE5D/hjqFmz8Vi8ij8
DE46tOLYW3TStnT/S4GL598DqtXrGicnqZW6adSA3YOpjprqzV49k64nGFHEt/1D
w2x0KXpNaRL0TEOzVB80Mv2rl7H4uaE+2oEx2oEuljx10Ja5GxZsB4ZAHyuon/Vt
QVzJQeaFzbpwq7uCGpZFDtXHBiFNTCQG2jBWudQyya1KRtupCyAuQZWbkt6tr88R
dK+vfgmRO3BeHM4lAsKgqIhcLPIKk2lFYzG9SgJB0fc8pYZp7KJtj46e0GURzPNV
gjbREDJ9I7lAcZ6nEUdyqPtodWW1gwx/re0VrBjt9K/77ItF9D3lghEYxwr/yWZ9
Hst4DKkWDByw4yXtt3o3rA1iOpb9YBxPJInnDvvJ91E49Tbm9VmD6t11Mn8q8sOM
j5HpE1AqLNvrratq80tK2lHs0yF9aOq9nrgOZCmtAKPrOtyO2uCqFgk9hzjNShHl
GaRvWrxrRcHnlLG72WhHkIvSVB8LJUxhkYBcG7N3hGBgR9n3MrMerGaEV72Zkx6N
4CHoKdm1SXaMGtEEhrlsVMFQgWIOpDW6u3lJ/nl8MCERfPodlnYrQQQsAKDnXBXJ
QRrElnFp3YQbpl5N47jSfTrr5YWul2RGfkmK9Z2qIlCXyP5rfedWdMCRRtnLx25J
a5k4a3d59u0E92PBBOusV2E5WK4gT7HKsBCpGASehZ3KZn/6XOYQxOm4xSqeR776
yFwAA/ms5GuFNm3ap1NOyg5sLHk7xywuI/Rssrw2iDFkSNKIZGEmwLROPup53JAN
cQ9FGCE+40Wr5PYqxG5DdijlljP1HTqZmMs0vMFb5uKSjKIycQxvjpuSFhzvAvxV
p7vgXmPCtsy0lJ3peOvlonnqhfN1CLn+x9Eiuk6ULfBevy/KS8+GmQBtZmLy7ZqJ
/hzUMbJdhC56Yy+eQJ6aqMPXWkkd/5c86CxDVmSglhm0QrbZzVy9TIOX1SUmSYDC
OTMxG/In9iOS70wH1O+ZB6GFO2Sqqe0Sq9/Z8xX5v+3W8VDO+GQS06ouFTloQR2D
x5aCORlhPw73VGd5XBfa+9182N+QMTLN2NQHSdNAw4hH2MfJsP6oO7Ox0tSST2gf
VepMOxLQH/GpXG9Z3j9JSjbj30agnsHDQJOmewjq7pOL3t7ZsOfBSWUQPI811cOn
gOtG4XiJ9Ya+X+Wt+jAqnD8se+6MPC9hFbx7AVZMMt/4XHiOmHybY7E7cB7sz4Mz
scYnjjCaAax9P92Zd7FCT8+fsWV+zQMgCLkBjAmup66m2OVAQyJCnDeXDcoKV7yO
VXbJhCputQpGVipTt9i//ZrjMBdCiBShe54J2rPOBGhxNByzFhpWVgocPqz9/wde
5dmi14UuNDX62FZqnnnXLJ18NZDACNfYuRajn6BlSxImAZTldFGpOgGavh6pOTas
qm6lRD9T9uMdttS1hwjqCNhqTBK8DxFYoZDFYwV6VvuuuRqGXwtGDs0AFzzRu7xQ
x1T2hB4nOi54g5iWdpySPByX6JlRtloM2GMNJNPs1Olov3D3pF+dqCWf3xS1C7t9
u8a/2iq5sInMfVnP+GfXddQuSIfIXitzYNYO9ZD9tqYj8YkKOuS1scK0JqtxC0Hu
XqySKfDZI4RbxRbgqKbz/4UjHub427jXuWS2PM+WsDoJCgb24dsrPpJM0ZcvWMuW
wxRYTKQWQuFKVh6Y/4Ukx7ETask/GymZunJ/WD05PmfeQZBAvwbn/1CaEXs3D5D5
o5P30jleo4ADcFKofZWVYz7v7ky5L97D4Zieb+khJhSqsnW2znVt5foA+5Rfhmkx
v3jjmPUjNYE5BcHjvgmp1BK1uTrkyONYsrz00lW4SIOp7DfGhs7aDfEHjRrJvRoQ
nE4Lak3aESyv8/gA7kafqUh47vbqPAT1nhQaGFeDwv+A9boJKIaJCyFB4JeZNyS9
0ukSeKqT/JCu+xfMxDn9GZr7ayYW/eqPMS54580RwBOP03+y53N+C3eGqsLGVN/Z
pupH0IX/B9gLXaQd/Q/7YWaBMzgK0pKtNUls72hFK13/hJfF9DSAd4MabCfqidc5
0JgUdvv7p98XNSQlKoIyyawHx4Djayr9RFl29Dn0AGWd4BIYIsCswkcfZYLa0aRt
2Mu3f7lsyahS1RTDeKUYRElB0eahUABWbGLUzSId1f4h5nuptwz4KJPpNJg7Wquy
vbuM2pRaegMUiYaQ8ZocYSq7WGZZJBfWoBS5V1CsmTsvxm3ciyNWak9aJw4SnTbV
wOSZ6V/L/SF2Z0DjeuHIlfB/j4Gy+BIFeLouVuHnVSec8gbKAIykWkvhme5hYe+c
iQ56aNMTKY5gnsTWPE841RULgxlF6alPtQJ9Ts/UFtV1eo/b7bKfJUo4+i/VzOQ+
wRaWc1ZZCYkvLx3GBTYSfsF1SBcnRJzo3jlcGwon8F/2jEEBbndQXDBiARdS0oGm
lWG8cvNRBrpHn7OwsVPzlxCHwNLiwNsY6qs2+q/AT/kskhMPVWzVLegUBNp1Orb2
5eMS7GYr2vGoUmnq6vLhI3424+o7VpoDRcR1WzSsjEqq9+SeiFmHtwD1zEs2Gu3M
a+VHahj987sZFvto8eiaptF8GNc7ZK3EKpjlypW9zWhMTfApbabhFG9HDNq5WdPj
rFmX1Fzk6eg9qvaNGg0GAGzlI1Nte2DpnWNSMa0E6RK+1ccnGsRmdLiKivPXxff0
o9AzSEZq5Pi/0jPno04+2Cwnw3fZQG4gArr5GNa82gfvmQymCwoZHr+syiwS9dvQ
xLeW5/QH41hOpfSwJPC3tFD8l4yIP/pfxyXWDZOrd6818aGpnszaLe3jkhvVpMfZ
83tcd6pKB8hv+rnwdFbqZL6boB80bC5/DeLCeamz7NtrKBqljUuDzhXeaGDB7VM4
kEHXGL6RYQFrtww1f+3ccGB1Br3uXG/0G247spQijxdLvStLCjr5AJ1mHbG7B4/Y
vZvXRy1O0n8KaIOJO/YkIG1MgI7JbBjV5eIZpL9PFVAkElIZDjOU0PjivJMg57yu
856r3hWvW2YFDt7vCEzu+8+AkRjSRQ7L5qdsY3KuTsgOTEWuHGPdwAsFECzJ3dNj
FrFd2qfVaZ44q7Ef76ilEBJbRzf7NMaYNgOebc64vtveXLewAUHfIkWBspaGb2qt
qj3K9TTEdUHT6TlGiq0Kcp7JS3yV5L6ZwWGD5ldLDbdcHb0f1tiXTONDwXsYwA+F
oqGWOftxW60AIP3A/hTKdKNXCJrYBeD3lquu7ghrlfjm+BH9qwa0xKjvvOeRuwuT
1fYSlWR+rUekZ+0syop8tw==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8q2c22QVGMe7FjboMpP3FJ7jpICQXeVqG6ImT6jXSEqv
950UCnpQF9anHYCGLezhLucdVpxC6p6R7yVU19tg51BVIMp7mh5nrwmH1qbgNack
mQEipqPGlHrUftmi3qvDavBDY70NeIsJHbA3oFBLPD0AAwD93wipGzpTvAAZUT//
Yf8k4FgL85CXdrWwbgc3EqQiUjm3gNtTJuUPiE57pMohH09s+b5jOIo7kVTa0rhC
PBoHrFoR2YGNRmLvivBket/BpMGCo4sZ7vzvJ3JmNged/9wDwIreVjqo/0+EZIqZ
v1ub1dA+Y4YsQQvuhY+NvuKOKvAE9KOOWmpWDEUfaf9afR9Zp4nFzUhkGAf5hwEs
pCUs2X1ej/VZM+SnS49SSBUGlo7YhQJXVgUe1rQbJCVHnp1tZxvcZ44p6mWoDnKN
Q4OEMP6CL5ZG6Wdj1RoONbqntaaB/7AG8aobLKbhnFJpL59bS0W2WOZsdzo8KJIk
U2OboQyRAWHkFo4RmgGU+Cdj6X05J0dmkALBXClHz06t25AEY9hmTgsB96vnH/Uw
D15JSSoPoGzYB5y8geVqzq0KmshVUzhvGNEPIjlO0IcfEYzlS4WnS6PUgoLfYeJ5
u3bwG/KSOuIXACi2YcoYxavTkwnlmW14/1fWyW7pUsWOhhQtZEMxc6t1nq0qBrml
unbcBsGchyVIi7SCOFM4ypMoIUJpXg+7rLiQN0pBFlbLtmgL95xJbCN4j3IBiC+D
kAkWsRp+EmDROG2sPyPKnRhD5rRwcWBvYjgR0+V6tq1Bcjosslegk4mX9Wno27TJ
yy0DbFz7LnUkO0SISYf4owkZbFuw3/4G92I31tFHdDjc46JtYnegVt7guFDxSvWK
71Jj/e6sKoKSala2+IiRKJCqYbFDJ0itHQbtWwAC3oBtsrEh98Q273j63ft7tPs4
R6oys15lioPPuqqz4KhXf9hzwcB5Pdt651uKa8jtq+2WfULF5cLWRa2a1+Y3E4d1
RPcHRA1r+wFAaWB8hVdrIQbblEaVw8bLP1L2MZwTwn7gMVaj7nqmqfDCF8VGSVWA
SQwpLSG75ndcRDgZG75nShYhgZeDmPdyGkc4Liq5F4e54CbpeOMi7MbDWwCMcIwO
ggVqq8+DImPjIKtRD8/jO4vo8FSXBcxNi0Q3NODOqqBH4K6ZcBx3OqbeQ/DmTbgD
qmgGzvkc+bnAfDWr71q5yvNEit0y0Dts3uvpcg5mVytOMVYXHf010TD3orxlmnXB
mXtnwWm2fFW9XUyyrD06apmZOWjxczVwKQ5DKAEgKTOuRYoW8PKri99HkH4+1D/P
9zXc9Z495Z7Eg6E0nKuyVOV0+rUVg9FIgyPT/UxxJfneTFlb6MfIRi7y2WerwjMD
OthG6AkVfnJv5pKS0UBlI5JJMp7yOu9zXXMd5kFqoeQxoIFy6cLti1BDhWvsw95j
GxVQIuuxqrXex3cEs2F+n/T9FVZlMDrfoX7Z18IEtjFon+2j0rD19KW+mVbezSeB
UjjePDLYSmeKhY4S0vUUX4oqabelpa1SnpjiDx8cqaxLLX2RBikaMYf87pqW4rxa
YhDZn1OxSl781GRoOUIF8RjDiteedc5LwC30YFWsS/01gPT526UFVkYI8KA11pj2
CPxp4Rdfr7SCmHkHenKoHRrobWY3M6vSkqN2nUFEBLMcyujetKoajayg/F4/iT93
RNg7InD+Rr8yGics1pmNEna9RbQ3IFdB37XiWAs+xP2hDebChu7PmmDDPvLSEQ+R
4ePp8g6nXAzAqDVWRAGuxhYHrBhLbNC62uGaeBq9ooz7gCRBG4koYx937vfRjhoK
7LCvW4QWJCE4Pp6tI1w3Em9hnys8JjMVuj5NU33JXp8TJBTmxpvwlfQ8Pp4UrTBI
7aXC5itgcVFrgbBGA3O0RxT5j9vtjMt2mFIKqKGrSzb4glQjO2nwJrc/LP6Vd2KG
pehDu2ENYW1NpJb6jotaNTFg4T5tyQweyK0TBICE/a/kXNJSbNe1reWNHFr608O3
B6INaONRHNDoE7mngwaWOqeSaeJer2wLbtOnO9hsJfBXLLxOsGLsqvgTbP369xsE
oeL2RfwYPOa3M4laTHfZ5p3qntd+Up0o9AGkPpjjbV3r2fyTbc8cU3ffouftRnWK
hQgIcYSEEDfI2EpbmdtNkl1t8NoyfgIm6kZPLw/lmbCkhrFkSBZrnuyXbVx63nIi
umKpdFplnhRRiXZ/bcA4InNMY+aGFue81a7h2LcgczBHIiUvjHfP3UbCziEMCiKr
d6co4vfzhzf9uqejNnR0cub3kGDaZNheQFCucY323rOCQKIhg9AZmnnpMFh5Lwyc
rUTxleOfEYIOUYIS6jaNmlHA8XGUtBsN4gPbtV6u3b3gMbITXCTR/ksvTjq4lM7C
rk6wSPeDsd2dfEE3wUa0DItNIgYPO54WqhBvc70AjQX3e6mBwGwTMuqX0fxAJlVC
nT7cVL7CIqm38uEDuGoQ/njN6P/CpQICirL3tBjilP17vxpEiRwCG3KA0HyTl2Gr
AtJpbQvoooVX7QdOG05RkOdfu0lX1VVftRv/xghL7+oQ1+upmqSH8iweNbiTKA5i
kvtFlJDdWZ4nA4KRtmoVi/3x69191krHMC+Z3JrAlDDsBOUbAj5QdsFdvBBTrf2S
fpQQ8BKe6k/9jIZ+ExuNmfawx4zpvTWYrdqEHJ4oG7VXVOnBtPI6EUVnfJBWxcKU
/9jDZ6veZzac3iMoOuoBzNzZ/IMw1jXHc9wUgeOb9grEQhrcmNFVTf41uAxYaY/S
CBkjPAo94WzXRqBlwGi9ZvevOpMA2Z5qElih1oakeZw7WZ7T4mBu04jl+Pc24BGg
L27896Py74pFO+C1sqnBrx5+u/KfH2I77hwrPSQmYH8DxKYOFaAGksQzJNVXqVdK
MRrhynA1R1uTjTN0UP/mFXoNgsVcUADF9vxYGqnWGQ/6SbA+2pDSuiCa2N9glPDp
xZEEU+4xxTGdqV1p32aA8xkhuSubVsM05koXBWhGKyYBJNMZfBBsVLHeH+vjxWbo
FuyIZkOx3l9H62oEkRsG52+2f594s5tDVpq4JOXHIcKNueGEO5t5Ca+nOwbBsCG2
iJz31C6qkYuBPYqPDuLoIC30YdxVYf5hiBgtebEjesQkIs8H+jvNxo6u9k95bjZ9
3Dn0Q63IZztzby7OGuwugBINm7oDHDQSCSVDIVIeGeDkNvivh0FseByloMAHJInI
NGrZYpEjeKUgNFnYpC4NPXl11T4ckJiLt+O2sQS2gxGchdVwF1Yczf4ipCSmh+fk
YbrQxSamJrsSDmgEu5XL00SErA3jOW/eJ477gYjK4yz48LxzP8YSlVIxQhuyBmzw
mQzw5qczF4rzzkahOVuUz49y04g38A0wHaBSsnKOUAlGAp/Ql20JUtgG+CeK6OrQ
6N53lFGURhZkYjbJ3Tvio8iNqX6YOTeoS/Nuc2pWSiiJKN5DPi5LxB/wtb4oMmO7
lmw9cUaPnLHR2gfQxCVZqB9RL3HWecfasSMUHQbAEfWDCn/w+Dm7IoUWTXrhAL+8
I4uTbSvRmemW1F1bj721HOuZLFGDhUVqvkncMw06UhgHWA97dxPAWCDDiaujZimP
LAhKaXt/02OZvpjUfRpw5MazGB2jMmA9Tyow6HnKeqNPyplfAYuyOZ9MtAN9CSVR
LdQfQHcvvioaeJAMnifUI+qRdCeDQ9wnIaFaGT24FbfFPdrGYMH0Eoui3E8MvavT
ucH/4BTcV5SP0u0cpNUBqNcn7uu+2DQqGw9mVJRcKW1J8SZl16C16+K90qn90/Ex
WCztrt0W9QvY4qkYaamPaQdpW2U4bZsvXhiO/jTlCaFZ6P2ah3OWlWb6DD3bQLTb
23YR/fABqmuDpCSl86BuXvBdgYs85RSiT6OzbfFpRm6A+BY1aAbBr/xBlATuMsvt
IYz0T5sVBUwWYEvnF/eD82ZkxWbmHW+i/tPyIZ73AoXVFk3vJepZD040N69duCPC
WOxQx4T5DKQkSUTFS7qgIh9CvMcC20Lz1i9o1yRz0W3yX53jj5kuOk5oSjuMgTGV
ifqW0Q3iG7tTrZk1FiMCNcM6UAFpEed2NuO/Vp6aY6yKAMIMyAVvJiRGi3xayid+
4L7mgv3mboKFjgEY8sbyfts3CL6osx1rgbryDAyk0fSAjKngV5iijOmCJBORtXyh
QHyQUZDnaa5E3v4GpzjKPXBxdOkkNbqAst65iPHbgNTeHP+HEroDKgEi/hHQ6n0i
OZRrOLqYkF1cW8Pkxhk9UJuso1sHnKklmzxXLXZ4ge0CmW0uxEJYbr4f6vewAKK9
QIjVVo9zcArvFLwrG4HM0WkxrVpI6pBaZ777eb02MYLV3VGtjMXJ97lkxbmjAIks
BbXoiEhi5xQjDkuoETFg81hKCyRha/ls7LyMOccERMrxi9BSYDHU1eMCRrZhUXhr
LGA+H90qUllGUEZ7SAIdG+dh3tkFJhrjXICni6CvVSdhwW6HzutGiVHqD+tQjjdj
06nO4azHkerCWeXvXwMVypwR0lLQlpCsECr9jWEVeeVfS98VUJxBDpwpmZFuDB0I
KNfz1M+x3524NWPJZVRxyN0/XY0Yz5n6gZm+x504yZ9PKBnNg2V1gw6j0FWKwJqH
tKWXCTrtB0gm97dwagG/1aeY2TNBad1XJSG4NIWE2sTga+EyBvrk/I/jZqmx+zZu
gtXob8ovAghDeZHGi1Jg1mZegUkrjoNDy99HVe2Ge0tGmvRfS2YU81bYjN8aZGhF
Yc0b28OFnbJMpMjsA4FjUdHFVV6cxVeOrPVSjD4P7qbzeB1Rvlc7tFTLRQ5Rf3De
I7iMnoDkA49LmilH3p2AqT8+KSjJXZJb3XftK124xj1iQnz8snVCW/Ha2piz3pT7
jqwjmAiL3VjFPAkZYj65m4H6AltqenxtmWlBm+zzhyahQ8qxu+3MmRPnOWIZEavv
sCssWJ6yUWku7iNzVYLEz6zmyy5qUzXVLPk2p7tlWVImaFaUOOKYzfbf8Xjp1loD
sMJMKLUY61gplvYkgcwt4TFJq3h0K083thXKOEn/WgZxY2BQumyNBoRe4cCpTV8r
ASpoijuUhq5FZLO8ImrEehB4+QH9fL4OKXyrZ1tz2JNHItJNgpH84I7gQBNbZsgR
wSl6aphz6toPUHtWc7zENI3qjoW2mnJbMAfSI5tVDMaVRK4aNt/nNLWpGScG1nWE
/F9JkJC1r4Fcz5y7rxNzF1P9wabwToemOgav+6Bv6WQ39tlRUs9QxVX0It2xMkR7
IcmjNao7T9hz8gPlJrBSu0XYCG2QQ6t5V2dGyN2y/94ypWL3G9QeP69RK5zbqGxJ
Xn0495TUtcDrHFRUbEdN7T5o+zLWUMybrmYu/xq/ops84kRXZG3xxyksWgkx1po2
ykm5SR9tmuXEhrcpZlJPRO0Kv0GyTjE5JSmuqhLYWAz4B28VATfnWqlDSSfajTyz
iPxJnRKmsWoBp8cWcDrh+R3HCcf61N6QWPw6duAZdXvdN+VU19pw4y6gqgu8UdFb
LiqxpiC+OzNeT3Wqe1+80L16MOkL/oi6XctI1KZMbh+Z5iTdUQtMkypQDceLehXY
+2VCBmw9SqQqJLj3xdKUUBOJPNikUBYiVIhFGSTDrdOLOiCI2S8Ove2CpA9gEkWo
shQ7bX8iR5OaODR6N8CUZYDMYNfPBu08wreNX6r8ZpywGK9q2NRVpje07On8WPBD
l1roIXOgIAzDprmUQ3SV17FWZkHTyDGwkj6vRW50I3vN5puIViwPNRvuVvU1P/SH
A+uP0rbRQ8MwQuVc0OYEyuQX4InQDyJakkBglP5M77v3DXJWYIpI8kW1i64a4d/w
oog2DyIUa7JbI0VdyWV2IdChfQ105s/oX7LdgEwSd7oL7pC/AWWzOaemvH1xa1q0
UqhFoenF07tzGLQMXSFGqRcSHdwxkR7dlm5FNOGwp3fBXASnViiUvdZjudxeNMWM
RtmxCvEAawYdlnonkeuCZ08W78RCarWbjl7P85dy/I3DEzCOeVTmVVQU00E7d5YH
pUr+qObkYM1lMWKoepzZC1Mq5j5fmnjb5uSrq+sMn40xyTnAxaKxjWH2QV/CTUwq
UgtB6R0e+ls5VEPZaV1XH8EdhQUDozYCJIZh4pK0L9Pstx0RsQF0bsXdPuNzWvRJ
biwNuS/qiejHn3gz0bypULv0TUIeeRE2rPCWFGaVmnr4Gnq74UWWtLX2eLnQuMpw
K4zA1lvV8Fy1JjS61yYdaJHyQJw4pQeQkOPIr7mddv4yfTrOfRg5PS+17Fno8Mvi
zCrOzdR0iWm9Ba1ZfEX4Nb6uVN/e3RBcR5LCbkOCX/gBnIsQ1XsVHFSpzdFo44gj
W4/NIrc5xWAvCXsMD+gmE/j4mtpe5/yquxv9j41yLyfvSv7GEKRWVL7mHt0wdzBP
RdAHW/c40b0d2b3Hume/8P7jbuSuf49UMGkkKbnloftSkSwNZWBPDi4sIMVxVWHl
PAiXdbpBRgZ+eHKb40BLWaKTkldCfYBi3O+AYLekeN3lB7hvPhGJypJNQmCQLwj+
qbC/FhdmFf3ThkxwwziDFG96xefVt1laHKTTgnFnbYSoVbS61XrawCHVJZ4s01yn
QkbnvLjHEOkyuEWSlJc2PLO2+tTyWQuYkw4rqTi9xVw4KkZ8Y24bLm+LJBo7s6YD
NWlO8w1A9pZQcDAYKAedgoYOzBgOmqGjzQ/1bMOMrjOMkadxwBdXXcjAc6t74VNo
/uzvPFyKC8ALZdgi8cnKcu3pI8PMbzqHy5JcXyA1cbb6uduN1sjjvWtqpgwzWAZA
jdFvl6vmxZIJeUJ9TaR3jsHawynTVbqz9ofJ6wLyUhhS17YkybR7ewo++murUz9p
xOyPTl7cUgiozMqWQ3qwwWX29QuQ4MI/eF/hjFEu+r7F4rrxnJ50s9rm4FWB/TYl
TAUMMI+cntJsITk9kwUMUtQgiK2K+Pt2fDx5LneJuaSap8c0qzf7jyqU7zf5RUnU
ItiZ2C7Efp/JAYsPQn8NFkJox/v13zt48Fg4e0bD74aNyhZ1KvSZY6q1OK5F79Qw
C4zhyw3/K0EwZGBdN7D1qmECGzgfDBMA1LAqsb6iNLXMPoEQsgoJbceqIDQbJOre
GGBZ7BkYOWsp5ioMQ3Fzo3kdxe/sRd8+Gd61M4Fv9sJeV7pMVXPA8yKiuSfS9KjO
KqyIo5qzsQvgp0+L6xTDgv9JE1lD7744a+TLlkoKj1ysFo8n3ZLM9ZYpRiE9gFa5
3hO6yLic0087e2GWv2eTVr3QlLvAIkUsnq31e0SuKY+E5MBX5C9kRrdMCElQKz3h
zoXsxCn+cSwh9joSDGrgarbSE7Op8K81VuGI2r7QagMPGJ8CVRxgfdHZi3qZnppO
wM1ZDUYKNeGIlm4RjjwaZIc6Xq2wcRp6eYzswn5Y1ncxF4dleptisp0ulpF/wMeb
XZvLqiCX9p3aqjQbnGouUqW1u8EkR2qmIkz6ecKqe9YYoOmAuG4y/PnUD0VfPjwq
SX5C64GZ28VHJm+7CRpDBf+ZUjzkAn19h35OVHKc9glKDQn7TO11h5f0h4JJFmFH
SroyNHcm+1aPhsLHkdP30XV3E7f41K6kdbPhaIepoFzr7XCNAfVo9h5XfQ6mrpfE
+1G+ioiM9qFsYU7qbAIyhQB/GrtcwaBUDaC5Ywa9AsZ4SNRlvd1cmAJo0200QPHz
6DHM/POU30zu3XhcHrAoWtC9oc0pfoRiHCsa5Ro+tdFp5xsLZrX4fswn1Vn6P3uq
Llyrt2gWphb8sahnNOmfWnSNWWzFQ1mDO6WvWn7XdOVrJRTilnBsVVpPk8dmZGax
5woOfcisHm9ADNAUAS80xn+xwgKpUYrjQPp+vmDWdgGjnhO4UQ57kIuZVArdZ8tb
CqhxARaZefTNnQ9yZhkckAJlYEypysVty0F3e6gT4Zs7Mr6U1c6RBtUj/wwy/Uig
UJT4MWHhRIR10qKPqsK3PjonKNA9ZgNzpWo7LrnrdS8wuzqeHsTzoPvm6y7zFZ6Y
Ac5c6zsUBumxn88LIVznqb1+I4+5/USTMjsP/vTfN4H6gIz5aVLvGCqxQ62UX+2A
H5aCFpXh3EaGWC2biQXdpRNqUheTfVj6k9kPhGW7sAsfvzrZRFyucaUbZ/h1j8F4
C80wzCuLjjc9eeftXwPkM2QXXRKc9EqtqkVYlQVMpjXoIJwSeZBOY9c2Y0qQ3ceq
I/I9nvkid+R091D6j1DzQ6XUwxqTw8LsxM99A4wUdfun/AA2JeOrZMTwtWlp9MSy
4PVGYm5aNr53xfGbGbZfO4ddj3/CZsMK/6K7Kn7Zlh95YO3wWAudhoEq0pX0uaHc
08ESxOWipzbwzf94MvQ7w//DSQ43E+1ZU4NtFvjGKSiF2XXR5+RixKXOQuRjaDDW
ncCnE+rV9zINJWZ2eITiTp6Zps+3yP7qEqZE+Lwj0RZD2GzfKd3fwGw/CcdCOOBy
iZ4N6qj/lr6zbOqc11NFAR4T10bbcvtS4t+sGHL+ObULL0bjyGp7o2qsPAST1kvo
LSKueFBm6V4gVPGOi/m4SRZk8u07dVs+hPYbGX9OHDKpdpBGlAzCPXY2QU/Co1MH
UD6PWSKiYG0UuxB6sF63l42JRAME6wlE0s2DZ+I6aNjbcKWUp80Onf9ox6DwUa9D
61zC+AIuYPPYRWCcrRqU5NzSqM5vG/mJ7R9d9s1PXll2U/RAgisk4DA+9oBsdpFm
FbxLicxhSH7Yw/JmJEx/S6oIts/Jx8hV3Nv2hYIkb4EzzMD9GQns42rb4L/9pSl9
t/1OphDIDL4f4NzHpvskbxlVsPiCcACjO1ZlkrwJh1s1XAape8B8vW+KHst6Y5Ak
8CA5D7lLAMri0Qgbj3uPNxd5+4UkzH07Of5xPqStRkZC1RnEVnYEQXkQNqTZkNKr
BNJgwhY05gqqKvOje2tub9YmUFd6K42mlrMYjof2bVZ5Bv6yVbvvsb1kfl4XR3H6
VCrCj6wm9vYI7DAprS+t+d8pPg15Rj89+ILyZGw7KFkVUlPMHoq5tDoMzboVg8ri
i6h0CH/i3GzI0Sc0acZKnu4saUxhm6A4d2+V0ZRKXES8EkdpLIEwEc4/4LAOP9pP
kxgg7f3IagBC8SLcix7iu5GHAKtwhL/66RvjEmHEXYGv8bBXtTS/heJ+Rjg1lH8n
FZFxbyrQx70nGjkG1/MSaxV3iwsR0seFVZfFWV9Ms1F9RthQuIAYyoSPR3BLFUNZ
GaCGJnkSyDBrWo4wNYqMiOfn8tlJQ2qUbtFkaDUlIEzmOHytbVAROChb7P2fia23
ya6Tlxu29ER1GbguGb4kXuFQzr4a+rr1VPdrmNdJtocYeY1lfNLz6TXb3GLxgWy9
j13xutgbTMbeHMqZ8LHKjvxaioakEGAU+SwcMEs0vErUC7PKtmDcCjm16PEpPqG8
G+O2LLnoRcDnVEeVJDeWHanKXW/H8HfUTNe/B24VfEtLKBobAiEf4bhXqz6frGGG
qyqPDc1vl/zUi+XOyezNfX5cdnmUTMBJVdVyTA1la418U40DLbsbnzVZebyh6NBT
0e+JlX4mtbIS0DXjRBvbkNrfhg53Uca8U/+z0clY/R9l54fzECf4vJW2g/OyfIy0
suAygSAhmVbOx4obuTUNeh3j1+wbWzrEv5OkaQ9cRVKE9HCNfKQFR8QPhKKHQM8w
V5YMUHPxR1+RK5nDMWYYk1V12sY9YPnIUsMLX4hl0yc7ReUVFA8h6S6pH5Con29r
csNiz0r4q5Y5H5JTcEmbPlU04xdqnl7P1RlBTZMvJgf0ge7h299xMeMwGQ9tz2Ho
N0HY1XmBTSmtr8qcm1OJ/sC4VP2oS+xVR4nCjg0yTIFH4DGcW1hsT2WdAckLI1VJ
nZq+XvVOK7o8M8FRZ2DGDeB+DFkPTVRbddSLdGtcJMwvV9YsoGjv0F2C9k+3fseF
LaHmRszUHI0JSocf/5F5IdCsuPvjjX4Y6q99E2LAbO/W2TJdAX6Tn+Hemer2jhvj
53o9e2HIcbX18OM3zTdC4eFf/jM3A/I6QYhFAvO7raE+o/OJUovqNI+e+gfje1nd
EKdhCgdv//EVLOkm+aI5w5MVASn6ORapMcgp9KYs8a/mAQr3B/GdTg9fB/KnNGOz
fDV2wihW0Iw9uk4SggJyI2VGmiC6zPtW0ggwGCiZeg6h+R9oxxVlx6KCF6wtkatt
pK0WJA7hwke34MVwfdDbarEYSQv7kEwOvGjdg/vpQw9ikxJ39faY7y86M4OzDZKJ
rbJw/9yak7AokJNZdZi0pSErxnJOFbBc71q1A4BPUndfEtxVOZPJ6H2kE5ZYIKgN
7v6R6QQBF6HOJYVEJSWw4gkF+x+/1xJnBufg031PPkGkC2wPNs28a+Aa+4lJUU0K
xn8MsBC1i/O0zgBJwrsuuqbyDeqVL7G4gOqST5qPem/4gNYIShszfL2FrW2qaqH9
NgUvjZJQwnk5H/5pcY0RKfNB2ecWU0Ue8rmbI9oXSOdI8wOsgkShIl7lo3T3iCqK
TO+CHzBISp8dcYVo+IU+LFhA2TmeW65BOkC77g2R6p7JlK5Fog0hoNQDTIdfDJAK
E4vLJ+4go9/HgjESwPlywuBPH6qR9+tluVLYx5vm5nB7cf2YmTRnL9iwD3mFaG62
AmFTB3//eSC4jRE++ay1DLv6OuH6tPev4i/EVkcQFPmhVrUzC2ItaTEfk7AZaF3V
aymdvUqYrWoe7iEGaMYNVyeQKgRZgl5bMZgO3Nr/FuFoN1hfTNZ8l6iqAb+y6UFY
wvtY7cWHjObGmYaoU+uY1XjD97WZBJ+vgfB1m93IBDMO5TuPNrQSb3XD7QhoONf+
8BcZWuz1SzrKSNe8Puy6wMclE7n/ICAy/aPA0s3HemW3KyNto6p1nyuzqKwLjQ0R
+xu8sop1WgHoUn7ezLaf7s0NXb+SUN+30gWDVxr2ZTHkZEE6YZNK8d30cpsSukHW
93n4QxCKSXRzm7cVHxzgNpoy2bZ6UyKlGp6VeTe099chg4WtIUqR0FhWjTeGmTt7
6gT9l/KRv451EZnDMtZlhwuGwIh02WEtnxH0zk/u5G0DkbhapmTvg0Cbp+tcTFvQ
6ZzYN6GeCu61ZT6L963UtTE+HjV5gbucC52+nG5JmKS3mGTovd7/DZer8+VXjotp
y3YWJyKmSL0uE23fQ5tW0HE5IKjoZp+VRCc6QMoM4Gg8RKms8Yq/bFi0FOQR7OMe
CELhOLopcTgG9cHDsA5jl1WZ9jePyiQB1PqnVdYVhUBuh9U2sJQJ5zqI9x7wmWk9
tH0XHUuhTBZULCzq+ty1gk/rEiK4kdg6GIuS/oQm22fe5RPImLvexht2tV3g5xTN
YMsPI6ny2PZ4tDZUwa2R92N6lGakekIh4mkSu8cBERBHKwS//6+se7J0vA/PALUC
v969/8asBSiT+K90uTAGKiWysWQLFecRKHD5/Zluu/ErAYrFHfmFkY+/ovkGddH/
B0aaZEyS+lqhL31p6ckT83h1lzFb0aV8MABHLqKkzNGmhAq/ClWiMvIe15q3Ap7r
2D0lOdJSlIimeySCtXhZk0gRP5RyOsc4BR2w6z+pER/qVvFNNdo/McGSqYmr+Rjk
LHDXlQ6q/YJ2Xr8TY/+t6V/hkd5d9b1wEYWCf3vf3gSEEr4isI4oxLKKj8trzISh
Y8ZFgT6HigHk/eI/Kz+F2LleXAQ83yRPNxRITyxL+/U80T3j/RbjTh7lJ5TFnYzd
q+UKGkvFKfi1P7OZtWfFhwRX4vxeHXs7PPz5WA26FGS3WUHylrL2gPD+yS+ijeSf
IUR94vxlg62YVxQhOFTqWdjdEpVyJyQrjEoXrShhXdG4DTpNxgDPA2ht3OwFggXf
cszS2nkdaOAnvmFvkOEoSnKnQM4ZoNP3z1MB3NL7PQYwqOHnKwhAGsTtq/3zGvnF
yShuCXBApeC71SctDBC5D1DR0nD10VTPsJp9vHdGJc0n3M0BgipsiF66zZo/ohNd
xb8ziz4VpJdm1tcr4kj7Ct9Kyvh2P0RIaKFj+BtFrpr3XEA3dpQSQe2lcw9bkmXn
5SBxBSCu6JSR7NT5YXAYDM87RMMG+rl+Mu5VeQQBWfrmBB1UYDzz9lbz1i5ECaM6
st2wWh5f78M5GBi01c6nBOnscsgMcPcZVDh2eRtgodFrqIKcvngkIPDo6ri3ycpj
AnpO2XOucPK7ob36/P8SXeXOw27tbXnrkTvDBEo4h9CF8hBZtjjQze8oqjuT3aGT
ecHztc7em64LpckEKnkYqBmFaRt7eR4SVMmAwS5FxbJTQ5+mr74YVQOvdIpFO9yH
LjgbXnGFFpPuJv7oNH+rIMZTyzhMQCeAJaB940Ud16TCw2FoaydXBhGkfSF9NPnm
YxfJr21DQeDG7nqelqvBWOyV/hFmM/WTbAmlNaLeQPWtECLEKcQ+wNEFDnbLeAwM
LFkO1vXWnjjib2g2O5T+pUf7kRtN9Hu6LwIFkmSRbWsB4wOxQqzebsP5kC9C1iN3
td//kzXc2qn/Cq27Kguhfi0yXO82jUjkeamzzUhukr5PFZ9Q9zUxjmY6RiMNcIeg
lH2p942BvpTt3ozyOgIhDG2J0Yf2IGYZ8JphzkXDBWYzmXz9P5M9gnoL1hr8Qbm7
FxEmB7L6z9yIAWcBu8NqiHzQ9Aa3Sf1+CFiTWLkZwX1OagB9tsrsMuHIbVcX1cgy
Y1YOj5jieZSvls7murdadVqTsWylGe3ElX8clhH2+p5u5Tq5KuyXd4/FEfxa4NKd
u84theuGNOOytONC/ftfuvBFDttE/Gdr5WaLJCfAATvynEvHejLHXOghvbsZiBNE
o7w+TP5yYVMiF1WvNvbvfFrS/ZZpbgU337e+WyTfPbDfH2ym9BtTJiTTbi8oZnM5
heORVWpDUu5bAU64nA3UNgxzkriFXZZPUE/vEgQo2Opx6YHEEqzDumF1EEo449F0
XYAYN9g2y8v6DdoWvMji3g5ZrqcIC8E3HyDm8iSJq3Nd3l1uM0TnAmfJkJiifMzu
ima32DqMfV/2SyHehFyqrfsOXyrDRFK1tErz0ON+QuHlAMTUo/xQTM+2oyNL5MmI
TCaA4ojkWbISK3KAEIAX0dOhxsyBDNLY2vC6u/qBmgTPcrx60DP6q2jNCaFRQSQM
pvIPMWJyBeRD8Y4k/X48cZpPyXkJUl7kHhZ3EAjgrFreslEwgQrjmfCH2V32YNFi
07CYVVvax9FVzY7ElYq+eDDiSSK6mr2pC1irtuMLZL+JCrOhirYW2nqLgmq+0+/m
FLka2+BgBd8MBMnaZu9bm+aQL3lvh5qk43uexLvboarJiagbqvIWj4q4zJSS+DO/
XOw7+x8d7+gHEPIB6eBSWoygabWsZ2gJzbB74Vj8AQaijtUwP3fVJfudZutEKpqQ
SAOSh4pNvC3N6vSptQs1KG9wP9cR742gwGWg9lQuJzon80IsvR2bUV2RBo55IB7S
XIpjfWmbbCXlBzKbCqtqmBS8j0K4yJmBBKwuC/ShCwUsKqbrvoP6ycwLE9HF22vW
ypeZ+IULIcY7o2w4V3+OXwQQyJ6FIkWfLK+01jDSTSIaMDyq+uvrco1FBN/wdRSq
P/w+7GmrMWPdWVI10pbmgu4cqv2wi07TxcwDawwNNV0Bfwu3tVe3C8D/KEiePZf8
migh/iSXjthJBPVFVtPrYNEWWfl2pvmYM2AtxwyW/7gLQG+h14F1rJ+dYidzy3FR
P7vuGObqkiUAZ9RsmUPBlt3WE6Ai7oY9++IEmMdkK+qQUvIG/6/KkVU29jpydm+j
0Oor5urfsdPaCtUmniP2mCuoGqNTeXCUS1KxWEiFYhfM282PoueeZ26txu3MB5dt
tbG9IdRs3HzWjeXjUG9iNQw34H0YTQVe15NFqzfDx7jJZYwnE1dGClMR4sTKqQNl
pf6pasBM/n90d/O4MDWdHIvAdlxko2sDY623CK7Whg5H8G0WUzWtwgtnw9F8kjUs
qRjW3sE0kpsMwBJALWBjjU9S//OPBXnbDanQmbNBjXcesRCiadWKTXd9yVddFRXI
rcnvCZDvzlorRFGM4pIKcu9wSs77u9zBDAa8IaUP8Id8+NWI5SERc1lJI2gOE8WJ
FNpy2BYlAa7crsc70Y4niFvtau5xT7TNJrHkP8bnCmkeAT5yU31blIyCVfFoaAyE
26uhJb3PZIXmbkBioqBWqwm7RuSvBdAgB/U0S1PcG3vOQuAtC32X9jX8x4JvVAji
xvroMhH7gzFSkAjdWhLCtVzzycoWI4jkTFsD80jvL1k+n0dem17gGqOEg9Uaw6ju
8CuV3TGd1+aXxWsUmAoAGXKwU2t8IgeulYmDb6sPwyvXQOIbOg86m1mhkVyCPKg3
dFUcVMNk6b6fAw8Eq4d++d3dd3roO5W02Qsa2W1sjmlrY6VBRIgEvvtekiYNcNsT
YLyhow3wo6oCAQyd+Ha2LzyqsK52jOWRB3JRkDxgGGjvZ/sb3sF1MrMLdIRyRna3
lDlomuLtJN050rlxRqGmfB5NEklPzz65sDnDzvc8umP4mYQ7h9UWRDoWjKOgPkOp
TQo+TkT1cs71w/XCS6q4BFiA1Ps/5WHuS8A/coHIsqjXpadOy5lKO3Genb9yfIkq
md/KfMphI5B0DZs9BdTpv4FHy+0gt+0HKMi6qjC6br8vmCFKP6XsOESt+q8IprsB
WKmThiam+4AGkJ1hw6RXljnraXKB1yNok+ZCk6cuKT+LOvLR357GX3Rc0E31+bo7
vpkSti9LLCtJIar0ixsK2Mca2HLWEUSQ9GmBejT1UcmvTxWrNdZCUIk8yi94XkXg
ODndhhL1U83BDWc2c1Esh2VBmgoM5Uy9cfx/orDklR8LGNoGI0lBrsrYjm+IcLbR
7gRLqt5DqP3HZJPsgDnKiK31GmFoNuD8Bg/s8NDsf4y9qmW3KadL97RlkpEnKI+X
b8iJlvAEI2ckPFU3mtjoj3lt1folZ77Yr2PfoCxEo5FTQsWT7ynaZNqoCmQxoJf0
wulqVQQKC2pLsIg95uxEyfXXcGfp8rDrkOWhceJG26aT/zr9kdwOKu3NHijpWgKM
d2aTgX5UZWqXqP2+f3ZXfVRYc9KMYoSGUmJIX9Mv2oXFbsqvF3tlddnGJaF+sTyP
wK0Yrqwyj//ZA+Knz0vlKB1+6J9ymnu+9oVGZnAZlIySL//UUnFQExXtN8URi7si
KiTRLi+IgfD2n8p8YS81JeRcfa1kE/PUco0Y4baBWCFCe0RBDIUIgEHLDp65drfB
AuT/M7xxAjCEX5SGS7MqS7JvAL9Sm18E7uR+3yTnlbWocXAc055nPXHkfUcnxhhN
MQ31ERHgf0WqKYTrkiDFKVH9eZvIMwQHunh83ocbfHRTo8tqdwpM5qu+2KF8qJ1o
lox9zepM37mAnJshrf6BmCo+CBnivQWEXo8iyVAqLK1Tl0ONl7LL8Bg9yWEPc7LK
2I6rMOS+GNPmfq1iKlHmWoV1dyx/jUYPFITWEAZZSNZ4SWHLQjo7GNVOjPJdeQFD
lnknd/uXe7KtRBD6pD0gljWN7fvqml47pX2riRQC9agJ9ce61L4Nq5u3r0FAGguF
woRvw4b98yAk8HEP0CwpxPR6Ubi2MkvQeNrGO3mu/plOraN6gnxHUsV5yCSHnrEw
ct5++EPbSHgjsmwMEzBV+2109Y1OEaVFDJnpv7CLYv3kBnuoTV8QIXprDnXBApiC
J3zidjKy3Vuf6XFBZbOZV4gGG1K/U5sLDm5u1QXXXIhS2ByM8wR/ttg8BD75FdOQ
P+44oe3ypFT+8W8ySwEWtwDqa6H4QejvHovudQb51LFLHz43r8tQJGXzekZ9KwxO
S+LH6NPBPhKEydhtCmQGW+uxooSGYxgSHVN3NA9ks4ug7wEcxF/cu+j2Rek92Aro
2PJgbdDAc1Rgv1De9VqdTQ==
>>>>>>> main
`protect end_protected