`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
K21MooLiMCXVPibvGUiGAVgJmvo94IpgywsQresTApRakLU6RdkFB8w0W1BYKtKr
+pr5hc19ER+4RlcFl6tNip9AUDoUK00t+MeqUpAzLFVlug07bkVR2uORoVb8dgFT
B0FZCFfC9DCKCVwM6zfbCmhsegcR6cyhcqnQA6gU9hVcK7NkydnDZnfDNMp5b3Ed
LRVjPWwFNalqwI6D6Xune4BtUSa3DgLl9w8gguFM4x5yPp4yqJFJIWRRuZWEybX9
fPFB/VCsVCzU4t8QIzU1Fu7vWzigefd5/V68uWAGVBO/PS0kfxCJIkJtyzXuUe+f
WuSz0vMb6gNV3Lvm5uBZBfns2XoUbjKKovhssrJTpV/fFQfxxSS0mDbyMackfT2w
6DnKsF6Dq7B8PVxAkLh/ISK+OKrsGbZx3F44PelQadR7KQ3IirGE35hfrUeVy6rM
DSE2lRAdA6UZT9sVX9/Jf63y3Xua1F1TJZF/7hDNhEi51uw8YCshe3TUAQNhlu62
wBlBZ8Yquq8SFwvTNoAfZjjDC9J93THkhg02DOMZK4bo+k4U55p+SDa0bLZXu8B8
xJVBE9Fjf1Y3UrImrbqTEARNchmxU49C28g+wfP+lDy0EUl38kyZXCf/cZCACo9P
cgDyPRYLn1uHhHLPFmuyc9jpmXvPOpfiIQgpeRThxbefo7v6nFMrImzf9Yr6rNm9
lGVUmKYJv9b5gWr54R3rzqNAU46vhJNm7JssYzqkRa0gTiE5o2Y2GmrktpNTV0qR
jzqk2mFG3HKwPPiOcv43m9s4t9aCU31l6d4qIh/EVehR9Z1M7Dvz6eDFxPmBREZX
xAlPwKsRvCF1HIYOnBitSmH7kvcasTXh/u+ATEsx1HQLI4xEGIODrFvrZHpoFjCP
SYgSN2OH/xjh8i2ct8th2sSrr8GvQj2AEzYc39WBStYm617usdChIj/xhLy1qguh
XBAgwIEfK7z1Qejc/d7uSupPUOIG9MP4g5D0TweTnuVELccD9xa6OITTiiLIhISN
0gxcYHovlpxnBTRFikXIN+VMcfqGcLSTDdkkjJIWZAXjtha2odDkJMBbfDjEiVKA
7pcZW9+xTvzuRJ9Ix8ytozLpjPBdikkmZDXHmMzVRM+uPqQ+ZzDD+ZU7uYaNPmia
mVTS6/4PSXvJVfhXHYqGFFT7l8uajTw4oe2eAZTQdAvxIqB3n6JX0dHRnAQDowGI
/76WwqR27dirfwtsahk8wg3RcQKk9/hpVcog5PXHezBw7Pp9pHxw5OltuJpNdqFl
TwbANph5pSLHPebbnMxsdvH+nf+hRvB4/ULSwNXyrk6YLzyfe4NfnTPbAPQc9hXS
b8FaQXr2BZ/9HJCg6hfXLA+8n9xbQuIiPgaVCiUjVu3yODrczOgvUFG42VjOOz1k
hqk801pWRAkzZh+n3TVhdlu29EkyAiTYl2i+oe0h9CdiwtjP6e29m3RIJtGx8o91
2Xp7W9poPqTWEQjTEh+2iQ8cA2iNZlO+68TrrazAOd+nPuxi5BRfrwTOOnlmojSx
0R5qV1Y2I0s0pc8d9AI2lyD01OsnavV1XWUkJtLPQSOTfJ815+ktcf74bCTj9Pkh
zR7/hVdw6QvIYW/sVhgdzl3aDcCxzNV+Wf+OM1xOP+sZ1yJ3M59Ri5nwmtyXlQtG
JI6kgfCpy936R1bcDp9CoCF+gJhELVWq50kLHlr+ezr3dn7FwgjSP6BPGbUdkDW6
6wKEmaCQGAwEXfKRCNko14Q4tlzoxxK/xGrP3NeuYcRP6dAF1JCrmwnCwBhVFJKs
BMxgJ9RiErNaG7bQPiQsmZ3/bS7RjZRzNn9kN8qBzqylNv+HqYKT2FIHfjQnmj43
6Kq4FCXgT+SAy4L1GjEPdQC92blaZV1a8eXRC5zzYRXGFmYGxbXvpigiTRGpzBIs
r+Y7BGvHDNIh0At6E08g4OXYg7F3fnRpmDMT/2iP8Eeiv62fhOJxWdoI+Gvr5YEy
+DvlN719Qm8F1BoIB++A3633SAtj+AJ8kbweptdQKgkq5wGLRVU4iO/TlTdcfY6o
OvRMQsxl+4mDt+FkSkB8AoxFj2sfanGy9bcNOkoCKM83MgZ2ZCY9aRngVGBhMYE4
owtUpzZVE5+sDM4fseti7om3XX2b6ET0YSRpJ1bteOkJNh6WXRPTRQCE4jTM0SfG
xsw8x/OpkhXnW+sUdew0ciVHktCNab6dc9W3Ra9FpxKBpKXzW04NfqGtW7F73OHp
hnBb5Ppcch+SepdOiFyor/9c0DZ/DIezpc1M//NDjt1Tcq+4K7wNWuFHQT8+GMYc
x7WKulymeXLuwKBJq1Pbk4cKG8lS1EcZb/uZQK44IinnBWBq3Tn1Wz4DkEjJ53xV
ixiwAcjS1GkoQ1KaP/I8fZ9S+1YG9JCcB1QiHrwDP0jjGFwc96Tu3A6IrIdYV65D
ZHKyggGOdsFF3nIMw4+fzIq+4DaGbUqlr5QXUs4TtiFqz/Oy6/AZflWP2BcjR5tp
KgLoawmIBCV8Ims5BoHKqXTbwj8ya9a0BZVoyngi1crgijmPqNDbRsjqcK/QG2Te
Pdb+6WQHrV8d1l1qjJyHFV44lCH2DzqkQh8U6oWSQAAAPY9jVDaRcbVQACwgnBkl
ourE0Wf8qjZzOdAcFUPcnBn/4aGehzT3E7qx5MrKvXY=
`protect end_protected