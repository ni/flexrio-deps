`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
XKfcKMLWLY4TfubABeEmfl7dfXW1qGE/uHJ6TxR3H93dsRTaWeW2BlbFotSwZ6on
+Hxa7TZyYKFpMXvPGNH/c4GDa2einwzS9PVj3oi+Qsg6F6vTgBjeCOSo1Qnbejq6
NmXdZ7dEXsFbntusL34lq0NV3aPkcuQbYjkKIwql7/ycn1y6wdS3n+QfoZgJ6TxG
7vWCghHQfn6/yZ3qPB9cn/1OzkjymU9mP8U7ADsJ+AEuGQyJ8LWRNwfEaQkPfGay
mvrzvWb6iEj/J5YnbT06fIZxcycEHjN5xt9FapoWPLJE9LgAa/OEsXEKzSXacuiH
USCLH95OTdT6hD1xYykbTcBt+rSn7NUvtUm7PqicXUe4KLrfloJVCLcHfNVVtI+j
tch06CWVaPpoR1UZrHHZcOQZKSs+n2/hoOgS/+RIR/boo7p4z7HWrMdisCz11BSC
uZo0Wm0hicA5NNsBfjlziIgzbFB0rsA9FHJ4XLUQHFxCFGS2mZNCs4+TosplX/Pi
KPJP9T52Z8RcHKbRp6Wc/iBTzc5FxhdkscceIAQ9eVM+CAfsouBbWdrt/043N2Sj
zhVmenfHFSKcYCK6YgvVMFtt2nqHjGynKGTPPWhS1jIPhlJ2e9MqWVOUhce2wfOW
pllpfk1ikBxyPBRmFe3bE5kVZijKP4cgXZpehj2tOvP14If0kWk2Zmp3l2H7YMZK
BF6T56RjJWhWldC56UtxXVQhM5K3k8IIdxpQa5B0gd8fPUIDN671QPGpKkduCrtt
u27tX4hXpAHy8LaBfnNc/9rp50FbgKWE/lX1k0UmnWtg/agzbFyyq5j1zW8B3tDg
vIEJfFBIM/uhr6VouBeT/Dez99veVPhqh98JG89MY3o7iJHr/mxTb1Dq5CXwtYQx
t3/9FfbJB7/wqtrp853nSuPecYutkMb7gcoV4NnL9w1YTgJIKaBj1Zl0lflaUqJm
6admR2fdcNKnQA1dEikDhLKrmGxx8qotlJK/+hrGJR0QwTkfe/q5LYvOCTjUeTMf
wcQCMFVYfcaQmzSg6XHdYENsHWnizL33H5rraaU6W7LW83XCPcKnR3zFL5f8rdyX
pRDgZSNecUvmk9rAZiZPIgnVDqhwc7GU9nwRrUjUAi3picdtGimIxu8lf1WyxBLt
YZwDQSKlMdiqcCxo/JZKPCddbfhvC15+4yslKtwVG3g9CosXpeUApzDBEwDF+FOw
r3UvFHa+f2Vr499EpDfK1UTBunr1btjbhrz/MrrZcqv7MUD5WhGKzDCFbtVXWR++
rytrY75NUt8q7jEUPToQ6G3P/BAUbe8uhDeu2N9QaXWXm89vPEAJpAtjVgI3Fmi5
m0h/CrrSA9ZyNIP2OCi4qoIKKp7N+v3xc3o6gkQ8oxkUvUXpJibxBnNMStbff4Va
dPyyAOf8VnbVfxbDz1I2FGiFV3IPomDx/JetRp2oI7Md/Sk4g/UNePVi/IGXEvzV
dUpL5WYHxqI2so3k4j7AFBJkJlKr094IzqCp0S6kSmNZRuX3lOWwxzG8y5wDtHzV
1LhJDzaB8Q28ONS1Y/mO3qzX2mVFQ4ASNbWbys9OIgfV/7G2XwCy7ZfvAXxyQ4pg
0MfPxsMxV+S/K7sXn2BiFms8sB5bnJWya0LoeDMT0I41JTwl61ERV69WnmSFwClT
7UMDatOY/yOtMMDKzc3x8vU7Qq1NwDNdRPAoFC4f/44ft1VDWpw0yBHMIldFg1gx
LzYQDAnDHSf9v9oFXbtlKBht3GBOhuXiocSV8kJn9K8cnWJN0zAgaw1ajhKLYbnP
iJq0cvaubyotPxihmHNiKPumMs+8RUF7mvRapHMJq7hQYUJpNnEwiNvOLJs8bEqK
YVg8MGjRaOdSMvG14i38DRyMcm5R+FOKsWfojyGeETeniXAMEEk4QVdmT+HZQn66
jMXT/w8nYv4M13AWK0Yjt0MoIP4yVlHNmD1zDWjtFdw4cRSHZPbRnRH6F5KFG5uK
X4NeQndXVbTlAfidxEg+M9mohO/dZ3gU57nxCO5sukakX2jW7LPjtOlLAuzDfRNN
cUZmRqA4p22fkq9WNvcLXmSv/f6xlY9eIs6uiAJdglIw0h40N99RknLHHx+U/au+
1w8s/SLNAifdJUC7xkXTSFmg5fxIEWhjWlO/I31+Q5+2mTn2nLqmj79JkUa2uxtH
DWI31sj1wfSzT8j+9Ue7M6IUriFU8buvdFfTbBgA0On9yJ6hxnJyRkfAd9DXqwMf
Ryr7qfV8UKHP0H5JsD3cJl5kcqTUpsX2FAFM2xRXJn5yuIy9feuodr1LKHXg6Wwg
vPbAvZjRVdHvaear8rMB83H776i9vLhPoCMhmMr3Zl/nBbv8/d8NWwAlcen3uWBC
pqKECLUIx9JbSm5ak9Ftwlcr2a8WgVXYIyGYlbhzGgaULI6IKaH94+vnwvXxx8uZ
iiNRfu9klOa/xsrTB+mg2OGRAqWBsvJ37Pux0qMJ5m9ktGjPdCKc9k8MrkYHUSst
xq4w3jW/MUOcNKhY3SE46WEcfKvMO4iHxQby313hkz76JO09MuOc7qECBxWzJQ+W
zcMviRPrUEfJkldVNYgkoORgLnoh6FyQ5zp/EtXdWZA5GAN34s4mCzZh02SkcO09
A/bizlE/eH0L1sfYmwgxzeGsZKOs4mrPMv5b89bEV4+xDg4vwZfy/jYKbGKEuQMI
ccLeJpEQasCFIv0VjzfpmFTZxWU0PNoNYR5dgRqMIjyBuUwaFPtDGeW9Irt7SW61
4a4NCJRosrFKKLnold8azbpAV46/fPi7AK/q5AaViMonx69nQ6uPTrfziAsl3ycW
WuakzA+2zWnNZ+KDwlw9o5GW+3Q3yUNJCcdNYw4UVSBbUSlEu8C1hZo0whvwxdRd
NA0ASxRIYsYnZ0p3NGjEM5diJxVxXUvaxSHWsayOyKy516K98YeCh7zfLa4zbrs4
oBbr9TrKkNOA9DSmgxbvEJlua5dKfFsbaWfd2s7LjPsiVywGf+x5+6sCPM9lOkAd
43oRByEcYkmxyxf20bvUj7BB+c/GBUd4Kllh02PXUB67iARxP06hZ3AxXsikU07J
CrUokC3c/j/e/ATWWFnzmxeQ4i5AG8XpIGaUfwLTaC9iaDD0rqTLNni+32yMHI+S
xvPMN2MYDUoxZi/AAOD2QRrt8wbVdBW9rkEd88pM+MO75noOnrj7pD8uHlO7faEh
IUoYWwK8uuVO+9zFr/0nk+zSjguymkUdwW32hx94cR+R4p6LSMwVmE4na3koOZAm
Hsw/MP/9CPbxs0x8sSETYmVuRLAC0FwXMN5ZgTFhDFLO3Tx3RjedPSqD1inE449/
6mUpq4M8NmTTriKHYxjdbwcwLOKx5uD4PpN9QE3T387AFYLahs97BVBqgpU0Ny9R
Xo5B8HThF0izLw+qVcBqCnbqLwCAWjbP7Kd/n0BiUuuT0Sw0Jmw0BM1uYtiOFcbN
Q3/nmtIbYIP3adAlnApsVSxYWXxFRghjSqQRAm6jQT9UhHn0clepqvmi7+oyd+wV
S//AXaC+YcTh9tVSowj02lPWqdxD98A/laHRq1F6n/z4Mpmc1qcE2Ah+IlPEOFiS
fjOhcyuOHdZ4zMqsEI2va/CumFnnM+ISxEczV4A0mQsaLRBvXo4NtchHSBftlSeb
fg0iC/36xE3RQC+5mzg52SkrStbnM5cTYkBADfClno/ByO6/OwREjQDck0bDe2RY
NXptqP2lsFYwHCaA/msgvC5bWZ6OmxLKN+1IDR1VLF1Ab5ia3lqBo1ls9Az5+GCj
iMM9k2xbQAFo8XQyX21lfLHJ2mkc/XGaR1CMyV0p3WlGGrsAL3ZqodB2rM0BWmUk
W5wwY0mFlavZNg8Amd1Uq7XhUc2wK/Y1jiMRAn81Fa9ZXI0aDPP687KoimwnvHJH
za6OFFu1aG1h+Vmk+tH22UFshbiO6dRnU2JQRGQ9jguHDkIwZ4wdvN595yee10vy
CShfb4DyqYtJLrm0GarQjvPydCq17EBMnRRqHUHqRobvnEQiubL7WHFBDMBB0y/H
knGCPXb6Lwqxi3DTGEwsjTIU39fbplbuSrnMtmJU5mQG9ZlD0iV7ZZYLHf4LYNOx
HHv0xC41mDdhVIfYaTBy271Z083wJCReJakh+xli4dJjbTZO+k+t3k8Ceqiuirh4
PLU9vkSiNEJGmJdGCK5PJfWu9V323f/MDTZYYkQ0FHGG7RQT0pWX29U4Aa70jy3e
HhG2rp0oOZpJlqJnQ01WXsTRq8ZxaxgshANwJNQC/5upIigZfQJVoJFSOQg9NEaQ
0OC/2PGHaSnP0AvQ14AQyFOYvQt5hZVpwUAxb4ZXkqsY2A85J7KhbAqL2HltC7y/
/vNLCS2lJ+r0gBuEyfJhrpVUYDM3JCPY4MK43zhKi6xPaq/EVjdKBjBfMNVcxSxa
utJeW3k+Rx+QBaT11ImlR+rm56esEK4XbO7rVkDMtejMYwyKLnl7ZL9IyFzsa20v
F9nRcvv8XcYvf4lkRHZ4CKVbdUM4OTSQfHGBlW3HXB+LVYMnzsAB5XZip0JPBC2x
BznIA9fbjoxCV6qs0Jk+ZRNoyNgf8jnFrwZLH+oJjlLml2Fbk4IE1jR4YLbvVBjH
gM5U+Ju65Ge3DV2sOHqv6zmwT1oyodbrjbK7urXBuXiLduhpvo3wqEci6JlLgow+
priJJmsny5dcmQ/w9gFH41BAbPcwEREn5SqbXpKKg5ANQVpQo3fcb33x1hOUrmeP
CvBYwgnM0ZPho7aMA6A2mzNkEshOkgfOp0M0AEgLa8wc7GBAqpr8ybocBzoASnL0
6czVdpKPQ0olReEvPrxEw7SgnD29cDMGZFY6XiZXQMrss1/X7j1XRlZa10inM1lV
9tsPM1VVfdltGYVhwE5ogbieR8spaWO4tjzJ4Ce5hIq7FpPI6jRqDEZxc/iQEF6e
9QHa6lXzy7qY5uD5TzWSaiBOnQyWRPmvwFmgXqCoMgexLQ0VMOhFSInjWiuwzS8g
ecnl1+HJi50Zvd7kQqw/TNUUFygBgc6dCDZ7ExnzNSRWJ1Ve3IQkPQVJmYGbGLYL
kulbOG/yVLnup5YDjnnTIV7LKsIBgn/seb8y8j7vql2tK8bpBZEChmK/YRBGNS8p
L6ElP4cqdOM6uuGGTZ/XZKx8mwM+sPNp38IyKHCvCt5jCTvtH1xjDA3MtAiMsLKb
Ioe7livYtHpZQYGXUxbozGtM05UVoI5/dkpPmMJIZRNNl8JRaWr3fT7NUDAQBYZv
8hU7HovA9kxFYVMCT07jTPjzFZLXvHA+maASeqe2unaBknlQ3d1IPzwm+l/WgXrf
aLwI4iwdkCyNsy+W+gTuNaHeDtMHR3YrRLVlU9d0aAsaudxo4MyjLH2oC0SmknWV
/RchvsNjnOSUNXvQEAiykDCeu7qNFpKE0QWGfn7NfSg4tcw4hnaD/0JPjdObjzxQ
J2r1MGX4wUZ2UK64GjCvQwYraIRafqN3J8FIVjzzXLwnBnUYyJOpuSKY4ijbUvou
/JCr5hfBx8XhUVDH/RXZp6b53buTAUDqcQyLIHJ3K8fZTqOIKw8mHUUuj+eCqgsh
CIzNum4NTxz33ov4vMPIisTvBeq5oMYGzjjNI9HHgb1GTzYsp4GOVU2urMUkqBrF
q90F3F2i0u2KkTE7v3fs80AR51/F5wVLtq5LKZZ/vqvgrZkG8Sb6jugXmbzOdugS
7Vbe7xlMsZSpkC8QcwNTAQgz2zI0XG49Fa+SYdQMOh2gHBl4EiMep5UhBQIi8eWY
r3usucTFK2uJfE+oLDQqRdZt+6A+ZpgftTKNkwfPO0Zo6FBQ1Np+hntkvxnPH6ak
IKn6wgqwY000kh4dcFL7u68s5lUYvAD8zmOnfGxHSOK0L9AMZ5mB8mEBveKepAi6
+D6l6IUl0u4L9U7L4FelDTtQdv6YuEN3McMwBUfOk/jDQZBEQ+jHc4Ij2mR4M/H7
SlskgjcLpXBAcETLD/L+dkQZrHGO0VqWiJnxErBntDGBLcgspKkMXxE6+Lt9Ouyy
0wC5cYgYfOoCMz/HpLLZCDUL8VF4w3jmRmBEJuGTKG5Sg7kANrnXMm2BqqO0HzAE
9ufH4rAjqWU6BVp3f1HdqsSfCXOVAluWBF+wmE8TdgtO4l1sm8QgC52Qih1WkOB6
CeQYgAg33PjjplPpK6QDEk+EGGvHYbbDBtr+mkCgWkM4vWzP/frujBFHDyX5bGBs
HBaWVRtsiMZWpb9QUE9q/0t5BnCk3A/OCP55zWWRJNCrSi5GDLTwfUEaNCX7GY3p
fmjjYmuHXeyjKK3fVi9KZThGmTMRTPEPDfyJs+vkXAL4D5BTR3Xa4I4OzqaWnDO7
rg0dnBycBNYonk6wuaFnKuz51v8Td4NIfUcRT9dv7DQMeDYpYw0YRQx+zfyeUQWK
PdaXiHt7uCT/EiaDTkN6CulMEkxhsDtfpBd16LJ/g1sfv229aURP/BMkAYTTCX79
2q2TY0529MUWxAG+CLAk2zQZeDZvLVO9LaRvudPcrgQqBtVuyio9zXtz+w5nEYTK
pwnhMsba8GFZ8F0jo5bjD8pMek1dNtSYPrkCVgy7YGtFnAPEqi0MoE/+Oqy42pAh
sBVyQZd47RukOC48mfLISl92O1PO/LqByQt88i5H0ZJl/0WFj5cJ6s3ZZr8TMQ/p
/0uAeqmbazw2t9mXNLWJWBGmu+9qZ/0cw2Yl6fK38t9AN61RH9ggWzyxWmewT/ZE
ZMDfQGGSLLWwniKzLqOUaPGpG+8sAWxqif2+YvWHeK+lszdwB6BQV2b1qy6ov6Kw
7PxKf/vWudw5qbkU/HdFhVSVy/U6lqOj7AxNZiePjwQMP54hnYtHbJmr4SHvPdNB
0XZ3v0gpVumr2PDAapSTdPHSiLmHZ+FZ6c3sy8Ha5cL8qEK5ALgtjOjIMVONqmRV
LOWBASpk2M1FC8V6fD3XII3dKjTE8wB9vwX6M7D/101AeD2PtTbi/adoWFTDJNi4
2MxF2TVIIAq1gVl/Pofwp+IaqyJ2up1k2EG897sxMof3gAa5ttQbdT2ID6iJhQNs
FD7dpQoLfK5T8109sZfIkTFlkSKuh2PiekxYDt/ESEE=
`protect end_protected