`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
pZPBKDWpw8SI9CeQ0UEeIYiIsHsG9LgtnSh3yulg1qEcW9s1wYXDLmQy4FxEL6Tn
7nmfDWiHeuLZrUt2HR4En1FUtkufI7v+TKmjOYmuxBJ6gWZLrvBv+huKu1M7yPs7
zMqdfONibYpU53t8YWLD9j7uB35jSVD8Krn1E9wepBdHgm7uomy9KEQxNZc83ITY
fvjzVqLgqdUrXzt9/6aAJ0ScX2KE149j44Wxya+51qPWbqYWIOH4KI2wnJ4ua+mm
h9T7Xj6oVYbhMjg+TZIOINNy1rOg8BI9M6wNMuU/J7+YiNAy8uFVFQzeEvWSNytI
WF7AD7gwQrWggt8EQbObwKU3sFO0MLwndhtspHX3R530JD4YkBLPJuuF9/JomwRC
5UU9BHtrEC374ywBbr1jeCeC4Wgs3+xHIM+mK3uw1goAu42lw3D2YezbloQRZiTQ
LzrIKRG2029hK+xgvZo81vg08dbmSljFRh4dK8lMBAP8MVdz5vUPRosT0yKDzJRu
uX1HK371BgY5rbNIFwe9rGYjefFU/lGrBGLo0U9kRhuqIEkQCI+DxJWZRlmpXx0v
vxeyMmT1rSzWZr3+EJdVUFfgsamBupDxUw9THd6bJUi9jCH55ozbd/2T2HSVh2hx
MKO5MrWNKqesjATR33Eqk6TYTFkgNxd56TgxnELKxhGo4oyJ47xb/J5Q5BdMmZ71
CbSgiNDFKf9ia26adSJbjlla6Q9Ujv346twXSk9LN/QRBeOExii7L7GtQMZydhnM
fceQZMcKO8/Ja6OJx4P7o5tr6361y69B9U3WjBjdh87LSbGlWuJ8coynEdy6s2Vu
AOPAXcLGhs9x9ENMt6cPIApYxaDFuSXC1HCh4xjdeZkFJj1tvzJ6OuElSXWvGsnU
MLXAYCkICQD+M5AVtC+o32Rpu9uCNTH1KVxxdZeOPJ6cJ455pYXaBif9g/t7fGzu
oLm+rMhOlPgIiRTJ8QreRmUHnAXeffrkOqntDEp+gU9V6TgJbus0xfNkGyndethU
SKyjufxjriWqsj4IpjNnV06C56AOci5pHbXOvc0Z+Qi0mnL2fOKzhJk7jlcvZgpV
p4cqyIdG+H1flzJg/CFbk5YF1UWwtfnn4XUgVBVQXTKBD6YYbWY0VfXV91XCqjq+
wTmxgCLyZ8waLJF/UksQe9Uc2ff28RsExVlDrXZ++5ZDA2Qmf5hUU+nuw/apc7Jp
1gzSF9c3C6wBRmCBEvPstLZyEPlYGV1rrm+D0cg/770kMkospW3kkKAKounxbnBk
3pLtQNh0eX0PBb8y7dI7CevVPhUxcr2+lQ9iAuzpbyF8ssxAuXMdOnHLDheeaArO
R2uxmXH28a1NWOcLqDObTuRBQMWyzqPH+W8lMo5KAhTuq29pY3KdIJyeuR5kvC3r
IO994rDdHb2L0l6H3imUxeHAz/dKtj7fdJJAc+zia2nAimttfjyE+O8gQyKtuRoW
US88YDbIGRrAxEMQKv0KJIwH9S5wyjv0ZidJwESzfoAc6Q1JPL1JjZsm1wN0yv0S
HdbO7wcYRLa5i5e4QBDDwef5/U5wwg5kP4B5FH3tKGZS1u/Zk9kgaaBwws9AEsKO
OILCR99QEEpTET1O5yeM14WsDb6nVl9JdLEnWULAZTmvygEHBT+m5XUk5trKUYkW
2GC7mqurSOFwfAnUXB6FypGdg3EhqetHtqNaEd4XMJ1qTLZ6XnfJkxcqnoUQaG2f
iDXF49bc7auZirFGcLq0Ss90f8assl4LWPDW5As469xwt8CmoWtRVbIVHJR43fXE
+FrgutvezSzFTeyq73bTKRwsCf/Cg68DXIYxwdRj2Dpo/6eMquybPy1RKMnJ8MWV
WDRdqdbJX4lwgsD3KaRn7CuId6xbhMc3ZBfm5Oy/8qH0CvYk/M/EBNLPaegmm7Iy
JycF7Wrt9uzP/CvockL/UmmfeXEasVOj4IUxR4+fuVFYwiIIT5nkb3itwKo0K/8o
dbIp9BoFq9I2OBgx1ksUAdrTYtYMzyO+WdLMYR+GvW+q40kuI9uWcIHV29GhbgcY
WYxO5IAArbvY8Xp4A7Oi+IYwmKW4F1lHbVlX7b9zpwISyQLE9uZc0F6QDsCof7cT
kGsdI28u6ebe+NJ0lzfIL9uC8tCG+pRzZ95oq14CPneDqCTi+qwLnrV5njK1uou0
qJeoWmCvn+NasrLStT2Ndj7sDnFQTZ0eVj+7tFDbPkx4+Zi2+Uku3nE0jbpSiiLa
ELtGgQoktcPgy8/Mxu3c8O0OLc8CW4pxKuxsUq7HZGPJQB8/XLWh0scBqqjNmnpo
G61EzJ3szFjZFrYZAxt0k5o1TMa7elZ2vEAcEHDRwvx6eknGh7hH+QZlhm35gnWf
NYOL0eEcLivecAu7krZNnoBAD9lXicOeG+xHO8fKMpekCtT0HuEGQEUxud4s5zVc
ciS8nHHqSF9MIh2SEgu1Am3py48g7NwVo1X/IPrCmjqMcCv+8sZQLSkti30SlLDS
osQb7fyViaVVs/HOa8h2PP9Gyglrcgb89hfwVQLop9P2KBZQHjxvL5WYZ8PWs81r
dJpXmjdJNMpORW8Y9N8u6+QkXzCLP8NvRMI0pseKUAq7/FtpYc0t2UKhq4xCiTiQ
UHNC/hiGIPWhthYfeU8fpMJPh3V9zJSg8ns/sDbSquqiCQoLYO8qNOruFXiUiI7B
eZSOijdqH/NJboSA24GdfdFqe1BeDQoUlrTQLScSS+fLzE2kg6CpRy3Mr8sGVYOY
mkhuQi92FwWLg/wVKXo6eMoFN2cu9ikQWdbEbX7Ve4AacR5fFBSaudCTnOGLs5Hx
0vZXd9bZjJT6tZC4sbtrZrr8psFPhulE8sqRLtE07xqANIrKfKA3phzwDFeuQXFi
0sZHwSvSRQZ1KSiBUjaj/EKEujh/+V1flWfdw7Kbyv5p1zgNqy+UylLIRcL+S0t3
p17CoHQ6I5BKrV4xp+zQDE6GG9T6Rf/oUNN60d0rPC9U7hxRj/RzAjLUFu7whp/k
uyq4vhB41WxFphX0w42k7lP+nqW75CFYXciq3CNbWwTSZmTb4GOD8uI7SOnV6+BI
wH8oxOdiiltBT2RwvXQUBsuw7CmU9qRQ/U1HrrfFiuKN6q0eIEALBUfaYQEQCpOO
UWmcqva2ZEhT/Rw10SYLHlB6CJvSttyIqutMqdh6fXsD4mQHEjF4JlcqjtjkFXlQ
EqAb/QQtkaKEYWCMSXaHGtux8aCw0ai4wNG3uClcV4PL2R0mo6OF99t4MM6UEFVi
P4BA8ET2TEt7reFqq9hOHcx7qd+2mGXmHNqOTvOq+RyP/WZ/1AbCLDMyrnnTYg0y
Pj152W6X12Ipf+KJ7Rt2JEH81oIzQsc/fvbkty2HENnGi1oC2xhP4EVmgTt/g2Za
2JKVRiHPOf4wxbU7bA6qRgiPctjFAwrm50SfzjCHrakjTj6Y8pn/+BQYoybiHOc2
0B/lTkxt9JUQY2h5vDy3lKrE/DDROUYcXWQmfiswaFdQDW5mWofbF0roA4ZYtUpq
vfSU4Na7FVfUfEewMTRzVPiahljpKqKiQxdUL1mquE0iP7tMnavMNre9FpZ2rThe
kZxwxy43LfUxIL7vMDJOX2k7fEcRKDHYb+Ka1b2JAtdHe8RrvMFjJvT5NdeMqzOa
h9inGyiRtL4ymMRYZkRmeeceIJB+PzRQrLLdjoYJoqexJl7UIX9IG+764eUEPp1W
kWBH4u75dMaWvh82qFYG7HS9w+kSpckbf0YWLifxlkSFfcNJF2RouQ9VMNuWaW3Y
9XTmI/kexGZd3u1upYcwWZKII62lCGr7rYnwdIhLWygJVWbtlUelQyuJMlkfUPz3
YmOz5XmQwY120CCaaoaMK88IAZdDM6uZ+5dl6JCy/tXAU5XLHwJ33RXDoHrMUVay
JDN9rrmne9DkVLrK2m6Ay+yI4i9snkn9Awn62SK1Gj+yCpipZB6ZFynGm3O/6mMK
kh85MFilH7eUP81t0zLRZlx8nbGCRwDv68FU2dzcA08Ef+PHaxk9wFGfYmkERAfw
5vWEUaGFP4HolnjsGbKsxulpiv70GcVQNv/FU2hSwcQM9b3hMKZGiOIKaPXVPRk5
0Gcko5xxo4yIKA7WNGdHMcnD0XzBhkP2bzaUSSD08PHA4VwrdAUAmWRPp5Lr9ldc
ioXd9tNGBQ8bNFq9lN/wHRaaA9qimkh3af4qR/JjUmHXBuvMwgeqN8coqhbX63dy
c4F6rr7bPTrO9AA/8Lm+EnCnfTF5BIu9hhukb4hE8oFFplwCQNIT3AqT1VbSXi++
/2Vt03BuNGHdLxvrngLWbgFPO/aoserxJ1B8BiPCCFoRwtblX7gtsx7HMa5Y021g
9Bv1O39I2IQNKFIw7yt8+CpymNHcbpzpr3A0kY/PAf6vEX06xG1LcL+dkI1AXea/
9Z888dwtbmCXhJRUi80u52d9awrag8vMZeB57g+OSdMaHAcx+8GNLKI1SOpnVVSD
qqAdaGSaovJWBujbAnDDZULSaBgoT8DxiiAgnbTvVgBGly5AbC571Jjf4cfQRYKH
P4sOcqfiohog/hcPeWGecJu0fPmSKT9DswgJO2K9727KjmZd/2YkgV5FMdPG7OK9
MDYUw5+KB+KqLWvCsrp8PzSrMVEEVWKmW2o3X9kpB00/iYgPWKMBTHoBSDEAL6L0
nutOfuH3Jbnbla405bHhv2fL8jQ+/YmOuu7hzeKdvPpf8bGhFNp6sIKNzdryCGG4
GHFDs8ztUUlCzHnNJBi+K9sbkrIoUbfcm5M1xZqP42ib13cv02Cg53pCTmqpTfSs
zfTWSZ3sXQaW/S5cAxsCcxA7NYTA1F850WnxWa00ZvoGK5/Hz3qOAsOwy3OFWthJ
cgFGfStfU9hyaWeelPyvMWPJ7PD+Pcp0OXyorUOYA26OR9zpqlzmCY8iuEs8sjVL
4OlBsVFeDNAaILUKBDi2GtG/PB+9c7wSYjzuGtLcabVP0WkFsUdK7IzHizASA7R5
8NRdmnUk1Wkz87M25mDgMRs7BGRSrLvIv2lBQVgvwLyhPi8+mG4avgXQAQNtkZv7
ZW9n+1vFP4lTdAv8WMYdBbHAErEYHM87icigHrLbu2eNTwYoDRCYYhEcTGcDOWUj
X0bwTI03CFvjfniwBG+BXrMVGDUQ2jOs0V+PAaCuh5msDWgjCQKQN7YL7usoM1lG
eJ9YfZrznQgqw5etyVaETHDkWmifkbgOAhuk+SNm71R0SQbaFF/5DUG/okvtMNlc
gf89NcL8vNM0dPpUDrAFya2pLbQbVxXVYBmMgVqsbiAvbigrIjK94jYXkJTxa/7y
u+XFV9CzSBuABS5LHlWGtjbOZDq9ZbRW682YRg9y4umrIFY5vWPUzYEHjEdV4mJC
cjkq6GC6LQ1WOxsdZPVnoyeaZxeBPcyqGBA4mKJBjTxxqemeUybASxTdwXGv7JVU
np2SGgZiQlHd4LLsKd6ECx5pcvz2E87ioOSjeYEHY/V8tRV7usprdpyL9b25Ti5C
eQE0xM6KcdSBVbWF8+Qwd7KYKQChKffFI4gsm5fUu9zMPCzLbuJQahPMpa/GdKjI
r2XQXR9i97WVQKq8Ydn9yCjO+a1kO7oeMleaHOi8gL4sSyqvuIXZS2VIw3W3vXg1
J4yWKfY35WZP229C7LdohgKIhz8PlL51p/AfRutx3Wf8CnIU22MdD4wER1jC9MdH
ccS6qKMDD903PlxtZWGxINnug98QIHZajbfjkVYF1bEpu+P9YIfGF2VJ1xyoDjQJ
nneLjOs2xjh56R1F/bNYYMGaHO+AQwsK213AyfmKK+qo5QO47yqUma3pPC/4bcEI
tw3tXfl9zhYYJLVLOzLg2vsVWfwuI0Cito4ZJwx2i/KfnPLmf1S0pkJR4iA9LlwQ
8WGqbg9ccT0OvX9t6cuWndVgR8sfPMl+asniD9K1mAUFO33HsxiVlBTQRdrc26QM
ucxYvqu44hIo1edhyTM6V3RRjehACjqB87SjqivCU12r6ZVaNbaIqeT51hbaKWds
V4QpS+rpfq5uLshaa0bB/q7RM9B6lE9zukhdeeGU1XBH7rQHQo4hp1A0OuZ3Tt9d
ejKkwJkVaJGYmL72+Pyu5lmoSwE8DdqE0ef9LrvaSZ6+u1DnK95JTtb+HH53PDzm
VHOwh22B96X6e/+jW6VduaLvbg2xD6jwdbAlfIl1AA8gh9SILnqS5eUSTQz2O5tV
rjjYCm2tFHfbQJFoFkAcTBWpdxTf/cHCGR3hhOm9mUKiNQdse/v5S9Uzl3R9vs3Q
Lt0aKVhaltwtAM5MyEZSF04EBHsO3m49ye/bjgdBKvndCzbjrkG6qSgSZSnIRp3g
k9lKV571wjt63NHXJD4yr3qYSwgMt8xg84ImexEFbkrqcP3adP/SG7d+xfOuRAhs
ubv7c4y4LdTnIDZG9BRWI/UK4VyK76rdKu7M4s5+0ODWklQ1HevWRfpwpiMYxjkS
AALj4iyJBsXRzXJ56ss17qBsVpHk6lLRJXq61JKlWgFlAT+F5/BshRJc5Tpr+6qG
1xwaX5wnrsHeJn8D4+u2FZrVpGCkQC8D3jRitJoUGT4ugPACIo4UCvg3+QOisQPT
KtqVhQXR+nOC/HHMtoZXUcNrh0uB9jlMTO4JHcrM3+0L2hdg90onXUqAATmQ5Hcq
+q4I11eX9Lq0dTEya1JybO58yrvbRiJXMJfMkiCo99cXOgqqbEshkZtkrCxIycSl
2BbFQntvocn3ATVkDfjPWOGUYRS0oSc2IvDrvL+mDHsvCeMUdb2j+08GPOHfHkRF
7dBN3ZudTlb4kqM3OeW5dWYhsB7p3oIwJgMQq7JSzu6XPkCCM2UhUDeXZjjInHrX
7CnsYpiaLFtLR1LVrsj/p5vcrPmbej+V1SItJ1A3My6MXNRytc4DKoW5h+yTuRF6
0xGY7bZZrf6YbC38U6g4cn8Yp51NzXkAbEhxX/yz8XsBk/nv7NN1LKK7J5Caz9GJ
+m4Asd41kFiGwD8Vh12zaJ1Ei1xaZDaMO/hqIHNtL3oLlbuKK7RIxZFIzOeDuu4U
kB4B0Q8NWc0MVYn/Wy25cDzf3tQg0I1R+X3ulBHR6yVXge1XiVM6QKRNotIrU4VI
HrGO7Q8jIaJVOmq0tW0kBIJ5XVgCd8c4uUcTmeGGzxx9v8zXQ2xoDjwi4N+Hc8pv
tKkf2Zv9JxusTMNUmkyOsO6fS+iwCUSq6v+rrvZbZoO+PVVvrDhXa3K2K9V9PLC0
AjWUUXtw3fsGiJOZHvkj9YmQBOQIQdls7mTctg0ovNcPxi9IKn+zcKgkKUFoXKu3
kjlBIu5z7xBhwJqM5GRlnaFaSDB/VCWxdapbzNppExx4sqp7VFDzCTUMi3Rf9Zt4
hWEShdhW/6eQxXivvv4ZMrFidlMigkqpRgWhcvdJlKwiATPUmHB8F+hLL1+sujdP
EKWoI/K+weblmzlyREQ2PPUKdL3MVuZEBShTQBAnN9Xh31gGPUcRVIsILo1SoY9M
jgzdzdoGitzS1KMSMgTGzT9g0O6Kxg8SzetyARipKMAg0bb819eDVBG25/HMNEWl
9mqoS3CJOvbOXdDRc1Ax6e7qaTzvDS42ku3iOnAtNgK5/9NfplzISFjrp5qQIyJo
qapKWp/S+EmfxZXHE1CKJq8+5nccGl6DWhWfz7AOjYVxr7M87I+oFArrQ8GAfUYL
V85b7LnOLIcbmLQLIaNm37HCzhSq7+9UAVMLo6VmMJokBOHK5XkbBhrVWKubvWfA
oZK/MdhwVfj9YVdHWiil+QKUdDmmg8JdGVnDO0IKiYVOaey4vQeqbgb9CNThGGs2
7BrBJvpQ4DRFjotbgS7b4Pxe/BleF/BDBy8Q3gXUH/NjI0GzKlTgmKrgY7K60CTj
QuEAAfKL64FV+9muBX1ITEnUgs3nnK9ny6g+YITZOHSjwsEs9vWaZwLCjSQapg04
a30iGQAhdNqjsuENpPWSBvxZTdAdRThVdu6OoWhtLqGcmTmI6APfHH+y8MGrUGqJ
JG/uw4z2mdCYZ3ElbquyYpwKIcokhJ0VyaDR/2ZmGCxch8PtZR8uXxpJ1KdN7AJt
MdyQHpo3Kk9xyQsLmM4XVOUFFU8CAMfO0msg1RGWNglGBhHFDCvqK6e8LRC9vwZx
VrfSV5S/5Mt7jAdzNVGbak55HYVpONVBNGA8T5i0kaGTjQA+KPQbPn1BgqEstoMx
3oqoBTIITb5wBXOODj/l/KiO8bOujg1THbHLJNrjhjX6sszBsxNwLYb2lw6KW9Cv
6iiOhuYjXQnyns363mDjEqJwpV7EJpS6AD5Y1ZlwszrdfmzEhlWbqlUCLbBERix2
62yw5UbyMx6N33k1XZeKShD1JgeCJL7pDfTQxZnayNgjJh2Ntzav3K4x/2I4Uqdp
0M9j42RblvbhA4P/Pyuzo3VDPSEyZ3/4U1I6Qog3BpboZgQR1XTnar5o6kKBM2Rc
1MmX/hD9M9h06aQdVabtrnSXQXS4f1DdJ2Cmuew3ypHSNpfHuxJGKoXBNFqXm1/K
d+gZcNtPsrH8aPZNtS5cQhbJZAGS4yp+Mwg+oYrLlonsergJzGSYSG98JjVIy1Os
a+AaD06zdiYPYThHrt8RueTjdZCx14oTOSLyUrF0/S5BYa5/A4RND/8GCyRbC3A9
SLV+2m+x50TbdXQTdiEHpnaBAhGjKIqCrAG5U8AP8oC/Zkkb+p/1e3r/bXo7oZJC
INnB4ew1eTBaImKnFta1EeLeC0Z93MNkYRHm/EC20k3sYClsypJU+LYY6S/i97qA
hNUySgaHUnqh2iTwEGNPXMZelJAW+EFHefvaFNCBr76+GvRzqn8Ff1DMgKfIvnWI
QIGUfDV03L2kwfWlvRASeNNk9RPFl6QoEIV3tzsxDmKjBoTRtfDdJUvKGXDtCls9
eqcEc0JEfRqkQXR2LNlJ+yZV3E4f6705WlVhZQNEheCkXpzgKIcN2p6eD378lFDf
4Mpbwu9/mvI050oB9UdDIyM0OxAoUKxZGoNL8mROLZhhLY+oGEZLvR7Mrn3Vy0ZD
RagI/+aVU/p/EVP/WXfZoAAEeGh5e5aSQzn7FnGQD4Jlay7POXLSJT7Fr7so6+h6
21BOWAQfkWjipJRGSXUT7IAJMQQQjzcnh4tL2G6SB+32C+Jk6DVLW9pN2IWDzOZW
288JAyHw5RE6b6R1hJZJqsyI/dHQd8e2RHdGU5lreKjH6d9yzQozwmRIq5qwGxJW
fioCP2TxUyQmtsaXHrhGZCg12DAzOIpujcxQnSsuKPyzNRW0HLsjjuJEo1fMXsoy
uuo1Mf7XPbM14PiP1VCFdVZREreENPxXKSTV4z2F+uX3PR6b0cAgOw4aFEaNFS3M
aJTXX32ZhrU0LkMU8BS92IzbkVvzS7p7DVzKU3khsRzGoIJyqUZAydj7AOaxN0vK
9LTFzqBBN+ogLcERBXDdLWb84OQXOJer85LKaWShF3lOhr/t475Q1RJFF03M9nlN
LX3fUz7NqJ2fi8i5pxglxsjPg+MQUlU+3mWP56fFc3wu3mT71xwt9o4jkNgt/lYE
IzfyZ7D/O/ei2LaM9YHmgEDRRsZCGUiwDk3VYvB9woWmzoNE1Bhg0WTdwo2lyrxw
OCCRJy0yK9LpZUshrBnBuWuT2XszTNCyKastolGFZZnRHIjBKhj9p5iL2EYDae2G
2mvCNl5U5UiGnh8DpT8gKFGT29JvFUaIH/xb/91VIIQo+9dvYBskiczxfctYC4vj
S2wgZQjBIRL/6KWrRN2LHhJL7HmVS6ej+R+FlptYJqeKV+xazYxefz4NMbrgDGzd
KdBXJTcWUSDn9No/QU0WjqX+XKlumhU6KjuPbK6mzsz0B3cPXOQzY9fyVjhDkBVp
In/MlIMT/VV+Ofa0ux/sjywZswgrWWf+B511BBr3Nhtq5i66IomIYHScD2l59V2G
+zi03R40njL/sltQRKDrwgCs3KxN5UEvdBTyqnCFQlkG6RuUwQKfL5vrorDrVsSx
T4ull6K8U8nJIjk51j8cP+gipjmn56NZ0DEn0BdKFxHoOengAhgazDZZZUZVaDgt
0AQpl98+V1X0BsujX2UXDLR2ameD13ZwcM57u2NTFaRoxFAaFTbom1c2j7xrs+xj
IMuUP6JOnHtxF6MIBRwicnaEtN6gLDSlFicVsyHzLZSw6zhn/pgRBW48LoOvFZz/
eARs/rXV3AZ5l3Iio2VTsBdjlMKUOWGmuaVaxgawXGsQLQVx+/61Tu15d6xoTQLC
JitujTVdyvjvx9EOCuuxYLcxPcCHSropQUnNKLuLsk4nrrz8cUYojfJSfEMQv2pU
IPGgs8DsZILtDKnSN60pmmFoT/g98NnEko4nCISbtKz2cxPoJfPJpbORGCfPNsPi
jlaU8FbsvSVRve+wLLk9JIg0PQXFfqFpm7lF9rgwm+OeaHdCVNhnh1fRAhcoKghJ
g1mDt52A3wlyOb6nNeIFz4gOJK8ri9bCMsz73OIk2smJWlBz9fZSNp8qmM4bJ7Dv
mtqDBKZ5eQhkRHdp1hpFFQTD5lfA/vNK5Nmu+fyKWEqwzx1JDPmYPVuReUXdCPGG
wxSQoP6UtFwlRMpwVohczDkYjRhAnfBE/6Jfk7u0cmc2NMveEkJQZvYd5eCzhSz/
KZPAMA7+m0G6R+EhZeTcrDh7Chq6FT4oJDV5rD0exwXlNnTv+lMnxM0s52ni54Ti
cMycWoxnU85gmS5e/2nqT+EZeTdV1w3mpVHsRGtJuIYv/2Ge1WV3jXxzgxN6xhXW
qZB/PL3lRdbrfY6hEtXwuSAtd1LUZD8Kb7nkzsNqEk0wBZ21QjFqRt/B+T5xJQ3T
cYm8hw8wigxxmmrU8fwyqQvelCCRPVJhMJvI3o8sErygaKQBeL0+o40TwG5Wuglc
NvK5Yt4uM+MjOPApl5dWC7VZKsqLbixZybl20iUXViEv+hCI3Dz8bcVOMHyZRxV2
UUdbpos5gRlIJ2IFUX0MjD1hTGoTadveHq8SAgwrTjnfg9jFdN699R5o9vKtvzRJ
NQiDAQs5YixPDZ7ikA2W6JtBa4V4JMYuZKgD6S4MBvQhTkLw32TDsy6ocOEFGGGV
5HbNNmAjnwWf3AJJu1d2S2VH+SAS9ZTXOatbQPN6D9//UAhgHQ2sod6/dNjJ/Bym
uO4lV74HggPE5yi9ov8rMyXad4J5JF3ZNhcLq+AxTYQD3Toe63Ow5xF8ny6loOda
G0WiCtBYgWy3ueQT5TETbv5UEess/onPuw/kT5nFZ1rwz6Qw0ZssqHiDxm4W691+
9sNKOHECjmpBeMRmriw+SsOmew7CBi+m9VQB+a5FcQd87EzdRuq7sCzGqwWHe0E9
DPwysRQFJkKj/7pgpeCj/DssdPRDS9otLoeACyVRmMQsBC2e8UsIj0YuBTGvpECi
qZ8ZePz0A+2L+DxXM44+gxlJQG2dSddCVEvjqbNLkf+8HbNzdf0WUL0IpCt5nE+2
EAzrgLBXVNtutrKs3oOo2ykD0dvSYIZAzrdIJwkqjJoFlULUydDVQ43UDo/EnYs4
H7sQ1JZ2TDVb2isSjZ2Gv3ZvcMPNqYc1JdOGV823drDgI1O5fMR1SELyytiTVAGu
NMWKhv4IF7TWRrgP8WrWqLVEOxWRxXxpNlLMqhiSWC3OLxwlXxDyU3rJeN0u7ZWx
OfMTgEqLpddcZO3D5Du0f2rODilFahUUXTapcPExlE6q5J2Ofc53osDRe59wttlS
LIZ1XP2t5nTFVPfLd99lafq8+cFeVSiSTR64IIndeVCJpDW+rTU21rCfYONsaLUV
a8b+zMbVjAo6+vf6eGoOcXfWv0CtRrELpyYElEIAHu5TNnMBrrHbO2rzvHtZty66
f1q8OlVBEyXl9F4lO5YozPnu7/0QN1I9nvLe3/twn8WvVZSXfssOchP+V9y+gett
fy1fy6qOV8q3KXe9alSahoHLR2FaJh2WN0B45FP+jiXe7AKts7SdAe9M98+HrumG
E7E/lijxHvW+1yQ1PcYeJjbyrWvqAbTW9UL853gtjuiv8POulgL6aTVj676fwzJR
+7QnhBurp63SuwThG7HzyZESWXjvu5PYSBiCLQhO0HzeQ2wbOMWQ6D4mPLR9s7UQ
PjW+UrCt928kNqMuh/N9Bulvwp4wDYT8Qass76kzCyM3DM7WBeitDSq067ofZkzS
FB6O03FblvalETVFcfzoBbjHV2qGBZ3u959D4I2QF0Snx9LeGP7ABKM0nha2dW8D
SlcSI0SGwoNqbRuo38fl6b6e1CV9fz4kK2qDDzifzTEvXgiQyJIwayL6WpGYRU+/
SKLoorX6CXQXuRp8fNV67jOAFLDAYJOp2QkI5e52E/aPTfT/2up7iEGweoTTfAEt
SpnWFcC96LnwrAhSwWR47M4qur+wQ6zcmSLSoGKUuFgVpkpBu5UsHXgfb9r8x5QU
nKgMmv6JTlcbErOICcSXaiDzm0y5IBKZM+mxcEx3RgFPnXWtBkH+zZIhxTFYqXKz
TqQCVEsFCsZgA5/zSqyebLI4KxZd4EiiHufyAqrJvZBYUBctKPdyUB/5lfIxO9fd
0nX3r0sx79Jph5UB28FnAWesNEb60/HL7Z4WuC7HRFkw2RX0JxXHRXEruYfglT57
mb44fm3+gAe7UaT6B9dSCaMpVgjXMW9dajbuVjDh5TSv6ucbDDwFfC2T8GNHBCyJ
Zimr1vYrLoSCeC6RJJX18wQcYJ0vSMcCZrlO8YHycq7j+VGa2pN9iMXT3o3IEvbo
/xPwi9C9J0ENsNB3Wi4IFtc99T+E8erdJcgrPFXhdDd1Ayv+lBaw/RiNMJq6/CfN
PK96Oji62+6D1O1eIYk+3gDdtOl+V2ZHW9zXNx53pPaGR1qZvyvrPSULneARneFN
WRJbz//a/o9ejRwY2GkOTxVWrbiNp6j+owGKqLPfpx36B1gSkYNLiPqKpcOINXev
Jys/ULyYQLKA4U8/9gMuOzBmR5jfFrbXl+fQYQotP1nF+xgFjtQ/vNV5Ob6S2r2H
XWP+22+xwVw7Y9TGe3sgPzJhzmw0HLcCiyU/4gjiOnH9VXe2M0Jxby9W4oef0uvM
CXAhWfWYt5/7Al/6/qJ6r8poYc4Y6ju2fznY8oOZLI4+RUhL5s9n5PgLtNxjHTy2
kqSEBOWRStTQ8ofearx7zRXnTXuj4uThnDT5r69Qusx+ovnE3Bw120qwshCcg90L
Hw0uTHT+y9tC03ssQjlwEMwrRVCL1Ll8vnksrFebIwYh2ua/zDjTZAJ1tHBdeyOA
S9nQe3IlQWCM6URjRnUfGoWin7HP3xDyWbS+76+HXRojQR4GNsDWoBjJpcf2UvBq
+DWNdTZZ8YW6C5LfPQBPqNDOW1Cv/oPDyFcPaqGlnfFYMK6tnd55+fnsOqDZ9sKo
l/SvFPw9L6j8tJIRHF3be3m0IegHvMD02DWYQxwjcso824eWAf+QoPaL7GmsVlnE
FvSTaP7JegGLVZ2/4tvQZuAd3THaUIJThLumKJpoji/h/SejXmhN6HoLebpgHFOa
YXpQF9xM+KDGBQdv32QtmvdsXIzG4J997TzzaA47pO3Biwmh5XQsvKzze2Abs1sE
S47+7MOQRow+v7hXakWUs6+3EqiCjX8S1EOuUbCLh/7t31mfus0qjoPX5Dhd2UTe
riFd1swsYD24xWF8/AzncIJ8uSqEgesUEmbQSE8wDCGtOugD9DCs1pbrPXnCCq1R
6qdz+Ql/DZdcvEWK2O6i9Cq0pyYLA7SzCb8ihSEm6NJ8fGfkTq+uq5sFMqCIER8R
42q2vSMGtHcJyG933sw83WOWZMYNVAu3AArKVmv1D+2XJvHytEr2xS3abhNO+NRZ
YbN2IkopYHLPY6KgpYh/4DKXfKWM6rdoM0WddBKRoGKrtWKnxRy6bVOCZOoyfsQY
gmZFUmeLcZzqKJ9dGTZMhktohSzv1RoYbu1VBKUSjKTXheeWYEgncDyC9XrXlHBK
cb5xecoxdANeZsPBknMQJxR8PFSis5fa/nclhxvXnhtEQG6Y9hVSuYMej+X/s+/T
tKMWpdskUfkhaImj8n+I2YEenGkLhlAryVOg9D1BcCDAhD+hjIkNFmgOzBt5EoBD
LiY3WLYOEVP7s9BwO9xLI7uJw//g9DhHd9x9KqD3aaVfx/h2qkVk9HCbDsZSDXuO
HEkMkL3cHbog6UR0X3g2b3ow5NpRQgPveZdBvH9VwvVHnPfoxd6AdfOIlhxR3P/C
3JnutFEUjr4Acbv8YxHciRT+tV4O7Vi4RSN6BFfwPR7j6ul2z1wM+gjNFTuXeLIr
OSqpLVNDxKjOwuv4ImOwYoQX8CCrkVCM+ThiGMi9VD8m0fwN0PmpCGeSxGw58q3K
kbTkaRn890UWELaIpf2q3QASJ7yj5DY8G1GIOIpjIE2YBUIBAht6pxD13RhHHZSb
u/ic01JYz0RH/F/LVYxDnEa4OGk2cZy/JSPk6taYXTF0vZK5wSIEqcW/FF2kKD1l
aaqE8NgHW7rBrVkAHFCJaKBewtG64/jvR/NKmgCO4hyXWRc/bCUjHnthv3bpf/aF
ipYAdYyBxAtXMCsN2jpIHZ7oSdxrOhoQ4Eyh4btmhljUV8Zt7fXtw4xDKsk3KO7S
nzCGSyMF+xwdZ0MehK7Z3kBgS37ICAbOZcoRxVpVyHS7hrw0hyHNtXK+Nra75Mw0
J3+T/DgZrqdZ0tGw8TuwQqa2Mreq8kj2FvloTTmDcjmM5M118QQyAB6MlIUo5Pfy
kj5isGDNOcGc/LiGUknv3YYri9tbHMHZ+ZsE8wTf6SNzkMc+1/1kkHDc+pfr/a9p
uCW+twaljbz5a9LVvejPq7OYgL3QGmpNLE1YdMxkmPiktSQvDY3cjpJZtntaybwV
zrD05X8a4VcHMH6MEawisz3DGo/xL91uf/5WT8rAgcyDaSE+vwkHvXmGi2XslxZv
2e+ZdsZDkmtW9xvr15ZF+Be23999Ga2YyUe5bF1gWp2VmkWOVnDdU3Ly/LchnvQc
mrWzWfc8WbdqsmmaF/0tR5SwXVh8/DRUkjRIGz04WVRieNMoMAhy5nV/yPLmraD+
bnQ62zzMwfdr9zEax9WNO/Evn7t2yQ7KhwdNRkiTrvyVJohw/jNVGk1ds9z6JRmq
CiBSugOrti0/H7ylUxdP+lUG28NYjbhley6A8m/zGmUfdRr+lCerQPHZFbFg/LcL
9j3iZ5JzGr9Ok85vdQ79q8cvoXLeaEsEV6wF6X16dzA4XuSKkywr5W65ELKiRsk4
onYTT8vwOCopxlOZUcAw5SxXo4pSjtofgOn3sB3DubB93InJ4A5D6VeXorENdh7c
hsilK2nbZbYg0ifGC3wPgXo+KXWJwab+t5n2EI1Tw4wKNGT9KyTpZKRh9p9esuij
C7/Ht2Mux7ZQBm7da4PUCfTGMpbfmSiB8e2kXyiLAO8u1ziwuvw4gA1E4CvBuEXu
faKet4DevF2hI7XO5pmhI6r2Z4SGVHJkq97KBOfH7Eae28DH5M8LxNxPhKlD8H15
F57KZUHsP1Fn/RMRu18FRVWiRD2hWfx83iPSgteE7gaFxTChqdA1nSQuAlmGRA3W
5tXia5mXTPr19c0GyExuDKGAmRylk9prBpyW9XYpSlCj5ALVAnLHV6EBK6St4QUy
uhdf8DHrQXU4UfymTr2zPN/MTCDfvlUBJ/HkQzQFgC0Ts3H+7dREB0ycGCBBzkBv
J/LhkagM6kPqC0q8VXsxXd71/hB8bP8azIFic6YM395uo+dTROTnKnkm8PDqmgqw
gJhXFQzLsLetS0fwBk1/xnqQUL8Of/Bv/zBsnlO4YsHrPgQUBgD4FRZRieOKyEWd
L4u7+uuf/aReQrIUpGLyJRjCYbnBDbW5jaB8SekvjP+IpvJ0ut3zZrX4E6zx1EyZ
T6weAOiwlu+iysuR6+28mDQmOdvJXX6FOv/SkMMuu8pcMP6RYsbd05SNMPunS6Pq
ZmdjOPC2u8X0JXx7UndIi27wigFq624TT3hL1+4x+g4syAvs9JW3zUrXXYrS+ej8
rL63Zp77zEFO1qQLZgNAIZpQSz/fJ/3gD9wxeACLdBXjFthvIrzW+LAqNXa3C432
BiSoO8ZDC1RQcQJg5ay5N77rv1k4S64sZlhVRrC6NbFki5pTsdAkqqMz5tRiycJf
U/tfmyoCiqCYnNKhGAfmOd0i8pJwWrd46NAZ+9lV8lRo2L/QnmuBQfyxINyJMIgq
red6Q5XeC+0a/TFXDubprOUNl9bjcVjgXQQ6DnoIZYDaHeNg6cnVt7lesBJCV/M3
KEAH+clUls2uzkCTCT5VgdjAO6EbFolV9LfRT5u5JMY4PbOgP6TI2JDm3pyhodQw
DhwP64AZmqqakcT50N20CfaUWi27ttvc1ca2MWCsUoQeD97S7KkKkXSCPMphFg0q
Gh+CppUDwwf7I/rVBUBwG8eOjwNyjOCA7hjRRY8pe9dx+wNxibVyNwYXcOFX/xjK
pkpBXdAcR+64yT+lkTtfhmHSgHAMJEehQqTK89yP4m91OFM1ZgdsKmvDorqa3ozJ
Ub3mqiuKxHNnY508n3mZ/fsTMHSA1SgqqvMkP/u2XDvrT2Ztc8X18snwV4LzCQQs
ELcdVJUqGno/IQulvXlhSN+wOWWaOYzDGw/KvLPTZQAoOMlbTGgH5rqoLGu2w+Ux
8VnTkKaC6lNVibyUMYUwvp3V6a83eTK386yXb71ZkwP+vZMj76VPK+QXgXQFregK
4kqtcsPBSxiiHumsaW0zw/GL/pK12hbwwZdurAzF0lMen2oWGlW1aaW59t/rGPnO
USvEkQAP+RcDwtBn5d3zqTZRt/9aCtxfrdU4yM0G8I3LlIL9hs/YH58GzUbdRjg3
3HJZqRv2qXir6je04itYTPqFV0E7JdtBpfwjkCuuWzLCWu1+WcoNbpwPZGfouzqy
8jUswKQXKig5Jc/dPmqtVNwLhMGHYQPSzXUL82OjjClEYGKidw44MHy14t/kyKZI
SMxFnGMd0dc6oEe6NQcIwXpXhDww6kdIQgCYGLCRZ4vCGLTimRcdTPztU6cSY1MV
jxwRYe4eioVsEZatw3ohHN1zw+G3dgaY3tFFo2boEE56JerleIr2ppYCzgCNPg5z
Ab9iHRsn3yJYsUd23DPt7WWBds5KxMKr18gR30xARGLlbzleMjf8TObQteywFstq
+uDbCN8UGNr2lXKXV/pqXp1RrWeudpVZNIk0s3hP9AvEDLNXzS5FwE7lQ+cPOkQY
PXmZFnC7t/HAIncKBxjHQ+OLS1ZqiOjOvMcMFQ7ORQ3eKHXYADZfZGmn6Os1u80o
HoMG2E3cuGwpj9CNB6LF3lznhh82h+2m3nUHzGf7Dj5q9mrLzuBPd0CE01GFoWck
+htI38BzKjw07uW0YWgoNPEly+bg/Tg7OtG/w0brEfJzT0QcCq/SyLDjvlGif4d5
arsjkiqU+FzbOuJsKPWqw3jTyQ2aZC0+4+lB0QsPvY246Jl7GPjKNAk4Uscr20Et
mAXd5bjNQtFqwHnAvdBjf0fGHbmKYebbj4yV9iK7olvrhID2sSjw14wa0bXdgiCs
zS8MkuxN+Ydi6O9Pnpwgn+6EyLK1FKtHbvSaq1Qwe25W9yOqBxmOGKASVcNfZcHd
aADMIaPNfZN+cwCMlOG1FxkbVZBvl1Hg9x2zwYIYu2p3InAK9pHbQtVXnWz7SBwS
s5PZKfmFpKUhM6WvmIlf8RwMDRkxTx3iO7e2H+rw2W4jSuJ+jYfszc4C/mNR6YHr
LYSyhZ63mbYG4BkFh4f+OUNjF3gQAyBRRo6sAoNv8L9GTb9OsqNdebx1qzMCAT6e
HqxRYeVIveNkF53e32RIoQDkID2DCb29Z4e5igtx2EHOVCsRR0IlTWPf+lKvYZRr
/ZIxyrbXCZcFXTywvOGPB081W2f8nU4nX06D9LbkBmEX8rUv89a6foDhfWQNmyr5
EEAl8YjMdemrrvD4RNniH2FGrRqJPI1PakrDGImiLKYgJcK9ucShC8JeDIcoD4hL
GBsOhah433QciU0zcL+/ZNsFkCKv0gl+L5IiDJxlo7wRUKDwcR1GWIKHm4s3RVKG
euzt8qOlBBBwuLK5bpiIvnur+O0Tsn/87DxJewY7vNTrQO7PJDCxDwq4KAncNXKf
E66hBvuXJfP7WLfsk45qYRm52DqUhbK87/thqTLW4KKwM/F5Zoyt8u5p2u9tIVDJ
ra+5f6TAfCkp2gmwD6Hy2oCAG2wardZnG8FK+sA8ShqyjW7TcHGr/+VswN2aSvPA
VZc+FEhdaHA1PHrObANeSM8sdsL0UExyCaE/ORJeTZmLvkoXh/nr6K6adQHu9/uD
AzPCbSsb7H7bDICwUKbltLleQHdGXLCTZcgNka/livNcIzX2n9h/dw4qIUpLX4Jf
CQMA+da9QpyDB0G+uzkRXi4IUAxPdYoEdZ8H6CxBXGYePU4K7L4C136wNCzFcwaH
HirV4ugHe5n3DD7qw7NFBB4COFyDRbRmAgsak3n5PgcUTr1bcodWsm0RoscJ967z
jMGhrCeQ5bgqhHii1GtkBjHGwX7Z1uRp5sZ0QSm53JA9R4vjopFQFc+9Wm23HsDO
kX1/1XQKFFQpQLCiC39+GpvI5cnrhYi6ITkmeOn59ghnyR1ghyPwVimDu4yKO9/e
vKlp0YphyNnlJjGefllpIjBEQ893s+zu9/q6R86Qwr/MVS4FY1ibSOk5ctL1zVdB
ZOTEeufYsIZ4mhnxLh985il8x1xzq1qEjDVVV2vl58DKAmbTWOx7rccCN6WeBRcl
Dc/BlZfkH7HxmIyGNzlSZZb6YWLEtWDVpEWnFnhK6YvhcIAxU1bz1/+zYnIu2QzD
78zw8IeWH4UYEc4B4OACTbU91hbdw2+C2SluCp1sZhu7dcA9QYjacn6daZlnfpFX
K/pZXYnyxxKH3VC5rTrRCuUUBReXRg4D8awcHoT1fV1/tgUwuphpB3QhUwvrMlmp
xH+pse988xUWwqcXKFcfEcJu7d2GudzC8bTlr/KGWVs+G/VO61vZVktGuNxLDIkt
cguoao9SZfKxe/EKLxyfemRPeopen3cyyVciHEtdpT4dTsCERZTT/8RKIim9h5UP
OmFdhNgSmd8d5JT7BXC1SBZIuaPu/cm7mNFrhWk72OhXfyL2SagIUayCCOHRSIw5
Ftk8dEFLZLdqJxvpdJOZ8s7vC5Sq34x4FqWRHdhV0CMck75PfkynuD5y3cncQGu3
IKoVFLeSWO+Y4nRYEko/UVHVlKgmAjVBVqzSq4Ze71Y0SjDS8yCtMOq//mrJoB4P
MZWnnXexfS166oVH7CT+qB5jeWtAyPfPDt8PObdztu887qIoya5YreHJ23M5QrWV
UcgWZJRHmIL8dg3xdhUpuAAjxvDukzMQVymUu4W4Hsdgu1w8Qc7G24DTIdBToUp2
BUrKnvsIu398o46DLb/J+OFUmHiWAKf6uVf+nvTesGTqxkwHShysn5mR9Tf1oPEd
EHS5vYJdJgK523wTk+U06QmV0EI0tuNmXMDUa6MI2iEuFA85JOT52zBHFrPQ/4IZ
9YcxLHbZESUKksH7EVqZYbaH1YM3crv2VjoRUxlwOwjJwqUr7EapPb74evQ8IgPE
DrQHGflbMxwEvlEDDbL/sAzDnTohW7RPpnCRQ2UUka+fzE3c8ukB5QwV8wrRaLOp
d6X1UI4Zw0nq1D9Pp4V0ZPTHS7WpBijL3nqHVELs76MG2QJVRzHzMRFasXd3HrWh
zHdn5w6bjo9DlqEtXwAU1KJ9sfyWXNGO/6AN4yfsEjuraMs8yPn6DahjBaJIZ4C5
0yprs/iCa5LISh6xrFzQFpjO6a2Vk4ZVwIYyJY41trlFi6FSJJV4QQ0Ty5pedclL
2Dx2VTdYxQaI/2//rRX9tC+Afejc6PEQOA27ZOW4zJubwwOGgCEmtGMd9F64kIpV
z2u5imjXstTgrAi3gtFkqAtCeQhMNX7ufROM+MOP/oj7ih+y5Z1eO5tgwUxYrP8U
CdTOIk1UNQTQW4cs9qhhEi1pfXoZ4Dy8Sq/zozP8MHrhHVlQxrHds7x3Eo6yffWW
SnvdpCWCl8q3VyDsxP5sOGat61k467AmRMj1hL3BGsFTHjwWODXTGJQ+tpW0Tl4e
qrUPbZmeE1QdpG+EAvgxqrSL13dgBIqZBzQqlXjTVKAo7qZKpu9li7/GMM8LSrpu
f+A1jdzS2O+D06Jn7xJDrbBjwOWiqUBInXvUVf1R8K3Qbxmt2zsj/jG9h0nS6afL
8Ci7m9jQ92rkiZqhJOU6BhkIrYwaumO1wAiDNe2ESDy6YvOPhfVMkxT1AzaOVrSI
TYc/NzALKA+LLnyLAz16tXERqDajI/tzVd9+6SkQPREOhyuyf/YX+yxP938mP81E
Pvd9wEbbee8aDRHx+U4jVR/qA03KFWnvtspfX3N+0X67sHhYpozdbtKvrLGEMlEp
HwUDNnFws5B642hmW+fkNfdk3YSNBTF2u1Q75CYGu4acCPLDLwUbSB12IO5Qc4Ue
rS0Kyix52qt26eegQBe8Tp1rRVnF0ZradqkbZ+IivUdUjIYeO1UKZq2m7fCvsG8t
soGWn5IyGu64KsJK7LQDqO7bkMItVsuhS04wrDgosfxOGIUB5IWIjqNPJJ77RQSl
zfnmdjCcxd50tH4n82c9N9rSSFs98UTR0PLHHEnemEa2vK8Ob4VR9XWYG3P6zmr7
zu156vxMI299tkdM5OomHYPPtCAsjSpIhO7pItQ0KumtAs4wsvXV0VLv2+1I4UGw
1PKcHF7t9HQFT5cAjtNhJf8FplZ7jJoux/7QOKayu6e92WnPVdKp21lscQwFG2T7
t0G5aM7pXmGJWjDpHxERQFeQj2BRhc6pp6sAkdtSei237ScnWy52kuk+qES4my+D
+arqqxUKF9tBsm9u2MHdAYNMgWDeKXMgNyH03KPKpoBoFAK4vjiHjn47klECQgV5
LS3kbNwot/YwCKxFOZzV27M4hbwSdvnWjt77UXTJS8GyDCn9gphcwvjYXXiJadTB
eRdTMHm+6BXgqVb4W1+DdH5EZWRQK9OKcSQpopFWmwadzK8jutVQ3ynfWha8Ozm2
8vvL9Tmuv6QUg5dgnx0k1DeiT1cyf6EYaLI+UuQjQqVk8VWfNU+xxiAnNJJA8DUP
sceU3n6EuQWIfYgT7TxSHo7Es86F4ESQ2iyj8AySrtbiBc4GZNEFiXE604LgwQVP
60rFjURYC7MydXFgg+vsDmQkHBwZaveDFyAh6guALlrCYa7Lh8DCpoQMbKWPWWuz
f93Bk8QBxFfNwTPVn9cdzbUwYcLQRk+1wv04HL9FkEHRDUg6tDZ+5kFsguX5lAUp
w0TrXGzJhswTlKBS0caP4FvE0Jn3soYfT6mXHAfxAv1fdq7r6RyJs8JirbLf7L06
pyOcVsZEuiv3p96Eu97WzxUPWVw2uaOPoETuXPVIjhC4PGRZTfyOV1clEXPUysIH
M0cKv1ZfcYyjktJjK73sLQGeQESdXFokPuiAe1xMGddX0CKH5IIF9IDXN0K5ww8a
utXm/0I7EorWxNgaohuphGsbykFG2HIS6O4sxl3XBDCnTYrC6zL2f2H2HzqZ+uiV
jq4dQTWbyb4zjOdopTlA6sE04WYL+Jkruq7abBj3WaYvCmNGf/GLw5DzYa3nZp3i
r94udxYoLadFHqDaLmxqL9MOsLKxUFoxdj/A8BX5F7T/4XsmrwQngDyGl50P5hbH
wjJkt/hWnHxWfkMMojpmdgc9SPLUUZ+HDb26NH5jDieb/D4nt9c0pFMJm9GPKpNy
h+p8rkzlMpfPj7dUXGjheRbwBCLu2bzwjzkr9XI2YZNrIB8x5wL7HKlIoynXbzUn
yx8mY+R5C0hca8Izw4HzDsqCNc6ObGlU0yQk+AfGMldKSu7ktGwTe2wqSNwLFleA
PxVSo6tRiY14liBc7vzDmgtHeWnZsJDGkUmGxTYQbk2K3kQShMt9jGb1um2SHIpY
jalJAoapxWYbCa/qpfDj5URTukxooJSh77XsnbHf2YyNXKVRfsnMkSaKp4i3tLvl
P2Id38SWJCxenUQH1k2AeVA96F5M6r0ic6IC9TXPJ0EAN3FUArKIMpFNCSatGqQQ
BipCF/7qARnu7UpDZKGVD/Ehw647UTPnLN4ngn05fFdNeJvbzOowoeetp1F4Un70
OI4CtjYdoo5p4b8imLV7vZ8mj6YEFZ75KU+2xKxbWXAlBjwhoJ73Zm9Fxde1yI05
y8+5jWMdIjRkrevwCuNduobQhcc7MdElH9h44el07LXnhl9FcwbpFLOP0MrFwrca
bT+Mlf7ts5hs4TytmkOky2Dfyspr3+UUqLP3ypCf5R1M/4Uhv1V/XNno4CP0ZzmI
IUHrZUTEjEjw0syL41F8rsZgczGpfUsSmjlh2JJcAdH6J9FcqfQccOIbQrT5r1/0
cLHClU6RB+wGgjuzZ7WIgvG+Vm38Nekny0jy46hLtyRY69ir2EXxffcYf8JnWsZt
f6nKKYZOQJtsG0okHGJKYWsRcJl7v+eNVCmRBOsPp+inAMDjKQ1pH4ux0W3lbb3d
2GcMBtrbHqx1CqGoTfywTYhIFsEUdfexwTG9KWY5BUu11fbFIgfyAi0Z+WdQ8Sbz
cXywP1QPya8HFvHyTtjCNL8JaW83GaTWOy0+A43pjoHcLmFs7mSTZ8LIB17n+vtx
FOHMRNwpu4doRbJY3Xla76HF8PSkWbwk4W95QS9bEg9/P44w0fjnvXbOnQ/lU8ga
pBsHWBAQglsVMKglhhE6ciSOjzvFGv4fmyRt/uSmMzccqFIkFgIVNFb2vvDa/YQl
M+8dEwVdGykNJcgJ4CA+LbQavH6oXPGfWZyRiTfKcwISF08d8ZK/4jthtTl//i3k
FeMrIAy+Duk1wBEp+qU950VlURCJ5Uzob3Lb1m/AlWO17Xf6s06AkCID6xavrjV1
/bbt4oJPi1lt00326qCGz/xOBMU6/S8O8/1kjHDpBcV8GZfjuNvpSc052Zo71+5G
Xdg4j1PZ1L3a5hwYdhTQ6cJqB48jD3etkuAWIJRuy/44glx4YfzJgWCFf2csNPAe
jF5n8byA5nNbCjAwO6GtggLkFNua10UzUaQZFPWzlATJPXnzrRm82Gkb+hlIaYxM
pucpKdkM5NIqGZR56t2pvrZROTuT6hxHAyv6u+diR7+9ZAYDdWlWuW0vn71xRzf6
8/c6rb2yuQ0sFzpk6VlW0RT+3wXdkzT4OIbx66HVK+GAdVZxljEmb9RV2eBB69Jj
+Qgkrrs0pExtqCxNXnw7zhWKO69r6EA/f5AcywRBTKmfdEGjxoJXn7roek/HRP8E
PHQbvCc+IsDJbyBrhXZsyu2HKW1fX7BfIyq8k0diaU1jPgFJbyJ2477wYd3FHFQ0
0BFBrTw+6Mund4siEjQVdT+XEfWBVcXGKmXhhv7MXEsiIfW8rUC/lc0363rdLovx
v/4hFF3LzkjJ6TCMsVbnU1yXfp+DdTtZyMZ0MSsiqxRVhbtijhmyJ4OI6Wr9EuJU
flxR+3tfPieyZHtEiKr8L35Q+V1gkQ/TJXXvmIVaYpS6Zc4xBQx7AEqbomd+DVvG
Prt8upUI4xyJow+f4voWSDaBda6RZOUZW4z9TJFT1+bP9lSf1BHpqywjiETSaYyQ
kddQ7y4FhjaG6i4F5XhefG0m+YRIBXoJpdIfyXMPO3J5rg+sr5W8Vv6dHo27aPwL
vyVvtifd1kfLS+yxFhde1uC4SlKC3ZW1nsFMJBqwNVIzHD8HmbYHUHuupbgHrRZh
mbpcAobbE/71PuRC/JCJaxRM+jr6eecEbcY6dW7Au/kL8k7b7szoO2oijICItVTl
o/VSjlKRfgYz6974mxelfL9Ci6pDpY4VWtv/+zoZPt8oz7zcOc5gypq/s5c6FiHh
6/6u75xC0Bc6+LsMgSJwAbuzni5qxdJ0oUReeiFpvMSkxk/hHZfs6k80sgvw/gFy
GQ/VQ5m/xet1HKw4pNPSA44BM01uX997SljHUvdTJ7tskUNokl24fKU/X3ARVQJz
fss/lFHvsz70qAD6EEvlQaM5Ifrd0r4i62ZxxOLsgjRrq6az3DJ727gA/t3FX9Ao
O0HHV+vi1lHTFw2zgooBtKlHW4HgOVdaOpETS9xZBw+cPNWtWSLFmkr5N7USHkV5
P7OsotW89kHY/VB195KDm/38YY+bCOBGyJbGxs3hnZQ67RKPLkdSK07UT/06jzn2
4jFO6sj6hNIUIuPLOwzuPg9FWP1BUCZjx3L3OTO0RKjBkAiasMCa8ge4CScWxEzo
EqDGIKE6x1v2MZrlXrRKpFxvbzDRizwVp/u9+fceLoOma5YAfPIpYbqsETC1b0s/
sxe101H3+V8JRbDsGoy96uyD1rKe1xxrLaOZTmSanKUc8JUFzxIOk2MigXA2tr6s
hsqfxPg3hY4LUXdKnrPf0nNdgy106bBo+0JTzAes9O2ruTsp75T1Yh4on86H/U/c
uIxEBAD5kapAaNnZGQmuTGa6KozuEZ105trZl5oiuDE5T1La7bUwaq0y+4C9CrSv
c+qDfbUbflNJy2uUUp9kZO/CuidkWTXsESWPfKmL/V/oI7ZqRJqMrV6LuprRxQit
O7aG4IxGjmXMh3027YeUVgBLXLg4hjdcniHb0ZYqT9U3KfpjuS+ElcSXBy/tkvZ/
5fsZUNUr5vlBsln/imzbEPlHhb3hh5qof8A+KlMUrlXb5E9/FXbcOpkHxoyjiUpH
wTuDhZQY9zjcdIQL39t1IoJuJ2mrwQ2yb2WqfXHjsBWOphF8f5pNf6vhdo0fAYsU
CpJ8Jd3eGck8qwyVsbwz3VSdva4WpJVnDSUK9DN+mDAuL9DaeA34sOOzt43FuzSc
f5eqV4/vS6/dCv2lV41Bauqn2hsYgdoURXCuAfjcJZ3DMaS5gtSpwsj/NnNfXhuX
1DYVxv1zL4uxuJTUK7C8y++GdXPUWrFFs8Mde4PnRnKGkTSYLxwwkaJaD43zu2P5
MZ82+UwnGw4bajuD8OljXnXGF5I451T63hsNUI0y++OXhBfxkWd83fQYxwxpqFbe
rHJuD2q7lr1tcnAZuNBaEnBcS5zt5SCvtHJihvkNMxWWzllXxo+Lbz9iA89JN/UN
lae3/xWmceIk+2iZK/RC8wlwd2SKCdsl6kYKzZs80wEwknnrIGCVuW4+hUaoaSL2
+4PvMmIFMPLj2kof774cpM9b1h/a/lEuuoQ7+EmdxyIHggRG0Nd+FqPVxvLkkOoG
gwnuqqRx7BO659KCULUffaXY7Yf/M3nctAzzvthtseOZFitNs8o6/K/umxAVs182
sKRw9ZEwCrliRIV7WLtY4uSNEutRJkTY7jBW0JJUt3/bss2WF8zPmq7McgPXQ85m
rHiM5LDJxCkOhpHj/zNs4GTZdLQtUqchqnvgcqLrO/j7ep/5zxl4GNuq9VXcXQv/
deUw8wWAYl9PfaK/jro1a0RK7CYapbkBf1QvSXrI3OoH5auiGDroqZcTETStyhD5
++8dFNvpv24OlnG11rics5O+74EzC9xyA4TE3udWWmqrVb15lTUgJu3RKCQfXYvm
s/Lq5dCNSv27rIYNW0WW5VlD6VOnsdgUpwmKRqQk5VERSMmSHlHJmsdCB3FLh2Dg
/wPpyoFaiuVGxezNuczdjxuAo9UpbXB4xvjzKyfRFlv8ZBDzwqFxoJW04y3+aJj3
sTlEJmDWs6CffhJxnQSgug+ftrHmsi6iwVr1PT+viyaBP0htVnk+Q6LuLi/L/lT9
XsDKXPvrJhGjBQfWTDpqb3ybLHtnl8/hp33GmJCPkwwhrQX5LC7xBcnUnquTz7xr
wsrYc3r+AzdUC9ramXs7rEHhL+AD+ZEgR4nr5u4wEg7ytqLxA/KYgpcPFgpOkZl1
pVNIzV+CE15yP/S/wyhw0dW9Nw5SzBtw6u7KQ48PrXqNCOR/BmGx/07cBo8PPvlp
9QGN33jRh9LnDmZkrZhQsntnSRUCe2Z49UjnIu37gJ6tQOILEN+Ql1X1xlZXeeVS
vcV63KE1fHLtiLIkm2u6gYEc50pyvHr78Dd1hVLlFAVOKzlcW+6wfJZgQVDt6L5v
U/86Vi1buNAdenxUq4fL69lq8/9PeRrsXG74bkdYRlAGHT3TF9Bvas56hJ5mgWXn
vJHkpA9ES8PGsFiGmyAad9mWpjD6KnPzGXyV0TesyWXerkRZXpJZmXLewGLSQMOB
nTj/7nD70ONBzxtCRFdZfwMU+dJUlHe8PmFGjKg4+QHHR8dnlnYhGyvuHXQ+9cHX
j/UN9nfa2lUQdLrGQlHNeVjdxsFnTguY7Q4Dp7fymHYhyOY4ch68OcAoHqHeZdmS
le6RVwdMe84Gj2dcBm1y+tEqzN19qEJsHq/ooDrcLlN+ufDe4vQwTgDPo4xGDdBi
e/x78G+FWZvsaEYJyhV5Nrn5YOp3gqelTl8zNv0anZjlCfY6uyD18fGHQn4m5Vvy
MbOIdXuOifkEymTSafqJeO2B4Bq6zuhlNQwd9pXvISB5qAXOgGWmJEFDL8NpXMYh
5Lfjgz3EXwz6qlJ+syVusgmaEcG/vqC5S4L1g42OLJvNRsirm2IBmm3JXraWVcsG
6/xP3JJeG1zOVxCZElbGk7fRQmBNc7TsbKeq4dJHrMwlOmOXU1PUjTlxEhW1FjG8
jJKqhj87maboV6cnNuoZLSC0w2qFeA2ylEWLj4GnpxPbQCS0Xk//fjSAZiXar+8O
zWiisULE9ofoDU+BIZKk85C6no0XK5trmj8ObaudSHxQt47t9sBEfkricvkuuQMZ
0u0gFCDL/sw0Yg3/evz9UYMgxWypRXN/weA8MsTaNXsURBNi6ctJdVGqkSxhRi/K
T7qp2MUthPFrBW4Q5kt7moKh9yiiLNwOo6xMQR3vQDjEgGnpO4cf76Aj6ipGADfc
SN9dxICOUDpykoXRQpIb6Bl8XBvvb/fn9BJXExb4w1iCKi2lh99wJaYYq23TLq45
ZNRewoKCUzSClXu0DO3hHck+uZIi83laxyUJ5F2B3e3aAIHdiOTGSsOo97OioQMq
zpXu1awbEFvMFcpWJn8yPPt7XrEjy4jPJv6igMukFDyu49663xiw8LfC0YFcKxP8
doGyqeqjrkRmZ9n6qrrcGN4d8HtJ14E5Xe01z2SXHCgpW+6nIC5bDS5cRtPJdUBg
CFsX4gYSdin30fm/k6QeeSQtxxsOBCwHwxZUOQFIMZx6sE79smKzgsJvXyQSRBnK
pbdU9vMZ5FG1cjzNzkIGKuFUMMYvyXt0gsj38GMSHlTXyrj3Kx8V5ga94Lc1Gcr2
8SwCDlMYzNBlyChMJf/E6ZX+INAJraiwsmCBGpjBtdZtKLEoQZYZfyvKupdiKYSa
DayYiKnXj4WvvJxCcp6VJ+2u/kjA59ngKC8DSB2wOhsFJWrd1FLj+7CN9IOON5D4
MgZtm51tVYRCdhcgjkhgYH4UXir/ntIf76UhTDrn/j5/9ZTTGD89QhwPL2+7Ar5z
3Jognhcccc5rGaU1/V7t9QWpS57c9TRRBBJcePvzJeQ2og//gSZxnCpYYXeshLYb
bdFETOUcjalAIFU72MYak3aa3Xa8vY6YJEO2fyOUwWcj0XjwwE6LaE0N4Ws7I+G4
fLoAhja4dGu4p+cNaC5czY6l9c2INslqokEbPaWkDHkNohHjHC6Cfnm33+zr1uFM
Lx1cDbHptq6Ut6RV2+lJe5cKlkSylRueDYN+EX0E/bT/ImhXZE2VSOTbCsGXasci
0t493926G2dth8NSNXyO0Q8tfldB1rABuXoenIhB9q3FPozJDPVn5a1yIOP1TR1S
lx/xuwnWJhm5Hy7fNYGOzuMFaH3FXIIJ6VLD9yv6EcskmsxQSs8al6tZFG3Bmrzq
n8l44qqAImCnY7aCndasgdrWB8NrlFEF2G8Hq/dmLPOAZkLUcZo9XYbAutMne8BC
0kNqQ9BUxtiN5daCn87rEX/uc6qpGTYM865sVpcmjyy/oEhlLred2WK8xRUE4S0n
PGFgPDw58Z2DUs2BjAab+z2uZ55YDGPGZNCD6As9Y31N8v0SZbfQo+7j6OjU786U
TWwZThyWf8LCPzuQbO5sQ1N7KQzJGxRn8melDuJJP7DP3VC7OxtV2nrE+XmjGeod
k1VmQBXfZbB0J57/iTAmve/CpbbGPH/nmYJM/YfLY/YYKJPSxFXOn7pGwQBjJ6FE
sWB/2kBIouNOQH7wWGxlzBU5LOLLt+x2YXD2rdqqQXVg4KZSMiG3uomWPEsqlc+R
AyI81cLcLvaP4QdrmhrC+lQgXI0xuLPpCAbzDZzboRvgBnpTzdLRdyScDbHZhKPC
ZtSkYsu0T31vpXxk7LOBt/tL3FcQaLFg8ypsJsaOSAcsJVpfJkoCz8bbKo0b1f7w
ObVBL/LN6YsMxEhVWNSSIT5IUIcKlhxLLCeJVyfC0alv8yj979l9sIGpDEWbR5fi
hrIMNUbvLGMqZkpPKvwWEzH63P2YWSezjMJCISyXS2Lr8aZ6f0xRg63ntv0lvmoe
oCx26Nt6phtqZE67rKYAZPhh1zlghZm2isa9EJbL/bSoMXp9RG0vfVjo+nnEV5w5
lihSu419SFZOoiRgw8/0IDqmQIeA6AIA69dHnusAFKHUJ8HwtftVNqdNfhwriRjo
HuKHLC0UE09djPxt9XIxL0yax2FTGomHMgQx9qUnEppQTCmOfdtZpYwpq1kWomjv
WlYJeQhooMWMvy4b7Zq73Aegj/Yp9eOzYyojRzyFKrce4ksBdAwEuGtfCTSbe9zK
CCQ5TLhx9eoQBST1cSZNxbsRFc3HMHlW1dM7bzqlr7rYmcMbTAZDJkVW3WvbZNny
re0FYyY2MPlUjFtiJ2ho7P6tpf1iM2qBlng56NNndOoBV7Ck+dxyVIxITTLcUSw8
+9NnF9NrLmtia2Wdtxt41Ant6UnyYf4FPt+iO3PLQL3/nr1mXBn/QqahwwBTUAIg
Q9XSjSicjU+x1sEJzG7jqiCdA2wNR8CEW1S/fwEZUy4vq5V4Coeq1PttOPYNEAVb
/hJZrV8M/IYcp1o5JAGB68gLK1a8wUGelQ1Wkb3uUDxc6lcYb3oEXTmOub6i9l40
wiDARbl/ScacM5g40KusGulKjpt/9FIsggUhl0g/t5Z393soPMvac+6FSFCGRyO/
7bRne0z59RDXnH3i/JaJup2A+gKXQAnhofPpJOXPeIpo9rHWfpJZQGXVpn9A+ZO4
EAd1DPgAG3aUZL4ZB0jWkZiIlPvJGCSm8HvSRyaKFyCmprcr0iDjk47RJqKlrVme
NaaI7cQX3kP8v+2RAA1weucfgEXsbJ/zgNJuY/bR3O9Pdu3dbpP5hkC4udEaCXzZ
2P1dI/fLiADPnG7V0AjGcv5U3pdbgpOVto+KigOlf3jKUqPSmfW9W9aTG4xp3Czu
slN/qLGg/3lrGSn4XosxtBTFkP2DknRAyZqhEsf7ANExhEOHpv6UgUOaZApdbEAA
XFFKKqLkxxp3ym/oCZYMf75lKQG2SRTKZq3JD3ZfncnQb5ggGiuvZv6ihsD73vNg
EEW9PUdBUXxDTNG/0GUOjL7tnRQL0oA2U4DzCgqawV3bzmznmDGXjEXNo5tCLe31
1Yynjy/Wo+6sdaeQF6liJQUKRA2124dlYxlpmHudfkXk3ahNHxhNVUp8BTAs74hW
sqySeSzh85voG6DgSV6Mw4wdLJOl+7hLYq7abLpDh7Z/RGRRv8SclRVCCIpSBr7n
UHNUL+8+4aWl2EYtH2s9udy3sY/N8fIsi7F8yc6lmqhO9Xfd4iK6q0TJxoyluntS
18KCYeV4t3on7AcAVJf1uH6tZS0gJ2kd6V4XhjMMaZCAZw+ZzGvTJ6HMqYBrIxqI
CChKCrDTxdGXOIahSJNEUaRj90B39ihxgpcRLihRkjYbtwEHaNtEORajU2v5hpkN
97ZTGyuXT0ClKSQtxSRnInGot9iYuj7jTvKMJwFE4jUBRo4O+ZzlpgZH7T/Jqdkq
p2reOVHbOTumEKh4RHeeGKSg7X873KNwq1A0ktKYrl4dbHTzP+p+mDIa57uaCXRc
iFqlFFfs8DBSJTIarIKWyH9wJfud7PnsJ4UCY2yxbMOcLvQAjkUW0L26PHZKIZb4
P+Y2kCtQwRbCU5ySbz2jZEN5TwWTgKCg92m1plxaE89KYQM/U51C++hPwNSrIAin
wRX4Z3W4RAd23r13P33cbdAWwalh/dWSPV/JHm+Il5opJGW/+O1ZZGMWxZAt7cfW
NkUAE7jaYzpTGKZA/dNhWBMM2smEWDJoHSOYp3UmtKCrLVrPYrXrrzIc6ip5naje
1jBxup04sjrA77pLTR6gOzoANURBeydpVSvVIwM8yg8a8QAUb4eF+LdDA6BhB4uJ
Kqpwnc6DF4xYiMj76Kbt/gChv9tlXYtSTfOcBo6cKJsPSQg0G2oTKNmopvnMUcir
ttoc9SeQo1hRB/apHikw2DavDuTfYa/FRqki3VPjmEiGIGwbaF4mWdfRuX3OQ8Wf
ykK5lfnnE+sXBfUNuFRikuGPqXnUKDZOxC4uxEpOw4TcC0uEARI80AiaTbcVUlkT
AhJQ49YsG6YVL+EDqiacmQZZASNRYlh9w1DOFuaiUpZgjojKvSZsoDmkzPBxR/hN
4jDBrb1huUJina2hpCZVVHFZZW4HRmbxEeHQx7T0/L0yripiEqpmNAJ/zva2XKkK
8MRytTOMzImE+BN55g1kGb77Iz7fcgXBZ/4PEX2vxtxkqOQk/SE9ehYqEq7fARLN
GRbWBlyFIvAmqmJVSvUcFBXzD5EZ8FMQneg4iHq+Hkr+euT27z8US9KyFtPYvQdw
HfLZISNJUTZsHUhfM3ff3M7KvHDsu2lCw69iULd50NadtvCMfc2SEUE/2tUCvQWt
ztAQCzVpq27sHKM4qnBpc+06AO2VSE8C5jrH7QAVZBfvoLEYIkcILVvsVS5uemMe
/wcMuFL6DG8GOvG5zDETuDZdAztYbgqLiiSrC1wa2fryJQx4r7DwFOBUR6I5zs+o
e4Ibhd7W4tZG/clMdwaWnCEI+W1Imoh+bKrlb5mR5FPOm0rqlSHZIaNb+6PcFEkQ
FexKb91qe2DhBjeslPFnnyzVmT5NPUO/jO0eALc+gt1rUVPr/8/qSc1p4p9j6+ib
CXNZfK5UOv9aPmJPYljLSIKz4TWmY4Xx9Nl4hboHB4h97V934ChoEmDBg661VQGm
MpbImXrO4vIHGYCBssWqniS+w8+yFEXnzWR0pd7WPk2MIwHd5sDCB/BrL8B7jEsp
bDeDLB5JTbr91innp+g/VbTRiT10ku/l44RIbnDwYV/Mtrm7Fzzfkp4aQzv+oFKw
cJGUtY8CJRiDr6IykDWKRK8x2IfV/Ymj0/pkqbyFeszJ4iUTR7Zs3Dk10KhwnX15
m8QFOu9hiGLkDem0yMWoj0auChfV2gzR64dk+sVB6dgVXzFXEtV/BpLiD4SREnZP
AQoFURwFH1QECSHS8BufFksDaba/1c223/Gc+0YMJd+2zkxFE1A0dvWQrp4Bc+ot
wU4Puu3d5ws5eOnLO48++RvsbCHTa3LZ2Q0w5Y12kyuqUdWRvNCurvot30wkndQd
2FJjI7ZnA4ZdVrDBxFvmRFqrL0s/KVscFvVzleeUW6QdQUMmsjywzNdnh13Xcl/P
D2cYk5Z+dDeogMY2VqucGDCA0o/kA44BY44vmRVBSnbyRBk08cLGpFtjb4o0DWuz
26s74ylgA7j0BJbrGHM2PezTo8f8LosdddnKtqvsUyr3eYZ+5A+/xbT4i5+GH8DG
lybVs+IDJqE0aTg+gELMsUDmUabkt1QawBvojLwfCGum/9+q6zo04g4KBzokVm/L
yhNXh4N8OyzpE+LVkI2lceGQpWp+rQ8czA/lDgU1ZMdXI2nW0OIS+aHe3uAsCod4
6yDn1xOvrQtbAT6VrP5nNVLkMaAXQBpF3zLni7WTUO+P4/PgOK3O13878gZKalkr
Px2BIv2eeEiRAQdwvug8jynRuTV+H3uj5OhvLdOnLi77cWaP0koL41epsk964Jez
R4x7eJHXDDEvyEOfKpvheS3NFJPKVoLEN4p6Gk/CtiTgjsNe4bWnerKtGHzahOKj
EHDdm2xY+YJv7e8K6e8GleWxbOoARrqSHfX+3ovGs1sDaxEi3WswZg8Hr5sBhs2C
yt4yS6fqKuh+xKp1fceF762bgwJ7q8H8oIx+ULDSch6rQWvuqBte+jNnYXLspE2v
X2roF1/ryHCtxQAJO4zaRhmwgnI7AbmCx03Wr+p7X7dtc10NWL+1dsAvR6nddU9V
1DrODf2V7ROoFmhHWzUe3nm13jHbbdnTsqv5PxxPWtg+8fHz51zRI9cIlYdXYX/3
XLQn5yf6hxpPAQNcpQEO8gTHhylHKF4NlbgLe+gLsVNf7c2/nGTt377b/QOjARyt
FaPlnCATQ6mwVwclLYtV5iWL/gbvmJHFuAa76WMpFvybFRnqmtJ3xfhwXLZ6ug4Y
LhyUQDs7HfVk1EDNl4Ij0Hz/KnJWfqTjEBznMAmEetYVia4ZkRybX/xUy7rgyEpP
rT9WyVt0lDJudvTRRRqrQjV6tObjHEamZ6jA23yb7ZxWB9mhfdD9lXCnWExjGWf+
H5Ow/7n3NMJ/FRXLHHoTShkMY+9XetosBz2jdEY6u1o+Ik+ARmf3kUvXVQxbBBJ5
ydOEmt864FHcHCBlObDxmpR0JNIZdiEEYkCR1/C2OHWTl04h10EM602bd+UfbXW8
7Fi5thXdmHziA2AmUaEv7GT3ugybXC+Kj3IrW8VUQ+g6WW+E01Vrh4Fz0Pvxd/ck
TU0ls9ezT8GIGtBE+DXyXoVuZ9V5geEqu9NfYRtyifyxHrXNJkubz/2wn+Ehvtyx
Gv5/NrPpALNr9W/RdgidXNJW7/GfKgg1pcEQA7/CRVCrW1LXAtZHPeKm9ZR84Yw+
A1Vvdg+ZT58F96UajH6ueVb2Yv8c1KbGw/5K+QuJLqnvSL4k8Rt/xRu4NMwU3Xlw
stQD8E1ukDN95DHOs8kW/GaSIXxAcKoWLOBIF2TAG6hft+/3pzYzvQWEU/l/vtwC
Na9HjK28p7OcDYLq6d/JQomHFIosZOBNpwKRxSJuHm2aWqyWj6l6/WpmQryDt1N5
XfIK1ZcvLvp1BIEfRsiyAgFolfboVzWnP8l21SrT/cEJJIfb6Gi7htSHreZ2jvR1
S8tpGZjnhkXlq6DP+P4O89j+VB/qtOsWWU3IrlI/bnKlsdfR4O4k6qnh/B/zfjaV
MAdVirmTFi/T0TQ3+zBnUxczNjXaDkucmDZKACkL+ud0xyCVN9HFAfbLwB8wWABk
rtLjlXhWS+GnRgPY6kqTulJmi3WoWZhPOaJmL6TN6dJT0qNGlPboZyikGyXrDaCe
afmQD0MSuV4KgAXt0nV2aiFODG1dI3JmFm0k7xbwbsqIWCq+ltNMLS2PqQtZE5h9
xUUSLomKNR6hs9fBam1CHQJQaPmFUDPGhXotF9naYHMhXt/EjWja+yBeOBt2gXR+
0hQnfAyyTcKnXOYPjMu6ZdwXtSRq50wT4pAhiPsH+VuAaDibXieBnO4a8qs/VcGJ
prTh8lBr2LQC2bi73myhBsjEhb/VtULbjSm5goi16O6Eg5fbEHgjtfblmaTuz5c+
O8WztdUpyaILoqKOBVvki+rKPJwGE608VDRMvqOAxwQ/2XRIIPvV2nKFp9Te51eX
3kLNVVS94K5wJiwGwpsD1J9JmKelLtyK9MQeQnbLo0vloS/pupzYC4LObxR0CCOv
iSquuVEj+n6XHjMARPVdFE44OW7SLVid541VdlIRL7zB2RyY1PEJKo9qruxY033s
DoJsun1Apd/1A3yL4KA+o2uTY24CJnEKNwCXJFqVGPr2YycwHCkswQjZfQ3pFWsZ
Ivusns7KP7Sv1e0v/hG8RGRLP3fUrDOi04KWb/ajA4zuNoKiSfgX8+UVJIVABQ4x
em3KON7lYudqC9CE6NpeN937lgSLWPclY2/lfiU1QnovyOR+/wEYS5nQLlWx9A3I
2Vlh//NIlh/4S+P/jT5+ZnUyfDgC0Z3lXzyJPF5dWZil1BP8OHtU/v/kw2fPvasC
vudRgdMG7f+XxZIQ5HDHtFv3hKzLNI6k4I3wwGNDT77g13gnIKzkNMkBsHzRwfE5
PV+bNdzK1oj20VsBOwGy57e0vUpfyIFcaXET8uE2sNBMUYZEBU4lkN1uKa+zb92H
eIS8nKrBIp5NVo+QqCrdVfO3BnVBFSRCVkU+ZMAFjwed85si9y5pnrbXJcBHNhFQ
Nrq678ihM/6akczF60RGwXxaLTBd3n5CHg8lkG7I541LZkrfUBq2Q1Kq8Et53c+t
CLg9jfEGGMxD0I3MYJTJjZod9xQoVxHdJVlrgJQT0J3h47iXyGzPFXFUmpCtBwA8
S4P9Zff2vkudoXf1OWYOBCARio5RWwQed7yIHWEU53CnlpAdXiTdwaOV1SD1eBtY
DcvRRJp/ov57tlZ4oooG6PqSX/345IXKZkOmNpUsf/sQFa01AJ4eppVyY5M4Ebc0
EJUhkOzdQH2Sfy/pFgBqB6E5z/4Z93KXZ9U/CnGB9gh0JZiDKgmcNNU+gd58LxOy
YUA1MlwYB9bH4WBz9s7Nu2jfQfJJw8udEuQ6zTKicm9wsdlKT/N4J1YBG/gih3eD
5Pqmd9H586xiLAss+3T7KjUcIsK92MJqYQ9IAYsDm1E9NyHdF2TIez+AcoGig3IT
3ZwXA563ptQiPBPpPrKrRGDxyhGlk+3zJR81BLsgX4PTdYJ0kDMvZwJD2w8DvJ81
3rOo72Em8DJ9h7VCkiHQvUijh0a+IeXlH5z36jHCybxkbGE/9l2d+o7cUlFQfkdd
MVmxr+T8lkPRGIabecV8kwAWvRAF1p3wNYQ2maggH5jhlvVhAU3uL7Sz0am+c7Id
5wh8O8vLQdFzyxmNKPPXcoyaOhdm5wJ1GTTxHTgjzj5HIgyUcCvdHlMSeEpRbXLV
6lzJcHrFHL+hPg2qSpYcM1/czcNsUoqvV3D9YgLH8Sbdwn7xtIUvTAphiKDNm0Qm
iL26fYV1PIDrPZ5UgkaWlxIXJqSzW8AKOrNPxRCa9XhfjAxKTHoGlhMgnTG7M/Tm
8NB4ZNh/VqpDYOSwWHn1iwccoVZ9kpAQysaa+h9Vxn7RGbIlb1HrJLIFlJz8so6X
5CPTsbOYffSdQKZn+d9SWZqpZzDGC4D/BDGyBnumxasymzrxkjICb2AHhiw1OlaU
Voni0QwV3Top+82PDKIIHI/I1YM2cCjiEgCpC5XqeAcmeBPDrNv/Esuc//ceVjNS
d99LuE1UDoejI8DIP1+ie/GGsdAPc3M+Kdd02EJjUObBUzmSlTH6LDp0kFYgncLT
1O5Jv5EHkFZI63uMsrCoJ9En9vujRmbD3O+UqMrprXdQH3DGVCezNX6hmE3A7kaH
oONPB6/RbnDZ+ddweI4kjFH1LWCK1Rn6z32YNXEdarBLTnLAjAV/eTpLBOnD0APM
z/t18jaovdJNB6NPzmmYDj5AN5a7/8j5ANuLN3Mn9fMvu2zmLcFxpZtKjlxvkrSz
XcuJf3hFswkgxqrhsaftQzHLpOwkfJPBZNDkXqOR1nzgw0f68Xkw377eVaBKf4/R
bCJt9TnmM46u5xcEE4RZ23SyP8aW1H5CaB87AXrJz7UEazVJENUDrye5TnVfkmcL
mx5iSXuAOfAwN/YT1Y9hZTSp8i/rOgIb6hX/D4e6fadtzKoIMsyx5j8144CIVnv0
Fk9jjcEeJBdykS3o2AFlmSLMXLjln9QJaenq5+G/czj8umM/JK69AHJddyYbpW1D
G3nlW9l4ayI5B+idG7x1ycoU/c3VOa2smicbnPvL7qhOXU2zgEjxqwCkzmbyFCkG
Ceu2PHlWJsgwA6ZFR36iPwbFUXrvlLBTCNt3RHJHIT/DTcE81bW948ilSFMYzhNN
Y47FcIRpsS+BD7lscui+edFIZrFARdtk15Mg7d8Ek2AtRE+mSezbHaZkK1pSAtm6
6fZeZgsHiwGEtB6s7uB5RZtEL0XzGnq3gE5pOaLuWXtSWSJ4HAKm8iGLeOEFniV5
SdO5bSjau+dLu5tMhxAV9nWhIG4vcRj26hgfW13im+ejZRdn8/WI8XfmMTqOsdC6
aVQseH6DtJOgJTHJPP/Q/98hVN9nviVPTDPFrAsjhVfwrYnrblqvx+yV4lSBMSsf
OiXND25bvWM3mcJnSZE9D8a7FVyv7Vvbf2E2QSoXdlvjsSEeAhstzOLPH8XnPMYC
MxJd8oJJGar5xIqAj9yu4JA/0duTr9wWLhdviuocBCAskQgtWgQqGLvJNZJ6V9vx
3BUjSsBM5umGzsbK0mnYBmaMitrUvJluGt/PIQmdY+HOETkK0jgn+Xm1JSCJB/Wj
EixHyW09f8rStO+yGImkvH25Cyvuwapc9k0tfMwQJFG6P/FkaZdS2KRo9XpI3LkR
MCyXE/0pXjvGKL6jqWfkTNpRLSKTTEbdhkTgxKO/KZksCM8df72kFlQIxqr4+1l2
32Eze+n+f/w3/JraPL73MU6HBjpj/r7p4ghIo2aPqy4uxd7/yVq2VJNOQf3b14Cl
6bzIbuZWz+6XN00sTPb/HVJTxUJVr4PfkEKJEY64+6vXboE8eq7hyG6h1SBSqv0B
WRfqd0mJzhtay3beLxi02Vrbq9Y4B8YFd8pEyA3XCWVuroeg9DohJorOOwSX43OW
UacG0YrfDgCud8ypR4pTQQ0LjHl2ltSmNVTmck6Ut1HG8BnHKLtKnfjOgi+Iv1Ls
TVKaK2w7YNttJZ14xck4vyAKVvmk5QRQJMWCDDsbeSS2Q1/GCXzuAotSgxXt3JAE
RFih0F4QAE7YK0axbHwJFg+y1MmkhUi3haYSjvIY8xusKl5/10DzVsXDMi1CuKWL
pYhueZ1z6k4sGE7KnzAfA6xD9cEOYBCSk82TYI2ALXIxCJ2S1POXuDF+0b0x1BnA
JzIZxwjE7HSKzaBSvZBPoPTMr+rLu3Z2WlRmbNi28GVGoZUbzKJJyGVExNO+AN6+
2DDtPPX3xdiipT6Lnx1/+hdhB8r+w2yqy3ZpByNOlwPaqIZlZwPQYxB1aznurHe7
2VdvCYjbm/mFu4nQUSVb9S/mG69vQQSNyp1uEYfYk+KDOHI+nyEErLYxP3pdmKum
0b6cueiIthlsJ4NKrb0mhdcbAC4b/64QWUbg3nBFxuwmUSjsBKnmmHAH9B5FFFdJ
DHGZP1Wo+mUhMUrc+GiSDW+KiJhVDwA671EwuVhm68Ho74gTw3G8QVVcHrPRkAWG
e4LSs1McyIuD7hSE4ADeEONtHb/FSZ5UeH2ZEXHTBfBm1l6N0PYoHrdlLqM5Xzy4
9900cy8ctYYeJsWF1JRIxLchVkdDv523DiFuiu4Dd4qr3jhDnyaIkF3mEa8kDfal
R+jEMD5HoOxm7ATLzUF5iMejiLO7Eu3SlEI/XMFa/oRouD4WZVjiwF1X8UjQ4+mM
Wnsj8sEael6hj1I5p1f7IAgqgJdKaB63/v31zluQh5vM/x7IPOkKklI9DnbdLAl7
NklSERjP3n6GWzf6Pa2R2nG3eBGuOK/ydxjKtTQbx1qj4Xk6AMXVleFExoGAZibO
2w0E6sYSlrp+tkrxw8pv5gD+0CM2bGmdAmGXJosV1yFTlaQA1pienFH4I9yKZx51
fDd249+Rw4Y7g/sCMJfeVWY3cxBCeaLEoN8lhLzkkIEnsptQz6abWnau9y7hzrM8
8dT0PgP4Q9dSLbbNk0DIL4PeG+uqEnIH6sNJoycDpsiizA9tFAbaCozsZ3D9U1TU
ECcSUnees4HijwGAABztgP2zQlp+B/Efzyb/K1gwZYLljD6vp1ArrP+03A7EJFED
xQTTo/+Hf/ANd4nl3qBhglSJBDgXdU5yRQfnkjHDmnEphEtjE9dowRGs4r4JI0OU
7QIBhWAw1q1DlbYK1WBGYNZQvQbzFCf43rRSN07COkxA5IQ6MhjrsRWqHwLbHf20
/uUsPVP03iyyZJlLg9Gs0G3zz3nPHX1e+OkHruvbZTG+BRVBzqyRCV5AIvrdHU67
ltKh5NDSQFfaEsTkLaewd2whbsHc/mst7Bj03vcIZI7GsV3nvnntFsAFzuzdfKe1
vlYbbF1j93i8go9QxuhJErza7WW3W+C6kN9wZUdyuOzmi2Y0oEiup+7Ed1EUwW2x
Z+XWtARQOh2HQDhzVQjB2y6pVeQ+DtLOIMcSOoHG37J3McTfgeaFIO5HnzkyLDZl
dDmv4azcotmnjdbdJ/LVZD3B9a8hFteQzNXSIQWQz//A+YTOEfV6vGtCYCK3hHZ4
DyRtCU9d40uebLS3gSiejpWDsPKBlGDtmrNwTKVICSDjV5YioqGddHWKx/jfZIXL
axAJaQxriXFhA2eHN3juSSs4h5sf+izc6hcujhwQhE3AYj14N9HVdx48sbJmeQb9
drSNqxIajyZkunXbN8rMnRoiOlK+fH9N+h4AMUJboAcjn+/ioUSe2EY5g6woxCRb
UE7zx+pqWWcXHnNk1s3vp25G8wYCBXdwx//3vN/3KSYVaZJviplqianzUZS967et
ZUOyZlnwIKUfTyOw7awq8GanvI5XRbeM7Z13jIFHSDhzIzxE7+20i8o9g06fFN2L
Ge+mkJQhq1ova8VPXvT4r00WlkOWQpd1bZgNUzxG+96FUBbN57/HRJRgTnVlIJAx
q8Cxf8K9GM+KG0GbtlWAThoKobn+Z6BZG62BPXsKjvkT8A2GXwK2e1tZbNGc+lnq
Smqozbx9Amlbo21kHlqsmWMZ3uliU8e+/fOgNzCGwdlvPSTqQtXyA3JaN+RaVjuF
StXSNpSDr1n0IVmLQ8wGrhLTbdrNwlSzUodqX8w+CDvGHlG8n+fq1bnpb7CFZEU3
+5qHAgI6UVIavM+FF9g5swEtnzhLS+r1gUVo+pwbSKbEdhJ9zWzxFB0Ro1kzZfar
e2xvDhXnS0S1SungJPWUqsTsrDhM5FqQHn4Nx7wbBdChm6wD/q4CRiMadBisikaa
PnjNJkk3brJoSq5OeXWC5tCBZqm//hCzpjd2QBP6042Zllj/ODwCCLlpSBVlC4O0
Uqh3S5SeacwIy2Atzjny99VK9KqNFuD93/2/urdKn2G+wiklKQgCkRTBuvbq4BTA
f8CuiVVCmXnitS/MV313Of+Xs9ebYAyYALvmt0hIrSETNqVY+umZmO9F+Ev2/BjT
1bHLRAo2VNAz2TLW5jho1ZsjUOqoWlzZFkCcfjJiLA+C601EddnbQ7QC516Ibqjt
bH2xOBeh0raFhUCEend1/zgcFHzzocs9Q1X8Uzqs6LYjQeKnXN1y0eM0BG0ltB9x
zyutFy4O3aO0oP1a8qTIITjH2V4BFf4RwI7L7cXqOHeTdZyNWQmWboVUUB/TiogS
r4V523x4eRYWEDxQ4v0NckEuULEDaMtcoZp8E9k3aaJw9stlSSTPSXKc49Q29NgN
Ofqz9S7lbQWejYZI42i0GZEXNd6t3x9ERm+7bJ08mUwCx6FwQtYyznLiG89pegY3
55O7wBxKgCYa1dGEL4uggMJbElpJDIEKr1GCpuZaAZcsIX8cmxFx4xDRSJ3XSX9w
bknU9RP5gKD2981GARw0+Q8J9nuobzxt5eS3Jvwr0MDpvmRvJRa/0FgctH8/9SRl
GDi9D/ol28/oxy4M2a2mESv/jhbWynDSbN8RWpMuNgRWBj86kdPkpzPBrzCfi6uX
TaAsig07t0UHVzGTaUieD9VBED8HHfl1we7Yb3GNxLC0DgFSb7XbT8dr7kHCaNbT
0qzP9GK2oXj2LyhaaYF9EClCf/POcSO3Yjt/l1TbkNPXa4f5A4H6k7EMG3j3+SJY
UMU6S1tvDBdJ3qVAcuz0iRsYXZIhgLJB1eG9l+mY3QpIyj1SDmvGKRIGy0ZH1P5e
6XpSkgWmVngQpkZQFpLrwM3zrR2VAcm2dVd132f281mSswYDH4B2rPvdriGhkCNb
2c18vtnlvWJU8w9Op03iQIYwON1feszoi6gbzDlSscCOA7BxzH5Tuh7nANRTbrXK
vzaimL25pGIWWhq5SDSmdMFb2HV0+s2wyaxewNzX93WDiBwNY03IMdkdirjPj2s0
HB1TRZR6Qq7Pt1AAmsRRZcyikmOSZfZuZlr23cGJI8HbOR+ZVEMDmSFpvFTvcDjI
c3mmJZrTYmkbLNe8tOjRTD3xXsq+NgOU1RVyxosuUgXzptudPXCzR9/2pw3BJfOY
Daq1wKSeVWJ3VrkAZ9YdqXGQrrOFq3SXaass8WEqXmpvLzhGT1GiGIjZ1J/n4ufa
0Kc0E/o/4gz162s5sTCtyFjPWMxDrXq8fmEo8flNZc211DVtTc9xC4G6unPGNvCA
FpZbkPyOxBfuWB9+9KGKAuFM/K3WE9uJ6dNL0gMrdIrq45ITPBxgvmfT33U/Xw9R
i7tkFHnPAwnYSvNL1DOdLg9fW5Hh3/91mTOdftG4Gt7Vau0jY1r/SN2gwVc97EO6
IVfmlF25u7B8N5xJ/MTHF28eOGlCujQwXvoGmi3pkbTcZvhVvZA1BlGnZyc7jglt
oHB3kdBAlKhSGwMRkkV8hIk3zNE5BBpHHi99jMuWIYl10K4FZOl/z5wLqu8MRJGL
xPQfDUydeUdwGNuPAui/s+0D74rMBtApqaSrnxlRQawP8lmUZnz5jA7tgsjPCX/X
OGPYVqYcR9Pd2eH7O5uUtDp2y3OryikeewA0Sy/7vPwnWp5srVaOOzET42w4GCOl
1kqhsmKtp9jJFfuunagBs7Z21qTGJwUOHceuE6JEJAY8TjAzvu8LpSD/pv4gv4rL
jB57XkF6KFxIZVKFEwiA6k4GQSNoRKDTruQWGntpEzRl3c2SuVaZKUQUHDc64sVo
FNUTE4RCY53LikGUrljriwRerhECqBZOOgpqqVhNmu7jhN1h/WbWLqSpGBeH+LCo
SzWCP1sc2Db9C20/Pr8MrvUWP5K0Qnub1P9clARN/bn5gEcl6XOxG7X0X1PzcBkv
qlsjLzOfayvvbaJDxFBoVK5uHjtOG5A7tklmCvA0/ANjmeBOoerCZpgpYxr5QQM+
V2hLismA/PQrC/m1UkYANOMdL4I81IgxuwxPyVl6Yw3wjCjhcizRa1TClLids9CV
ACR/BXPcBjm7sUN0Mek8+jne6VkstNdzflcOh3KciJJdlXr4C7ehSqFJHO8fOyL0
mJr4V1yAixLhWGt2iLpSkcj8YTMXNXkk3W0tSMLW41YlCj/+LD2MYF7gqoih7sfU
IcsJpEcUuwWPWeDeT52Hn+lejilTUgaiBcyBShwXBDUIkuBiikgTe3e761tMgAZN
GM9MzTXimbfAlA02+dZbgO+RmRW/ZJ4kjt3FJ8NjeH87Tk/F8zox9vMRsBByxHs2
53/jCHhc+jx2qRhqA8Zcoa5nk4xj3mZSeuomFfXQSebP6oCzT+opnK9WjUsmDwu5
gzlunevjkT5osduvIUNkRiK1BVaaa21Gz0ybeREPSMVgoIQZMlFY/Nj7my4Jv7oQ
8NMtB28JeAgXMWHlj8DlBroVpzSaEkljUrHsrofxVTFUGntaBWF3h6zjVsENgN9i
v5l/+h4z8c44JKFlWD4P1rxqeZZ6FJi2ZWUm8KgWRzd7Z1aus1MmXfZoWCbl/7Mw
ETuJ70ngc5qlxI+HsSM85fb0N/U5v63i/xMRR7KuOLDlvb78+vJEeVrLuewWWGu4
uYxP8GrzWUmKA3W93sQ4T+atsS2Gb98MjgDorm7RxnJh3A8ieDGBQi22/sRaBpih
Dqxw4m2vTYImbc/21pTtK0jW3dQQgazqSCvkAFl2amKvUFGP72rwSGynXnif3gcM
RKlh4NXjDHPa0OOvYgUm0RA5vc86W/CbSJUv/AywdDTa39r/9eu/jKMpGEuYjx6Y
lZfMLdWuGUNm/9xzolbbp6Q3kQVLwj/Bk12nSybkB2TOp7MbZcwDjeMBqFP/kCeU
NH4RKR/YJqIMTIFzriC+i9KSp5gaXP+eIK8bR/83rQoRjyKEIJKUe6PNOa6CNR3C
MVeB7vqnSO26eAWmVJs6zP0f11PHJyFJXxluEHepPQCQs2qol6+y95JXcg0lSg14
PjVHk93PlqF4/ahLpQclTI44S6AZpgNXJb1FIcPiS3QI7yWT8XorJNbY8nbG2u7i
C7zXauVmokeTw7AAkZK0LwrqeevVjHOq1HNc+ONhA+D5XPClnpUVKYROIyr5CoWb
hdBD5SfEeVLnr9j4Ix/xxy+cIKR0z9oSQFUKu2+qFzvOSzN2BWkjLYGvJh3/OxIj
0GJy0aXM2v1k+xQ7/S6Uu2xtWtGE/QWlr27F3yY9FJ69D/HbEJsws4yJiCwnf+B1
CkrIEfqJDrraoNCC75vkVlJ5lsd787uBYXM7vmvd6p8kr6l2SdQ9LYSb1Kq08PdP
1kf4riwuF+naT5Yk2McZSiibskx/3PeWRYf47MOxZpDGh43SC9lpJ8rJG+o5/9LI
A+eyI3I6SkITLRLvJUO+5P4bpTzKyNN1/1lx2MfCFeJgQKjWYnoHi/+gU42e3CCv
2PUdaZi5Yl3eHGA6my8rrcM3gJamvbZ6zeg6Kxpz4RBo80TeqnvIwGNhx9cFoxpD
IZLkImbNBC8rtDinz2s4BB3NwDlUu4I99CeE1Qxuf2lET/sQWZ2ZjJIBmI4hLIpg
pFnIovWszX3a7pAgKdYYLd6bRW3Tre/f6VdmT5gmKZ6RzF0LvvMTG8F8NcBJTu8P
mwEk14+7QzniH3k2AuencHqAwS4gtweqi1rXVjQ6pyMKFk7Qy+zL/bmgFNK3Lkm6
K9YHP0v0jLapbFYlZNvHvrRUglNFkBgR0YfIRRhY0H1penh3YqyzFm0nWfRLSzLW
484NtPeuQe/JDXG60WISn6iEjnTVlBvddC1x4TZ1CroXZt4pdbLNQVSnqLlUsRe6
2k3PT9zsIW41rIsJkpmlZV64BwYptreTeMlaQng5Wpj9KW340uh0Iej+0g36/neo
sdRPe9T8pH4cWn0QpISlr5CsT74UVKDxcA0wxhs15B/yV+zlUej+eD1J2QYhC82C
dJwQlSqJVod0lxR79+5kc+XdNWZ1v8PYWVwu+yV0D/KasFKxixNn8zjIblGWWzA9
gDMX5fqNZG6Avy2zWNdPkGEgVj5SV+alI3pFNZTg2U/pIPDmGFGap06osEE+OC08
iXSIm3590+2GlXIGL62jqKLAQ0XsmKBK/8zIFcJO6f0NocKzEH7m3fgQG32QlGfS
sl9zkN8EpsHhvOZvR/XaSazCKbe2DX9wyQXciO52zrAFDuCca/YAeR2lw04TLYm+
FyIt7zvPc1ngjbgsKdivjP3i/Aqf7mu2kozW0q3yjHQ3/1JZu7JY3hKR2Cgnkrmf
a2aDGYl8NOsWaHscdUwRZA90NSn3xp73GAIo4ONrcbkHiylIYdwNnapc8zIWkAUa
HSzsnXSkGpWjwRQf6ta2jVchK6llnOZoPcgY4f2LFvudGon7qlzzUy/gJEIwXUtD
04qBbASu9lJMko+jHbTmP/HooHVCh1nVl1yGLh/ORFLm7yrym/7/pfvXiub4hRTp
WcfDrdjIJHJ+HIu7fHw+gK/YOLc/25eYqQOtPGWbEAqRMxhUOMxi/6GRLX85e133
S1HRet75HZGpESti229uzuWuZNt6ytYMpg575K35YtDZxwpo8beYvvWNCAdzVjZj
AW5wEtULBpw4IT+/m1Q3frOYqXd/yJ2SyxFDOpSZxGOoSqMAAj4pgBJ1nRu2CcOY
sLipHT9jDvOAbk/70ScEICskJa+FXDfVSXPHtsMkjPVWRpn5eyVIEsmDqvGshU6l
ct/dABEuBF+LxlX/mH5UXFxg0iLUszuKVPQ3qCINfvDBKZPISZ2Ok+axohhaVp1Q
5S5ynarhri91CGMaMIt0RVRpEyBUsIjOpo2fx5s0gv3Y0Zqf3UZ1bwy4ux0pnZhd
5O4L1eng3iaKgpt/mLVYT6cy5K77X7kMFfSmXlA0cvLViWFhSQC9VgxMfkFrOlul
o/5g+RtLSdUpMuK9e0/3qW4/KJOdshd5eEtgGCBiJtWufli+j+W/PfRgTIafSg+a
3WkaTWWX/ThrbNr37BvKbPraWSNEH3xi8ZTwREPanmSLV3v96es1faeqGDOxQfpF
Q7AYN8TIEjFhIyOcodffk+xcMgvlDc63KCjjOqdATFQtbPfL1cwV7OdL0uzKmo89
pSjJvij1awUA1iSIzFcsWnxqHWiOdQmD1eXX+Ha6ms+imIV/0XZsYeohs9+OTHkb
Oz+iuf7TsJygdp+vRP/8ekbVsq7LKs6hd7mAXl0Ft+11Ht4Axd2N6GkUbl1ebc41
IM8mb42ew0aEgtCL1iqWOR6ju4XyXG/ibb5P4bvVVL0f2syQwjSLS/mAblErJhId
Mc/fvB0m9YgwIJL7oIh8aYaOcndPWwxZoXGPZAsXE4/sXQGOfENm00PRmgv64wk5
AlwUtbOvhiYhZ2NnWeYFb8T2Jsph1OwJcllJ0TEbrk23FZEpKrsoQaEUSRfbOSkQ
DUTcaZuimVr+oWxCOZnSTInRGyvxhenESlcL4hviwpIFRgHa4n6CEvFgXyPrp/kL
+Fh+FTvS31KN8k4e7xMKI61LNvQGVxgjPT9wrTVDVqiNBstinS8EeHqOuXt7lM0w
Zxy04Q4AmUEmraeuk6kSBj9YryJBnMkAa0SO6sJPVMBKuVZElFnu41CENSjMtlTV
+u0ZE+8yk5xAUXH8bQLsfWA81Nvs/oY2wL+zU2u+mRc7vGUnaTT2/Q9osx3EpwR+
Opm9YR8jGxrosO4+WWimKbAWhOGfB/iEcCaRxwJTYflno1W+Dgljk3fOOrggP4O6
+7iJNBk6Zn6qkuddMi8j/e5Du02kcfy06B2N/EZao43PIrzhoKHjFc39eHo7IHja
O9U9tArnizHvUvFlLLaA/DLXL+g22HDaKkc9JJnszXKOWd0721H9UziPeH2xvxvj
n/BTGxkVtJ1AJ4Y1gJLLLy888Rq1VeHgbycl/1bePODFR+tafyKYfAhFYFnbXys9
pBx3wHm09hW4ePoia9m0s+7n4GAwJYbtVBTgiWw/FA9BW4EVyILB7lVKF60CbjGt
r3I1Xc9XpUjsxb+mwMWM8v3n/sLpQPR90Nw0kZUUQa8g65ogSv1I76VGHQn8oqnV
1CO+OU4psS2F9T4imFuEJgJ7XPr4GG2xTtwBVzRRgEefrsibIq/DinJ6IARN1Nom
YJhR8IGRc8sUliCGq0VaxjN4MtBSBPNpnD++zhappgJSNKHvCnX7CbDoyNeY2/DJ
G6UO23rK+Vmkt+JMNCNUnwmBk7+2OLCsoK2YDq5zfSUaaXcZREiMT7vnM0bdirRz
aUps//naTbiDKVfALKDZx5i0Nn3CZihU3C1I9Z84f+6ri3Q/iPfFkKa5Farp4J+b
atuowrMkVgVeV16LksRaQbKtLRsZ1UEYWn5Sni6ejDFvqy8p+aHRvlU06IXKD9F9
/YIZ2qH6S4BJW+R2LeghAVozf1Y0cGUBkZSeQ1O0mQZpD37Lbf28p7Ved5TNNxMr
iuxBfJsCLPOY+q6+6X4ONusfxUfA69bFgdkjkbT2x7hCgnEvNyj0lGTbQpApteDn
wBxPossq0k2ywjU6BAA+3A0010opQ5MqkmssKhDObQ56lVzdcsCNcacwb92JX8k0
HtVOS2FxDmiIP0JuAS4P0SRuYqxzUNfbpC9DfFGmlqS1+hh9FKo2RZDjk22aRbSg
QZSma/OXy/Fx3td7aqLWLq3qvJDKWcgUQ11icb+X0Vm+XhK9d/+gVQC8xOFlr5sG
rm17KKaVM+oytd7iBlhI5F1bEmmoXv03zWDsrWPjXgitSob4XJCR9UGCWJ3/lJEe
ap2jKPkKY+Ad/d+luo+FD5O8NE8v+5iyOKnVGYGbK4dWglirMQ+vG3Lyr/uDcw6Q
OhJ/bWd5n48mApnJCpnDjNzFUxEBEPM9KA10VBU7QzDqeQnSOV2whLDD9aLNmHta
1zqmStwF0DSwTOfcwK81P5aAQfSv9SV3+hOuJ8zwCpYq3j8UBx6At9UtvsEnKWOT
K+xKD7YJnE5ww9W6ioX3Pc7F7eQMRTWLL/Y1ftdzdiAW4OUBTKvrEt9eimITO2we
l+1fqfQmiqiySF7+fNDGKOLBK7+eN8VVofcXBs11hInqWSyEn2Tan5SBcLsgRcEc
5IvIn2+D7Pjs3jb7Si9jkVz6Z6XJbX8ESa+c43mvTlE/D1jLZEQtmud2h8QwI919
++eJR6FT94uploEh4gNOejWbMNkzrRy3cow8E5oEXuVoViNnjCQ831tnV3lHSQwk
fPQKqn0PVcotAVw3uHrY6MzUTpBquNpdyYhVtj4m5W5KhUThbYshZ1xJ8vSQHwM7
6k6Vx2waR1Cg1A2/HGzeQLYyr7ytYSgFTFtxZfkZgtWwYinyQiS/7Pz/VKOhSzny
AHaHY/DIDnJixuxZDsF4vvAvT/RDJ2P5HUbedwgI5G6IsP2rkkNN/FT9u7YZH8u3
lIJOvYpjtrDpFIHU6ayEoO3hhvKClMYcdx35Q1FpRvOmjwg42QEfdUaLojOtC/5i
zGqkc2xGlfRcDmCjQsOSp+sYb6IzIZ4BRlPU0f2m8aJ4mSowUlWZXE59lF1xa+0T
d6oNtXY5SukjbXKSqiNtHcAxkOaQaK6UZA24RXKsR1a7WGxtK19/i1HwhOPh44cv
hhzHpKIxGWLGXJ29tffX719E1gL8Fy1Luz4DK/j/Zsb3+K1LP0ROTnvzJSrPGlto
i0wqKnGrdGpr6xGWc6GfZE5DarOFJBt9zOjvdAfFL7SQ2/AW8lDq9/7BbgBEgWuV
OLPIKEje6slWkUrCRhIT1c7IN09csuWAkCau0YjSUMsDT+zBYogP9oMSg0FNo4Ss
17E+Ct3GqUMFqz2I04G2nOz3bbH5awCuJct99QuZsLBId0MG1jvNFWVHUN4veGqc
wl4HuEidJLIADQFvh7ODOy061EOBSQmEKZWFbhLHThkkYQLHzX4b003UIki3K96J
2jG8iKzH2+N9KeoCNR8emTS4yQhAeZZ3U+YDTfSCvNL/qT8ZydLjAMDTgNp7iI3v
4fTMDiwzLgTzka7eugWHwnUsHAxtDjHc6g/iiLdYho879Hhysl/TMMJRwlVu0+IQ
mKNvDPTP2Nq4xWFY5yOd40pQsAMJW7kjwa7HuYjNs12RJLvBzmcshnVH0a1rHk6q
btiUEnIAbhskdwaXfsUR/pRj4Fpo0w/gzAEOIP8D6ejq/lsnCrvRuYWd73WaKhKk
o0soHcqOwFYO3IlD7gqi9hGulxjmwsgvzjjrcawx7vZXmGq6hYq223/EFmVrAhBe
jIlazdfPrVcj+BadtZXnHGpdm6c3EXRfqStthaxdUdKa5cvcW/RkAL45noF7vhZy
mVqsbVHOIXvDR9xdaBSofZFphkhcdZ9QsemdhxO5hvGv0vyqn/ZLE8nlSHN/Xn+T
VS4ZV3qrfJ6sv8kNkM6lHl6jzftrJ7MYhIKlN5xNk7Qkfn7BZOX5BewnYIWL3TYN
SWPK+uw2O1XOnyTLWvlBTdtXP5pfO3niSFHP07TlWl6EfMB+b48dS28rStfTN+C1
dK5yfvKUTo9LzVD9lIZTJg/PmfzgYTtGB8OQimboN5wn5QeruKf7nAw/h02/sLYV
fVP+9g1v1M/BITjPaDhJ1rJuY+Hr7JABiGEGwALX2qJfhbGPTPsIgZDXf3AnIn0L
NTpTK3HVdBDPgvum97zD65BOvFqZHC4NzySbjuwp9gv8MXcDux2PO6WzXtjP32Em
eserqMTChrEdNLL4XdtSAuXAKgt7kZQulHIdTesbwdlIcUJdPQ0wz5IgrEh+yOrM
zgp7y2O7i4bouj9ajMM7HIv7Uqqywm7iIb8nVS5jjjfB6yt/YpW4xcAhpjSr/Ff+
lQZt+XAGBir0ZPdKdDdlxDWyxeO6rQCJputG9oluNHJhsGS445xmeRUYuBra8KpY
jrI7daitcVUCOjsYkpemkd8p9KOu+/+2CZWWUPrJIxGWRsWlfWLQ7JgB+YBAaTQy
X851ld8zeOoRcfozpTB1QkTtiHRA7gfmc4VnD78P0F3hg8X0Y9MRRXLVN1NwzB/o
K8PzB6hZwZRk65fAdeST5pO545MbfOdDPXoutkLnfRh22vqCqiZkmGIrOpM1mC+8
ZpHlQhMjw5LdRJZ0BQtKBVbrNc7D8pjlYeZBgfztZd7sjbH0dh/uUKyqqJ2qspoR
HxIKhoR2pDWjYdp8Klbl6ulhp+nisD4KOAPM/h+TxaciJJVkpNWDgA+LzVrjKpr/
R97VvlUlhirktg5tbDg5dvmEzrp1mnG0bJ5damD3+oz/+FTfWNGgAny6KCaAom//
R8nhnvoZSdm78gCBKWkRPKk3jnnbjU1gmUlhP1a/WYeMbmVkAmyqkBR6WlKntve2
tpyL7nC5ocUoayJ07j7O2nZOhtIe6BPG1LSnpW5e3V2nM8DOr9wm5C5FcuNNryne
KOfjrimnyVv7EhZNzWTk+8/1kg9+4aLzp1wEhuWij4rA8ft16bC3YKz4E1DtCopR
TNgnoKYLWIFmlVvN4DTY3nJIYiDOy8FkrL+/49BLfQx5d5OyMWonTAmHlIvP3U7R
1LOheZZAVEkTGwAGL/wTYl7830ovG+bfzMD5g68voBdjJs5oUJgHr87K8y4ET79n
bTA/4PeLEe8BE0SDDJBLF12DelNM3lS28pkrlRQjibnQ+Fp5j8+yRTTjQM9wwrXS
x1PG3EcNgTaOX1OdIZZVdu/qAN7trkRfHdaQyxsOtZQGIf41KHws+wYcG9+h/3Vz
Nbr6mKBsf8ayQkI/0aUEiFG1BWb19EM+M6nsKeRkBsRw2zHSDk/+mHoAPehdEIyu
zajZUiDk3xlHTYwXOEDtSV/jXWiaqEMIO8xt2rxUgMW/7djpTB+SBnpc4T8rx1OM
D385vGOO8Brs+WKu0xYwJ9EzXQoPZyU8bGnIGKcc9KFPTGytCUHk/WmaNSvbnPRS
9TTmxOv1jHI9mHD5jvj4MyHRyMLcHPuR3MUZ9wyyTHwkR3DNnhiNfsH1mGmA7frn
QC32xNwzQ2yc236BoHnTiKWYGqBv9wI0n0KT37EtPs83GQoNQzQU7L089nCerscV
1Dn4vufnwn26SXuO8AOHbKrjMk42Lz/PPddOyaJLeYrea5ASE/igapqs2+EsBTT2
4NDVCJVtvwAHcWZ816ryWr47bxKvTauL5XrTlwDq4b9gtsDt6s8czR1OyP9JEuAM
yMeBWOl4fg8wN79+mTjmp6u6DZUSngqP9uTWY0MZ8KwIQwCFvhit9M1BNprUopG/
FRsX28kIGi+sm+LFSvaAwsarjNqVgiNQAV5oH1kaL2F6wnzV1hyYbYQhSTX4JpZv
JshmlplHLassiv1pPA3XmQTFKM5ZKHvZMEAzHUQYJ8h/6f/3DKsDyGbywDQLr9VG
PryjEBAgXMMOudhNkTGbiAmgJeaX4yTR6ZvZgI7fNTE2DHMMk0z2O5XusBcvuF/W
0aTo7iZ34dzFKDKygFfnPDMQNpqaiYmyKKf9lAbMIBrKGrTyXFyvEendtspFe5kh
mbS4ldpWpwj8S9Bt9izmhtEL31k6aQAQAS1DMCNJ+QlgUBJLkfpzcz5SqJYkrASQ
hKbzZDgxGhzE+OcGLeQlb5Pb4gUnFPXi+DV8+PqPQmZTzrsrNMZvE9QVkM7MNifb
/yIOsHI0qYCDu4yZVaQniY9d2jbTQYtewQkwHeDGikL6VBRPek/b94srDX30KahE
qRvLTYuBjlh90OLYFV0E/SMjTCqH8Tc3HanvcqyT7DOG4wAQr49kqt/MfimsLaIk
yTb67IsCdWCFdpGmqsSyPiDG9aRreCn/XbfcpBKCsGD2QQjd8jyKQ7W6zFDPr98F
pTYAfzvSwDINj6Nj3MskKAMgaCf+cwK++ZQIg+eWCk40NuQbbN+qucldZsbWBri5
r+nTkkQwk3WRhAFCAKmUYD8399/QqfElKF/JlEKzuRyb9soiHLvZGkS4r8RL9s90
+nFzWAZkSQMRvTNquVEreu15EfKiMZnYAY6aMSI75qh3l753qXElsY33u2w77v/c
6y2RMUrncDlEP1mLe/G6lE/NaQdxdnQF8P9KJ4ReCftFhWEBvZm1+7TrYme8HaW5
eOaCpFBaPDoKphLjpoz4Vs5lM4Ghl1dwMyYr86hKVd+vTr0QbIh7erHMWrQXE7qX
6zc9CZd7TX+HmoBkRVqIQRPYaglvWAzHwSym2yFCTiAvO14k3Bx/JGG5kUrlRQww
FBE2KAUwLa9NF4zYONuWA6mRSyRKH08E0y8DNksYKhJjolCoPGyTeO890OPUlVcc
XMHb6CZskQm061Bn8ETTv4ZweN46WQnH/OWpQ0bhCdcsQCQuYZJpte7tKTrSGdfH
2TXYuWS4PdhxrtL12kgr+q1TCJc5HaRVBsB2wqnMufMYZ/miVtDmi0/wnh7rrF8J
VoJf7XxEuMPYpfrVihpjDOvc+DXhDc4FFe2mAVZhFm/h3k5vRWsrhKDWcahm02mi
HjNp19yJZmsCDwiiBiLS/9NmPXb2NUK7ciRkWwYiToUL7iWZAttygK9XF2lUhRny
sGpgWf+rfk4tx7M//gD3b4m+aW0XtYwFg4pzbLyzTqhzNEzYx2sA4iPiF9WhiMrT
YzI4VrrIl5crdyGFArDTFn5Q1o1Tp1zK/MHGSoLNMD9d5hLZo8Po+A4bxi8bQj5D
hqmm3HajOlh8fbMOnKrZ5GKBroQ9XpcHbvP4TV+uryoWgO6eq73eV5ZS2WpP3x7F
x/7xZ7mBuLxdWOqvfpVOaU6BjAY5ehRg5A7DNLunWm2Wupx79eOUH16DmF5Ry+sd
WZWxsWRQMSigmIaSnuINITYpaw0llb4+v5uUpc0StPInjbx3bA9qN8vb164N/bhM
WVf7oZVsl9DNyJEOC/uIW10id+wIbgntG9625Ga8EkFvH+5IiC+AqDsehZsElGFX
rcnTyl0RmD1pF0cno/Y0d3u4YsAFgKTU+abg67WrwqvYW4KPcw4D1wXfl+dSLosq
02qF9GmBI/QbJByOgy0BYlZz9WOFVTdTlqLiQGfDL3F7IKLbfzG9yn91TOlYh0Ti
QvFiby76dTJUXG2no72UngRwG90o+aosUaB2+afg3YIr2NB7KiZCZRF/49ULz2o1
ZQVvEYGdSGMNDbTosP3plcvNZlX/MHefQdBvvuYmOCgWMSLA+Q8YmJGfvb3nCqJf
LCiGHB9UdY2BDzvb2EYyahwCHTjt/vm45mHCrxEWeBQuF4vWJRUzAWdW3w27MeW7
GW7vMVS6quQ90YzEJBJigwnQO9xEmZd4nY8ObFK1gQaRz833mDjQQJ3cMjxbG8o5
UPXkzBkxzt14FGNhrbatVkDiLqSH3hjQ4hDht8n2HAnI93i4LOXuktW6ph7m6bY6
m39Syvtr/4ocCU76wgSf1Odgwh34pxuNgIIrgD2Z8bTcEeTz5ZDDauvO9L/LKuNu
SaIZcUjCgrSJDYZgmaXGYSS5dNV8Tc6WinhDG5KbPd9BEkSQfuhlNlNgLWxNyjR9
EnCfy9L2egiMPpvDNfFz/wwQau9FPwn778cpINW5Xj1iJfcwYvEI+V9Rbpm9uGrX
CiNnwVX203wzwLtI2ixOgOOVRbM0am5UdAAn0itj+wwQ2ZqNLOZXvq5hF7p9YNU0
7fxZKqfjmLsGNaCQpdiinonLZUKSl1dlzI/UXaQIFZ9BNeT7Jl79pv8jIbVhlKCn
b9BCjfWrzUDWkj+3dYykiiCoMZb7lRdAv2M5lrOLXJtkeyYT7GbI+pdlKcs299xd
8sb7lIVtl6ZUcI61vZI8sHQpR/VPrimwAvpKkwgOZ05WZqhHyvPZbimW9bihRG0T
zcr9fVGrttva7ZZI7vpTMomzXFgUgVN7rjwmkQSIvX4qVhl24jAzNQb67b56eKJZ
HR34typSjcEQHT1FMuhH1mdUrgcahqCoF7wiN2164oOzsbJ7pCt6zFQtncmk0xce
MicBxYcOkoxfrjgWZ+8z9IuRkUaJ7dXmIa1499V5PxK/RqYMe/szKIluZPKnVPJj
zvmFKo4djYwHtyVz32C4bHly0qBcbyqenacbmWZvCsLKt7aTbRhqTjCF/zbZgLpv
IKRtpYT6Ak4sAGTK4qnMbMrHfN15jQKaOtUCvdWqK4PDvyB2iWi2GpjOQ8dzb//K
+gydOtc4s+IXPbIMTzOTZ4UZw0YXAK0zOeSrzGKN0rinV/nzsoaRLQrjx2FCquKJ
kSTqTlfSaPYDUqE9Vxq9M26DzItkkUZKltCsG5mL9cq59xOoGNqnIsdgQfiM8iNo
JZ8Xam82Edxtt6uXBt0Nly2PilsvVXeOcyZuDHTn9YKSW2Uv10rkloH42ehim6GF
5XHwvwwm/cCBTrabjAoFjvjSMqjbla4yM4dTDGPUs/JaMeRi4AiaXP5wX2HQ2lpN
Hk3i9vQGwc5+kp2fQTZ6c7tLYydTZDbOKQenjkO0O17WkN5DNtcld9HbYgZ5tcYK
EgiAIpdqA7bMBxwjw2RV/ZLUncYskQ9KY5GMpDFWkLOOafvlj9uXpjpNM/Gxogzj
KGblkfTVA8P/FTvHfKViWcjsJvyX5xgVZV8is5bVDkrm/MJrcOI8Wyi4y7gFNZbp
6VHUnIzDnduli2IFwQcDkXBQ6bJgcs4/167sRFEhqaza3iPchuQ3NKQI3d2uXos9
+qBclfkwN/TpyqIU1xNPUEnAVpT2pBfcpeXUzJhq+fExtkK1hZVu7xqjUTiSbgF8
9CaTDa3OomB1dn8a2AczCpsyR9QKFg6aRCupdErgUslPe2Pbi9FK3ePXvqMojVFE
L+unaQ5dudpkLCBZdBkeA8SusFAMWswGGYohbbZpMgTwieh5SbWEEKRsggraW8di
8KLaOtMVXnfVf36j/8ThoxAwlppvndyvtoKwi5CwYzq+tkLJODPx7WhWPDcGFzeH
GnT0D+xkUPUNbkXfza4e6WoArppHWQoOig898PAWZ0WpoflXRWdj/n49YP6cYSsp
+kKeNJZhfaW9guvvThHmsqTVArUXkfHJw9aqmktB5fb9JLPKTR65VmTsFXDdkO6y
OBzxz77z22g/HPM9O8v9ZBC8d6bbPBzFkA9xmp82fgaFFypYd7pNzZBfzuozSTKE
KQXWqoWwcY2kxZVi7HlWd/xOR6dSJXBHDK5rjGRV77qi+IAXo7gwECc3StCMRmlq
X6dcT9V2oAzduLRc/HChQYtb797sJeAI+RaZfcU30mz+zalfKE3DLIqXQalUKv/V
26LF8AoXYp2y3NyIi3Sb4Gnd9f9aytdbXb2o3OjMcsg2ekP3kwXhBo8Rb6scSLau
EDSeqG9YcSeIDA7UBCgizkuGmpBe/RsHtinferTOOSJiyTw8IG0wBjD7+0xOxgVC
E3V1FyOIsvX9zDWUdJcYOQnu1oXx6vgj4KLFV0FihxshsxNPU2wv7dbNrKJcTDVX
26eEiwm1Bd+D7lAC9wBZD8QSvQK6K8nuv0VlGbzPYMk0rUAo5KxgY4q0XT4nWy/Y
KGB6jsIxIbNVAv0LjLTifxH04NYTZKjUqDeS6L9WcEOuxQvIDPAe28mNx630DGlC
8z2LdID0cGAgBjf5qrAWBFFWVSfAq8WNrk86rnohXvXTxosBaK9xF7sngQnyMuhb
j8gexwPv6J4xR0ubFS23EyCWdho/TdrO2vb1oLvN6y+Gpw7ZFxXrhQIATotrjlwI
+t4ipldvV+MpfBZIHBThqJwkSuVZn7HDHF/6tfawAHRhK9BFZdyf/N3gKLgTcPIc
DuFJ8JgFFrVxT94B0w6vYLxJTeDAEoCGu4BIKgWTVsbHwLbYf6j+Lz52aPtaPzgw
sFMnI+T9TjoSQRCP2bGgnuJvxq2ZKP5d3EdRr8anxq/39U2uyRrHFvHk7hlHJ9hA
kZd1WAg4kwgn2h32O7TsjbquRJNZy/b8KXiiJK3GdJ3h4o56c/2x7kHQLP27/knq
WIbtHRwulXFvg4TOY7CswtPIbiOyYXbLma6nc8yIJKhuhGJh0TVuenZyNJQV901C
d7+rqkeoRjb+Tu26rLXsg+gmr3ZQIuJJ9w62p75D0XXSmlToArbELW8m7VUCp3hl
JQq8MEqiKahxv0wAsUGxQp3SmzlzQZgc5J0si9HnNRm2e4iPrdNrBwi5qYwK6WBb
5sUbZOLqVDGzzPv69GbpINyuhOaAAgPhTYvm7rfkR18LoMfvEl4l7errWqDp42B7
9kSOVnjL0b+tGjxMV+jWnATBA+xnYKhn5v6HvWxy2Dkc+P0AhKP9K5qdN+dcAJtg
hxmPmfSucwrs5c1LQH8i2yevur1W8TYHAc9eL+g3yOAzE2LGIemJTAdRP1+aMGAU
0djFBX5GCc4nNGuvGzNDh9O88t26DdskPZkeVOKztWbVEw7YUe72Hr4LGBZKMPNi
Y6bp0+TxUVjUVThbUjWVHpbSczqiAE9diuuL4qzXLM7yd9LcVlx23uVq0NWq5da+
BZ0NHzt8W7ysTUcZGpUCLW6NRQG4mGMeayGr94Pf13L8ZwwtguLvfOBk40Iged7M
i8i+M6a4E4drh5DtdJXfW7TuTejPe+uhzoopWNJTtkRdNfi49VXhUlqfgdbRi5lv
Ive33NW8HMSanbhIQL9MipdedMC25PS50+5IAcNqnReLEyViyPUVCxDC+fUIG353
cLDsjNOPMGn4l2VuIE8ve4S+cA0epQKdl/FokACC5jKLFuRhVtodZHyJDKnEQPnA
jRr9IJj4wVY9PoZJiBUt2U2HMHdRgjJNHoLohHL6WFUhfPE8BCuUVPzhv6iircDj
mRL+7rYucj2iKMLGCF4qKA6s8iANxeZjrw8lPZLeVC8c8dlt2ygVY/tZjeUTNXVg
frA5+9JDN0UTFZc0KYCsVGMOaKXr/LzKm92fLivex1SOjGaSc641RzXCqsBcIcAr
hnmlzSDzIlAfBpM7+AQq7hAq4CTtpUYEfw3GMqCoo5z0rLMrMq1FyQOTdwmtOx0T
/l+pmW51lB77CuSzzFqHQ0zMfDWIRxa7wS0mrfaU9rxeedCpk6saO7CWeYGCCcsC
LmOqP/sdsClddRXRxsGmcyB2oUuZBX2yeDGTt0hcz2parMBI74k3pJ6WhHJF8/Xu
JeK94oNtVPqUSqxXdXvdtfygE9O5LCV1BPaboDgH0qfaN8QMoUJzYyTS8BNbX7zx
A96o7W6xIEA4dT02/SiStGWU+tmmQeSZAlEpxtmg9eIcfh7YWfXkl/OQI3c6sOQI
wK9M//qcbX6rYlR8KVQgVhcZYWZBbVoIrzoyUz2onKWCLvV/GbXQocnzKQdSYpxR
OZ5+lj93jnwfSGs11OoiX+deBqXN2vTyblO7lcSqJ53wvAPGTMWkVGXMzmfG3Yge
mp5weW7iV6futU2IVQye9yg5nK34M/P47vSuWqDqRjdspmHbYKaKHNGGGzHp/N8R
61fP7+7xhTysiNLIIaVXuisY8opIk56adKxRrYh+J3TxgHu1HXvzo7l9w2dBhyVR
bBTzvEC8qFrEQS2GaUCwQN3Uz30oFXiwsaXs49tGjOJrXvFO1NDPb0RCtqNOhysM
y95aT0zMkWmEDR/dSWt85T5IdcLsOOYdReF26SU0urmQl5ThZgysfl4XR0tqu2pe
pojzOxpVJ7vu7IVz4y3n4zSMPMYVKAYtu1CSpXLFpmqiTtuUfH6z5cxlRpGHtPIx
IuERALZHzaG53Fh3nzJ+jG5LnQsh7HpFGms1/X5oTPrYoKUcxScLiSTb9tczIzCf
IcRkIt/PI/l8UU0u6l452tJis42BKScayZhiYQGCLCOMnP9+s2EpZPrvNG+mFURx
BfSBK1XB5d0q/Clrjsz0hUVf1ijFOVNq1FWgPSQEtEBuuWP8uN1s+8/Gw1MiHdCm
jCWpB9BJFjcZAdk4RtP+TM21UGtqiMpc5xdzxv93GjwUcuVZUH3MJ8OgrxeQ8W3a
7xb6I4uaS9ufjmJJQG+URT0NmZcegMmXrY7mM8Mp+nngicChxM9UtgQ4fN1cj28F
Jm+DdDR/wAcxWqtupE4bVcfbj/76mZRoNi6YHfCpg3suR2M3VFG5YXgBZBx4IX7e
UA+dnst6/UkLk1/fu4c/57UrKde7wYm1gCjxN6kiuwlMvbmd/kC4ptkpKseJpkxr
iEhs4ObDds/rAjq0pXRey/k6HvzrtIak3oexedkQPf6LPNWJ46GMKCWnioo/C2KB
uRsBXm6DIqCzps3HFjsDHje91gRLqz691bd52H+LCe5NvCumZC0TnoHNbYo0Wo5W
yeO2bFES9m55doqfPEy8/YKvSSk2Dwjtbkc5+s2R3C/9fRwJw2zIQncSww1lw0ol
np2tKH7gXP0CKIjqbFKUBJIMFSU0SHJYJo0LxJd3IdJXCs2zzOZqHp0dNUkLtKt7
UiUq0IggAruOXj+cCTx/hrKO7JanwzK8T/N0o9pzzzjCoEmDXtvvJNUVO1/5Kgev
8OJdh+q+7E8QUut0yNxfpe+DIBrNGlGpkUAkPsUb5RSbow+IqmxZZuZEzOSYyWQ3
C672YsLW8b7o2/88RtxgJ2IejdcnkpRpCPMPSe6t0SXMmLNZiG0RB/d/ObLozzzJ
BET1Sn6G+iM+NctWOBH+JHTpifzNcijJB0uq1ZimSRDGmggeKAfudNBeSBV0w4ww
QokZTaXPPlf+f4JpNBMWLL6s6wob0+6P6+qEY0cg4/qjJ2ELCV5NLwg+skL8jz42
9OUVfqfgz2h8g867oLWtsDI35qQxoc5mRhIaz62VBEDs2FVT8HQ4VXy8FT1iN5g5
kQ2eWDSQwPP0P4eF9MXDH+/1a52ah0QY+eNqqm6+LnwwqXwaiNU6EOUMO5+4m9vA
rsd8Jo9RdxHMX3mai3lmIKtoCUgQQIfUqAXfM4T1gKido7m+ZBwLycnYZ+qcji5N
RNaW4YwcbSfS7f9XyPNzS79KXfw2GfNl5hDimHazl1qbDkXeWwH2vDbv9XH6OeP1
PBYFQr6SZiLw2y7X/YV8RGN36mAHx1PQaWjEuYJym0fdBCLY/jxhUvN4OoxUbR8j
dj4B0L0NDE5wHU9sGdWYZ3CZAAltql9T7Fma/gr0aShPbJPox0b6CQywrOQThBxQ
lYjDwuG0qyWCX5W+KlGZA3+hPatA/4hkPs5IZuox0ZHftzwXjG3WYYGiv3Ip/NpQ
2f6J7DvEnlL6W+PeWHbKtd1AtoMjngrYvFfxQLbiAD5Qz3+XlfKmh1T0uJ055W+U
0v3gFQ9orp53ISvzaOiabs8NaEYPBddsd6Wn7yIP4/kHfefDgtMfuYo1JGfzo9fp
/F2qPwxDryVLkSVmfxdl8ZPd0BUFKL6eFgMN+kP/VeOYx4FuPwus+8HS8Bf5vnPT
ixZp843TbIDjMyEXL8Pvklns2cvBoQY8GtoBsjkVDaw4PTQbGP9QJlqxuBh0KWIk
YfeFjLQfaXWagjPV5Lvb17g/txMmlC0GqBoPmiIU9Mf0PP5qE74YJUHjXKKEEgT6
f+aP+SfM02wKDN7gREjsdghcBAtb5BEs4Cjn/cEkLkGDBPeUo2CP7ODxfaH+lJ1w
2Mz98UcNiiNTNh9/k/m2ehZpuLP/KYqYMVvXpWVY4dS1wAb+G9hOT+j1xstKbnGo
fxQLlGrfEqUvp0PkPIzLyU4B/dnFxW2QCyQJdIRjQ0i4WrtqsCnvLmS4clBsgfRi
yshnyGyQRm8iyf90PVE2+dT0/hQB9G+VyDjb8ehpTInRgh54ZRDN1ww0fVI8k11/
OQ+yC8ZKSZ9ukJwUCUQZblTzO/8CLF7LHR7ZFUKw8+pzzDA4IpVkbxbCUaIJVJ1G
PeeoWiQegsEBzz5m8xUkQcpKAB5mhrxK2lYF1g/BvRkRiy2dRQjfSk5lTwvKkalh
f7LIL8OPyJ25uOVgZTV0Wc7z7NKZI/Bj5Ry3ZWT01fLxLtz00Sg7iUp/oZNoabGC
yTsDsvOBHQoGKv/LPrdxKIfwvL6uEGjjFPzi19YEYHAY+5+mLZctR0+a7VBUgkxw
Jhu6Kno73+Z5X10kFoAIM2ANQSJqGve4ys/ldsLZNZDNgIYpE1luh5PWo8w9Jkn8
cPkjprBlw5RLzNNJwhb8dTaP5/v967Ftb9VhIQjPA4w0mS/+e0/MbJL9GAJnVUae
IFc1Zqaf2zaIYGnDScss1jk//UEo9fdVpjlFaDpf3Cdt22lNoUMjwsiM3DY4dD5H
h1ya0oFZXt0gyd1dzT/dtDEdMGCQSzr+5Qicf3EznIwyvsiaem6FPCJpM3glWlU5
//xsNPFd3RPi9Hr0W/iCzWv2PFLzUu/cEaEuJ2+xVxpQ8EymOK56aocVOCPEsKMj
AP7Fsjrtn1rFSbzKWouZ1fJsqJYXfx1GPosI1w11y4QoKwkRy8lCOaHKbkmMf0J4
jUHTq7sb6wCZUq90iLvFxQMfZTOLUy/VSg1ynjvYdhjunikHb5eFqmtLnbfFP36E
kzR+A8PfHVde52/Jn2JWCGx6sVMWshdEkcuafQHhuIK/d4fnPNEJZ0zEeZjBfLYb
N89SRt2NA1+Jour4oq2D3qkw0bLATsnAXlQ+hvr3STQ7fnl/W16mcfbgQoqi7x1n
mPSEPjEv82WiaUWtBfYfzLEua0w0EmDJWxt2e7s+zacAucPNx2SXYoUvDbr1HDhd
jK0Z9DhwblHb8apEJ+hmL5S13aBtQy63oLLcOv302qHlWqcN+7tvcUKnZMr74zLm
vUooedRkNB/SlXpPmR1/TEdxL1J8TkBXeZI74BJy2aycheqKvWM+ckePTQ7g5FoL
vVe+7N3XN9LxE2Ioc7cYVpM1SB9neCcF+ZL5461MdpdhwFEEX3k6PPJE1Ux7ve2d
Yn57rot88Q2+H2pjJegsJTxXCRIuhGYueF14eH1AxcGq/+xU30xYvMyrx5gT0evW
kzYgzMEpfINuSgVrYIvKMAOD41Y+WeKWo1ybBXKqm7DABcWaEriZ5kG/TiUTOAHQ
4QVIMCtUsdOQ2lftPHF8WZYODG+ch3scCFCxw5hq9I/gY4K1elZz/UP8ckAD1Vrx
q9UJqxatSp4SPmfHNKf5kGtoY0g3tqVZuM6seEMmP3CRSJ64EceffV0N3WRzMpdc
f+cqTFdcCEB7b/Ud3gOMEgb74QiGZa7cc+jJBTf9XHnCNeEr5GvMrinFhbhK1bWa
t+X0X2yv5sm/3lhuD3e6e6UixCrQKWGBIWeVgm5G5jfjru1LTdqXRd3iBFc+cAFN
bta1WXV88w0i1R+po6TnEPNzBHTdfE+GVe6SVR0Sh1JZBcomCU8dQ3FEzUZsigmz
LtNOde5oKuikexymjy9bC+rmevXBwwiTWAEpdy64x1ChCE9yw2Ox8WI8aGRcIa9W
hqLYwWrNk3KHVLhAmugolAmldjtTf88Z7rd6aHCW0qcBL2a+GwgPncmCChiUqKUw
fJAHY7jiF/jUQF0DvSe5xdZoeP0BfZLs84xiXT0q87ANrbJXxgTIlSyqjzYSUZAY
/b6r7K7wFIXaXIq36QHQfy2kFLf2BECSKFrCEzlxIAlZQoVn4eRc9WU7h5EYGIvC
QKXnwRGmKdfghQuOIixW9WjQQ6ECx687aouRD/LkmGWF7/pWOneSyEhLYlaiSUhZ
Y/M1Oa7MILlH1wyRaoNSr/EuQSd80jid7p8MrylxxsksVi0yX303ktX2JWOzQazR
hOml1Vyi65J1KbEkCL8MaA1Lin2f3s++pZSI9fUNUM+lxrUdFwh1BvTGkR6reKhA
oWpcSWpySO1YUUL1anyL7Pv5SzRUJ8YzR1xsUL/3ffJjOekWXGr4dzdMCE24iQt3
iJJ0axgBbNbE3iIjhHSY33HKYiisgfW+LbAT3/eqM1VYG3ievk1g80i/vkIuHzRR
RhtxT/EQVKRT+xrH2dNJb1TVukeFK3f8CX81W3hize/1HfzpUPM2kWneA2EGXUmc
EN2qAIbOHd5ZOV5PvlQvu/v7dLpbvqK2iqo84QC7+v2jPiUWXavw8P94BJ82uHXb
ZyjRoldnnmiC4Ezy40VkHRqnb7UH4JEcHVUKoa07guVO6g9FofY+GUYP3qXvXaOG
23psmfH5jroMwXPkIU9qv56H7EWTbVsSDEF+SkpQETPVZgJX2pnxURUK8z0HYKSE
UEsPdxTyju2BQzSwHtbPDYJsL8BQnVG1s9JCOCEv3QR+R5DrhB72YzGFD6RKVvrG
kdlfdynCHbN6EjbqgRNLeVhTOIihA9UnqHpcVjJ0ZgEDX9DkzBxxAMleImi0I2qG
6ijDxLuGhJUIqvuBSU4H2GXr1GOCmmLxhx9hi+r3CHSSbvVbGfVFTeU/grTh4hIK
eiStQ0GH7jg271s/HiZLkS3qc/Hfdwu7O20RbVOhs6jTkxX4FtWscLtPTcKd/aZQ
heio9CiZmHk8M3o5Td7LrCuo9uoeCE+WoQeaCx/uBV6iNbqnsa1HiNOU9uZIrSau
95nHmt8+XAEYWYCYOZPRG40JOd34iZJhNNO/VuIvUOa2t5xbeSq/fNJSxvTA2Me9
Datj4WPaw51BfKgIifJGP89X4JzOrMMUmdpITVElHhPH//swCZNQGv8gZXLVt+iO
BaiRgC44rPj/uKklyBB2WWrJM8VNg0L25zX2VJgTiZufAL8K9KwCcalTzCOsKDLG
bvYYFCOW8Xq/k9VjpKrcUL2PTmHZTWhm9sNW9sI5TF+DHjK8gBb82ddg/hm9Jyqj
Ec5SeHNxAapBVBrniT6omWdG+f3jUvBDOFeuYesh3A2MZ3aVMCeISEDQNuRzZPjj
Ln/54Sm7SBCfQs8LBaSvj8QR1c1ExJzDnrkstGPgwy1765e1xH+Et58/OvvJEnBS
+LI1OFlZJ2bebDC+AX7aATMG01ByYu4tqddD2foLk5I/SEckpQvq4cA2KAvQxVvY
ULentE48BwxAVTSmHCAfoNoU+si4PCcB+9GQdnmm+Ia2HOtxH57hY7stGtXiTkOD
hugOD0DLfPrEBw9YVly59snB8vAf476e6BJwoO+IetOIAJiQLu7+6J+BB1n0pFxb
71vudLYmfEGcNYIQra/jLVrjSVXFZcVBIrj4K7B90ocKKdG7RJUdhxWtNEu3G7Vx
z4+WFV7ZTWJnPlaEwze7H11ECxaC3BVq9oQjxJo/m5Djl20xmdnBHI3huEnL3CzK
uWTOBD8KKT6d3XW58/L59E6vxdGjNGz8QT1stXspdVK2p2lLvTxziNk6m300t7ZD
3VHbMdoDgGuASUIQqshVWr7EM0U99J4q8U0Sl8TehLcPpxkYEQpOlgCTsJttoQAM
QzCM6gEn+39Zgjb1LPVwDLstcISJ0auCcPu3RVTLs6fyLQZOAOuhDk6nEy0QP1Am
a9uUdHC2imczVDixAsUg+zpGPffQMvMoMfdj+vcn1uMR7zcjtXfVi+44AOhtUfNR
ruTW7OcEI9qcalB6AaxpsiklfMQcvdACdVX/uhZOkxGrh7SNq4WId27CoretOlws
DNaqW2lkUWXgcZcY9ljBW7b9dvCz83xfMsv3RSNsgUi6PFV7nFnqiI9TgAxtW1mK
bQV2E7bfUmQcL8f+zmjizvvbR4mHrnyBtr0w8RQMBJ7OlW5iNr17pn3Og59q2FLA
efz6h1IaXVy5icXri2UPBzNnaOMVXH6ppDeQsfngjvPuHceHGJlZCARLxxJMoFjX
2SHvoHe8XSOJvL62MyyXTtx9Ol13ZvPL8z3PRbxzXuqrHUpntd/YxIMFRwaVF0yE
6cY9w4Qga77UyR6skfNIoXCX0qIP6ET0/QXp1S8H1nrGwncDqJLMSqWvpPUxM0tB
PQFVlizQMq0TZG6RMiibKGDhDoBDpuvkFX4yL9vw0SbN44kiPSpSBIPB8DgtKdyG
gmKc8Fwsu5cJ9zk0HcUzBl9RvoqLqpS2iptlVLUrnxvYQnB2gyLcXr4hFqhv9Cdq
m2YuqDKqhE+YbEg2x+xkdAiNw9vpmItUtJSSy392aEp78kqmLyY9B5DOXibnBK/E
I5CFdgu/M3wnqivOucL59ziUZIqD4jAY1ALolhqMHmHimROoJ+vbgw6/5mFx7+Y/
l5TSNmXdvC4BFpApCnb9IqMfQDOou3Btr4w5P5fvftWft9Drya2R4qMm5OQzOGuD
Op149czNsVOn/upAXeBXCwc10vh/BD0H0nJOhJri8vUunp3mwUr77eKDY3w66X0s
PDWTJ+aPTUOfdo8Gi1caFMPbQFrWjiejdhHv4Vmykv2iyyHJO9Tjbs1maU91sqCZ
uVGYonhcOQYYdXPVCuEGAqQGZBcxnp6dMtnJed96/CUhtJAjLT5iLdjzUUmEvJ+T
aGYIQKipVrulrkHZNPbBsbkSJNESNmrZEHddKv0b8dzfOhK3YR2UC4lK0zvROW5L
FLi3C6IGuBSmbhlySUA9V/kX06vbddD488XWZpYr03f9F97r4PyuPMGVEPb4l/jE
mYyTBdMMzlDK8Nntm5L1KtYqMxILEeOe1ng3bj9iuGnmARk5nNn6tXXbPdLuAEl4
IpSFF0u7TSZhcfu9za1EubU7Fj9rN/EqaQ861WQnjEVzjILfNuwQ6/kWPqDIAvZg
2L5LaLDX+Bz+H7jT3fMnmoNpenOsLIKDP4/Lbc0eIz5T5Zy3KeGVrtd0iYq2SEYx
od3f3t29hE3AICWPqaGYe2nHH20tfQsN/9ghqKDqVaejof+cRAj+piEP9Ku1TMUC
oVtyB1WrDOsEAq3DcbNYlgXiuG5O3YLm7WH7Wc6c5Q9shrfG2ah81vwYzN98X53o
XpZSckwFtyDKhOhTeWSEMiw3cMdKWhuhpLtvehG77zzQZrmua/8LX0vJB9sAYFt+
zl9dYl2lw4w5Du1P/VSwysnHP/1Bohe0T7wqB79JFn3+objL2XKLx9EdiqeABIcE
Zd3H12qmF/Sduqycg083QXx56U6mo5vS+BoTveLKzvtqn40PJI43cjtOHVnCtdtA
2wcLV5xInO2+jyulOP0d+xcLISIPta+iNSvjntl6hcN54nZnQCQ26hdmVAHBWw9l
q6Ni1f0hMKG7GHjCEdKKQmGcTMLpQcy46eVmJ3PBIme8BDZSjoRtb49cmKSz6wb/
JvvVufLt6cysrzlweCujavU3K+DYGqBwWNkQn6VEk7fpSY8yuNVnUfdP4T0XIGoz
FuVE7vNLYxzf/5LyDLtnPzUFqaZRasyIWD4G0GS1J/mg/bBoVOHsdx8haYImuLDm
1Z9vbRGBwByb5CncmCvA7XRvPLXG3hlYCthLC5wKdAKR6hFb9iKPxPDxRy1zL5et
1SQ6jGYupxUYVdC2wANQ7vHWAHUtwwrkeaqjh51BE8w+Bj9NL7jdVk3DqRKg8yxJ
GMz2jooeh73XzcDAzimu/IfCRahofUGqpQqffZlAOJarrIXBIgTMbZsRlbf0/cqu
vDnYiitGyDrofDl3iCzMuuvBVLSf+XoVEdQckaB5VtWJq2RHTGKOpnccX6i2ZFwe
Adz5djQRHtL8HWjEKT/JUgYQumBCG14ilhN7tS5ryL2i/eO54EuDfNLj9+t8NKms
USF6u+VGhHnnAFWGoDEyTGKq4aCJ/dQuaXiJuOzFDeAcxgMFXUWW0eZ7SiXQrpUC
5XhW4ZbiCtGezE3FvYxmMgM36KgoQPX/RATQKN/WANpGEYQVLIYcE7C8RpoMbLJv
s4tL/F0KzsBoVH0jdWvh/aK1RP4xpoQqfsfUz4ZGQAWI7bXPkTYHl86wAOwCpuzz
bub9MYYhTt/jOZWDPQGM3tPzcGtcqXS3KqPy94nQ0UrVKwys8bLZOgBC2AwKOEUZ
AAMfOR1tBYLKHAUQmKAcffkeLMN2lx3+IqUELnOAeZhqRzLRPla7/yIIZnBBqKa/
DpZvCEuueD5pBH6+oKAzG4IymdnKnu/51qdGjhzIYZGPKgK+0xw6K9Cjn+fEU2FA
Q+2z58pZzDAVaOmOir72ge55283nod5laIRF8yHwcMzFRAvAg2W8KaoW/iWp5ohg
/qYE+2z3Ju4Luuk/0fQEaz/u09QTWIcVjyXljTuNRK8BHVuX5bnHi9RQtbRfNf/9
zw7juID5SVscTajfwQhbXboVa5XuOD/B1X6i2D++sl68w76vyvSNt5uafEUsXqJy
4ulVaLX1ZfAwN8j2kfUgUPRnxJqtqXhH1rB2qPFY7UfPMFBA19MoJ7y9whFBFleH
6293x6Xe+P82OAOB60jz9tVlPH70m9tORGwlscn9Jxqn9Ff5KtWhJ2FBURY78aoB
RhhMWxPjNQLEwozSE/GeJeR65HMoj4Oh8hTI0JqJyNkhqPvT3ssy3niAPnUFsCeC
vwqdWcKjDIVZv1AOB1wJuItx+w7zx7OEq42uSN950l2UYYMGcCUwPfca94EemPxF
L7wn1Ml+cg+1ISpt+lXazFbu4ZokEEfp/4Ah4YdgZjnI5kV5yw8RvyVY0dkxp9Fa
eLNsmrGkJDXR7jxkTiaj0mVeFWLZ59Oghk6wajpaSkAu3fsTMlERhxn/0uKasKWU
sdkdFdQjQyKvKmYJa3QUiBqE2le5yPzhLgqqa48HmBvWrEcSxs/zUIlWORFHRfY5
X7oGf11rgNvO/Rle6kHlOSUG7p2XWVQkj48n8T94qwbQuEC7mq+MRpoqFumUcCtD
8MdKCrWtXjQgF7qWmVniWiKyO5zxyrpjlDtmIWnXlYYq3nf6BpVayXDY1y84Q4Xp
tGE0/qZRJ4WMYmhqa63Zmu3tKs8Wk0WnZoRXbD6YVqWmMl1zDtyAE/uf3cdW1N1T
eu+Eki1L1XPjZyxE+RTOV2ggc2wF9VQgJtzs8t8DQTfhkvhwcrJra2V/miAahyBV
Oq9BlhilFCTL6+ae4bOasFgTi5Wl1dv1j5oVn2YyJE0k1on/NsO9WRUa4IU5B0z8
h0wICLMGWzo6tTxlg8uR3CeI7OljZBiLSSRVoSgIh5wqJR3ayO6O1Ukzexg6qljo
2fh7HlIW+h0ceC0Eu6CHDHkDR89/UysF9kmydCqWP+TIBteLkvm44CC4cMGosRUZ
3xirg809QqnyAYpYdAARgkLYWui/aPvZB8G4WgNGoU4yE1rxNdQlL9IcXH4RnlqC
ObJs5NLkSaGt7KhC717hZwm0IoPFLJ0OtjYjAOIp9wfIqJLzrVpke4uuAd/3wIfJ
U7qjHCEwiIApPj5xaPLeDWSubMF8fVSqJ49JwWw6j2HKkmrbNaG+yYgOiCKI7beU
9ZACBEyxExUHuiPsw392TjhsZvlVrkN+/wU3BWUrEn+xCIozVcW60HkM8dLKduaq
Ts6mvbmN2+f9aXQ1Pz4amSRj8j7NaQ+UncUP0TKpqeXNbC4ZcVAlYBUzIxDCuQ48
5eKSAtG+UwC4dsGnDw8IXgoLp+9OaDYg3GPZwyyvR7cjjjctA5HBKEWP5NJA+Uf8
pRUooNZYv3HT6k90mVcBll8GQBwIt/p8cRzzyZ6anrpjy4bKeElPZgr3SX2Ui/dd
AAZ1wNQhzu8/TZ12u+wVs1avkJbrxSxek3GM+rBmH6D+LGpeZuSzKo+1j6qL+9es
/NjZySJ/8I7KqlCeG72+aP7uTVm+rjjPNi/05Vm9Lxn0Vk2sz1DC35n/Yicxdder
VqulwoXHXA6eyxfTzfpAc141Z6ST8i4s2pQZdUVfFlOo5RH8h5pxSP4Pqkmo5ynJ
1XS2imj77dyYhDDIGl7wtJIpQtKpcVQhhQLbNXOpFqzKcb7C0i4AWdgK18tbjc5o
/yij4jmXtvEFD5rbiZES3HeoFGli3pT2Sq0aMcOO5KFRVWAyufb4nNec2eEmY0br
+cLOQBqkdi7a0zfycY5g1ftIXmXKU5WzJuIpECNgB/V2ipOQZVJB0Li+R79AATfz
BvbdlXc0vtxwr8xBhyqTd3m6yvF9BdSMYNDwQAA0Wqmsl0KIVRlc2dKg2/bIxlr/
S0meG+sUtFfCwf+3fkgSv5r5X9TM3Qwl15RRMqIM3ogDpdYDzgAorw8cg4N2tGoA
1Em3PFfX/TB/5wEw4wgyp5pVr64KCwU3xlPKsI1nkYSX+P5y5cnaRtcPigok24D6
VHB9J7lLAJMVhH0Y5fNqjItMz6HQBNN3O96dOZQAJi4kDxrusmio8jlxlIUospDX
+v7VGYoISbkiJ5amQYfi4pSNI8IJkW/HnfXO6zCpk/v2a8pX8lxZ4GlHH4ulv6Zs
e0dou9lEyGwBXUmHM7or88Hy0XdisZsamvg+dP9bSwoeD5jAVCOZZdpLWsVR97TX
bqNhfGYoOP/KaTvRYqjNS4AuFz/ee/gbHcC0dV6NE8e5x7oRsydy0Ex+r0OMhe5/
LTyoRlqtViRYe310oItmG3nhTYkBu2uGtNQXKVmB7W7gFbpq95uM/xbyxf3BU7z3
KR+BGFcrMWQy3aUNcOKlD/8MA5N32KdZCx2qqoWM2YT6XgHmbWGzvOVvoeg/R9rr
b3Z9NtjVIiqmj81TSBGNfBFxA2CIhj/aRW+rauZg0Jv57597cKAfhNWrGzx6QbCZ
JK2qh1O3s71vRev7sVf5HtE7KzCbz5BIVLBcDsk9jmdpKRruxttcOxK7vWhS3nvL
cDriaFR/fGSAGIdCUhPzceZxPiJZGo/U+QPXefPnc3539mcKskKwgXMs4A3L+j5w
Z1gaGERFR24QZMkB1BTOobP9kTNTjcjxpO2MjIfFWkU09OgYirmQVZOApTz6DBqU
oqbyaEI6aOiyyP6f8VwVhA0l4KjbRaih26iO9cSY7Hj8JvTcKUpl9yrcyT1bWuWa
9cRzJ+r/ugv2Gol7+O2eAtzfUehIa3S8Ga//cStOyImKfYI825SCNx2WR9gZIXP2
++t3n1SpsQDnyfBlRuST3xZx1rJsXNZrIx77WwJO91DB7E/rquBlkp5SuKMu6dXn
3XYrCS/AIzWEEmjmnh/u5HWlJJX9YoplwjKXMH2rFT3wgvJ7h+rrM3dtf3DDWnVI
H8zJhHTdaF0dQyGdrvu4rrqWTOOdjXBYQZgnQHKDV0pS79TqM7H4U0FsINwVUJwd
8Nabx9Ttd5q32x5xrt93SCLezyIKlCW31GCoVPVs/m/jdYM86u303wKFVSK6gCFQ
LNyfg5A/sBBuc6DQkoZvQYUuDEdassci5/nBcBQcmeUZJLy9aZpRMR+qfovfS3TY
17jeSYOf8ZQhL77qft+D4y6W0FKECvM8y3b09hYpFpFE+PhAf+t5CKJPSohg+5Yt
fEufEzJL1JV45kZ/uWmJUUT6NbiGtcmU8aJzq08dirr/ITa5YB4I8gPhEr1gnICV
ti1ZEiqaVz4MpJ4cJgrfM6Q40/Mhog2wTU5pmZiY8c26ISJEn6RVV1DqXMN4ZQyI
juS8315xB4APgWkYC+j7gw==
`protect end_protected