`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79I8iZ3MaMca/r3UWOgJzbEb
4ka0j9adKevpK05p/oCzxAS33moAGJjJkT37KVTM5vas8mX7VkqSjFJMYUl+fka4
WRdIC/iPul/FdUMudb7ykTQPwTQexEDOyTnkdezvbDnTUx/+B6SBSj+oLpKD8v9o
VklXggyQZYIK8DBELA+HDao1h3ATNRyUeeosk2BaS5hbmzfLHNHW13fxMalSJ5pg
j9BOXXSWIMyZZQb7e3jBeEV8Vyrptawquod9TdE0pmh4vD6JHSdjjXPv01oq1ija
8Vtv075gmD/fCl70eEHc5tLQPmvuDBpjTzbs9WRFkcYKpSh01UXE3Mf8VZ698xXA
MxFt0iu5//8kdMeR0tb7sUaegdya8jaCuuwmYOg/oxV4WYXr0OPb7R4xUxPA9Av4
4JHY0htC0Jh5LhIBuvD7c6uK30pR3tXV0EG7FAE8qMPcedc65wbXEqyFNpl+oi9S
umRCqmHfdwFMrnWZ0dPBTC+4qZsN43YXeRjtHfWm3vSqkWCECWGoHaO8PaiGDxqb
E2jARP2EisnFE8FXA/vT+3ICq2UXCaly+JYfgeOfXCsQ3Uj2nytuZqrteQKs5l/H
vUXd+iGs/K2JOSPoX5YAlXkV2bYG+f4dvsAdmvQIWtYkKMkhgn+EbS9D/4NXpPrr
hePT4haaGMrpBmlXIAvPhfP5pRZIN0quObULsOhgxosunz2VwJRm4svWnAEfZidk
dSC2Jd92ci0uLp6ElXq5UsrdmDd3vGoRqHnILQLHsd/NgPV785pHk3JEpQb3sr33
/HAMIdVv3y3BqIpS3k3fIFQU3B+nX94vTZ9t1ELjWbrCdOWzTZYlPrBIft/TWIkA
026N9/MunkclKm+nUU87YRD0WjqlEIca7lTIsGlVh6LPWgcyyB6HTKbwNBvcgCIZ
kEl0GWvYIPFv3zpPeP7qp4QWONFH2rEggheD41qrN+AQe+ks4bRM3IYu0Q9XvCRL
297JLkkOs4j6jZj7xuwrnAbfvgIISRKObFtwknrD2oW8rCmisYz3j3uWwnu7+vyh
xgjmHScvnyJ8zz2UgZp3ugmAm0OnGLK4QprozNvHQZj093x5uY06V2U8LKQO408t
Aj7P3horwFaC3p3EBGiekD+BIzhJ383aHSSH/+x3VZYd7+e7AEjtPDkbw5r4mV57
yaS6xkglYFy8CZPvG8UAJKJn4Fzm5JUqqXtXvZZ9e2ETMKoC7ucIC1fl3G5kWAbA
srmrENKW0yMuxz82hBn4aTAdvzRAS4XZpSuOjSc4v7Ehi8JZoOC6+WPMOy/vWoDy
eGbdWEoMz3lhhge96kiESMu0sdOWbe2keLvIDZ5d4pkQquQfJVKEiU0bXA3BYWlv
MWc5FGocAeOKxTYKIUEMXmX45dcF0L1y/3qCNdw8tPN3U7ohw/u2azOoJrGQnxKu
QhF8hiaNs6mpiwq0IinsO7a74OQHZiKCOGgaxwKW89cwal8NPxfHwHjG4KkAcQ3x
3Zu+U/T68IGtpcj8uPLy+1qOmHTFZio0Fvm5ufJ8ew0bUBvzwTpCpID9hkL/XEoV
7LV1af0xBk4ad0I4EANMKvnTqTh6GMWDfjTj7zFanUu27pTz/nm+NCHr2Yc3kNpL
MR8HQDu/7Q8BqO5bPxbsZxkuwekDmdxYvCxvlgwEi8lgh0o4VudhewCmzFyG7cAu
sBQ+8EhxaiL59Ajuj3b0XuWHnN5y4228bdnEGVf30jdafjl73R5yYJJmnrB5uhVk
uW6nAHGBFvQ9cfLO8hg0NlMqeBMjzcy2l5ZgEFyMzWh5wSww0Qqs2G3Eu+/lT34T
4yndlXa+EfIOyGDURbi2nDek5iOOVgGQ5gSnry7thyGQ9Gu4WjbMXtWJZGTOSTHO
Lj+XxuroOweRe7nXLB2wI79QF7zWKEX1DMnZzUD7RWekUm2d28vt/gBuxwtbtbFE
/jcMIFfZHUK9WrAltBogf4IxxbQPjGyiNpOfp/g8AkeP6dZsaEGGpCfOQCTQ58r5
JUSk1j4FkUSPgAhzc1Ek4skspDKYzJ3uD7ipcxOH6mKxZZGaqBxRjoQ5G6L/fGkz
ijpE0zZCKdnxtJ4/5pZrJyTiOvuC5f4ypuMps68GgLRErml0oxF3SjnL82Nwmn6u
GMp+ztXm/5IUtdaj8ngxR53mvdHns6xJ7Bxb0psTB5/1kJd+hgdLwdf5WI/FAHDm
GXr7xJLT5rGfEWiYyRU1TkSTHg9QC5BWuZ9gk9uSaSCsgcAm5n6S1eOkGOcfGgmU
PTHl2I/E7HWqHygtlNDMbLLP0bW8Ezw/JVzUebVwBP+btC9VHK4uxWqI/zEDFf3C
AXBnlG0s1cUzvxKQ5jPlYAMMrEAMktXU2D1SqYncaBj7b2bIooJpMcUF11OaXjr6
OnA8Pk41f0qN9LZdIdta8uWzZ/Zo+YFF9U85NZm3t03hxG6EPuLIJsIPQwJzHX7S
ULlKX6qGdb/c7StuXUU+eFgnaQj7Rl5VMhJfi8pAUlED2U6sMfXhz6QhQ28aR1G0
Gq8Rs28lEgJxf2zGEPtLmkLdNrzqOTD/JYCGj23IZJRriFJkcE0BrWIE+tibR8ZR
N863v3rvkGCfEd+q8wgATXgaN2JT9G64KSHLpu1MN47sNxnxrQ/7u6NQDaEke3+d
fYhu9Rs0RIJp7VSw5gVPt3SUr7GAA3Ngay7XvRPrS3sC0ApDAdSmcA3ThpFIQMgp
xbiEx9ddG3Ib5no2uWnZiJW2rSiLdt/JbIvDtvV8QTA0RgWG2+HXY6jZJHz7JFOl
yUPN/Iv5OEJq5l+Og1ENi2YCv8thkbn+8B9cCJ8rP5UvsYcvLwsYvgjuTsutADki
EUimwCoNOyTTI2CI0LJc1+xdydax9ocA9achp8yj7LFIq0d4mxoR0rh7s3kGy/Xi
dPAZ/6QOlJPPuQaeE2OlruDvv9pqlzvairDdiGFRKGA7EAvTzzNgd/6Xr927VFCA
SZZAIcbKRpX6IcO1IcShXM4H1Dy2Fbcd2gDqA9h2Phc+GzbDiusOwESjmFAebcNP
jbOVokZed3OcYDXTNFN5r9S6Hr4GLVsqsplLlP6/JyTCN1X4kIxFE05VFrdci8a0
DMIteEXTwNf+xGTzK0iH+c0HeBMQHmN2+l7dRcdTCtB6f5VQXqd/D9oumNuJ8lVH
l+UaiCTUgo5ZbcQ8K8n62ZVmCRaX7F55SYEUFBFnKP14HAPKkW4ocuYst8ktNE89
ylJWobhda/Qpra0SYQRzdswCHUa1SOL/IbzzhVWt92nZmtK5HpdPB6BNGuYzOJ4E
h6RfUD0G1pCNRaqT4AkZJJqr3iXB1piEZ8DMM1bzn0kLVEGlBIh6TcVKadmKeQNm
Jb6WEpzN9APKfIYCHMNctTjnLroQDgvLgURikdMNBavYkMM5rauq5XKlziNFpzTO
5Iw42JRU0WB/bCdrkLy3bHFsVj+BbB/TOP0C0A1IvkI1KC1sepUC6Sv87reN8gUV
uIism3NO8wO0SrohAcNaZ+w3gx0UvRp1tUVAFqX3egzMUCqVvyMav9cOb0Ed6znQ
4H9QEM8NYccPaJJ6Ai3xMD18P/7f6Rv8l9b3oxxcFcpSUbOXfiULG+qSnPgs9KG+
YIyd/dsnqKZSunS5wEJK/T69S0Y26w7eY7YqH+LY9lgIwcD74QgpGAOlmuSvacBy
HQ4cugwErJKTNEFq9vaF0dDA/zcyY90FC6oneTyMY2B21mkHM6UQDwsbWLX94aLZ
xScTR/qTXHmKQ+w5sXwtljZRr4fVed08YIg3iKQ1SwiSoqTnzpAeCSMH0mUVwCSW
tYq309bNMwlQEl+N39axUO5mrcPMFA4yc0zxGyDJyxUNTPwJpZEB5aw7JYmQexUl
kcYnggLRoGx651Ie0HQdLbmQV8BrYAa2X1f++5koy6EgVpenKvCZZ1LnuzI9X9dq
1db74cpz5Mst/9goW6R38YGo3EtgvV2gO2yMizoNw1Pc06SARuOx9P0G6YBy8p05
sanRR6QH0mrchF2zRHU8JRTzv0txVsdT2PBDBb/S5qteUNq/f65tXOTpmKJdEWcO
0cm5gYeUTdnhXJoYDTP2fwuOydD24A5bL7L7Z3KZzXfs2klUSW/L1RBmIhvneleZ
8D9lqEiaH9nKAMYbgawyB4pNQKsJe+QUYdDzprTurNJrvtbWJO0tqRMy5WU+RVpL
otN4LkRCKdkC/JCjbJU0eibfM3sxca3hZkeA6onwSUNZHCwUmG/X301W49vAo0jo
fyYCUC9Gh/m9wb40F35+dVY2acwg7l0mRV6JoP2G2nGfoZl1xH9i0JCQXX3AcShn
8PJ3hhBlWnUoHTM8H6Ze1tmltRvjUjPAORVJa3pqTEOthD7ZzJ8BiJ9MSEJrAUNB
ZvCzkuVOPmLujnjKmlpt2PnBidPmShn+jAhYNFGbIXuYt2VCw0D3ZRiF2bOKpqCs
0k7AGThS4F6KFg844Q6ukzawYH6h+TkNcFY/hy8mVvY8b9grAQaA6crCi9siWJmh
ctaSF1KzBJoHIveaXvuj767p14+KMttqP3ftT2yfNbaYV46BBtkUzdIfFG675xzf
S5Is6cyPpMAuX0Iriuv2SL/cVZttU9Pto1VCj8U4+Y1lMFJtpabCz/waQ8kPi0LD
BngJgdIpkueYkGlWNyMvP3B/GhbWfU1yxsl4QZ1lvSutjuwc9NRIW1yBoYuO987p
RA0OGW/hQradHJnQz1oLxqk3SYDj49vkwp0+AEvWTdIZEJ97GkTMBjgnKl+atr6J
gcwHuce3/1XlJBLqzqBwh4cVAq80SljjpmuBxFmccc7o8jDt6Du5Wc5o75+061TU
Ox3FUoDoYE6Py+4g6FESl9d0U+XLv7I53dfz94gj3w3h3gl4/+RmEVrddjFb1ChJ
WDmnuwnx+bkVPs7s5kj4xBZcVst/6EHgE5VZh4Gb+0THTkEtLziOlPzerAapRAlp
qhCQrX7OlAbwDYnORKaRNC1DB0w65pwdYvp2vCm+b8ZwrIG4orN8KR/nr01siDjX
UEWozgsTMqS1KTHWJvGgcBO/ruWr4uxc7x0ToRHWhkYCObHXsoUoPM7T4e4g/dZ4
2woqjfrtCE93PrYiTuBlEcvRezgori6ZSxuyeDqUvIs+4Qr86zvwI5R6cRV9396t
cSvNbmhBnY7dnZ/JjAkOWMf2GLtAlhYpRRD2Q3HYKjYvMJ9r125zUkrYsghpILAc
X/OuqqAy5lPZZFibL6bg17l5QXrGSzfB03B8KZgIVN7Ly8+CajiGKPq+1FBhUZA/
uBJ/g6ntkHlfEFySBb5/A3LeRdoyUenF34AGmO6Judwf9gnjfmuJcbHrty9CEVha
hS0pezT9oyOYhJ4Nsi6Axqfpv+OVof+iX7Eo3Hn9rTZmzOQLMYO/C0Iehfv1wjYq
i2HitDf9h83doJ2qAssmW1ou+eas/7BpIrP1qHhUtr6LAThX2F7oY83ILmo4IPxP
1HKDvCLKVU9+JypOyuDp+uhCGsW5uuXEr62Jqrl1X57Cn4euCKbCq6spUXMAIlOw
RmY8FX9YcdTzJS9qlXPzR32eFEZVkD3qS834ErNRiRY83s1CzcCUpnpBIk0jhiN3
uiHEcbYfIMFAhBTcP+zELBDpXqtZQolDxBGf0pnp20xo1mklJ38SaBuHWC1GrqH7
OzxRyOAJZbR7IF+sajNDswv/McpBRvGFFZ1a+x5fLrvHowcm/Bi7HPxl9sQNegN0
tJIn3auuZgvUyOBjZQpjazoevs0jWDGzuEnQ24RpCITPOHFgG9Q50tlEe1PTNZK8
x9QXuyjG3FcKAlSBGgPrdiydox3dgX89TBSrSr/KD8yp6SMrK5cgcc+u5OexnLI+
iek6ZjE2RblvyYo4EYV/PXEJ2J62Otp/FNxmHGNnQor3xifl72uXl4zcgKvFypie
GOasHeI086RTNZd/rN/N40t+HGLoWazfAU7aeHdmZRrCIokqVm4AlOKWaaYCyTgu
SM3UnFNsSUw2Wo14D59nRx0cTYxZC1mAoA7XCSH7DgCZ0gU3/RdbRSkoa36QHhIY
idHDMLKrEAawG/rrrqGkCuYpzA+V7LGtMZjxdrk4/14WLwNtWr0m9E4QgudP6GPa
eBfTaTYYYWTsOovc4/uw612gWtY6vvrrhY39L9/kSWW18qcGjtzeco1mD6gyMlQc
zr0p7L9XNyOeyvF+RU3xE047/1QdV0xeFViG6axixd0b+xrIHBkyHhmJEiPxNKLS
GZgIwdtHlDpF3Cc6EFwGCVyZptoM9Ji2qOILc9/ucz/LbVp0wVe6m+0zlSS88G9s
eZeG2eMVZmlgnACVcZYermbP/JlkFGM8bDLBPF/ELclHF2nX05aej2cgfdJSmG57
TDhs6rV/PU0R69MvgCQ2oKYsDCNcUk4mxhRpSHmT4Q0iHmfRItKVdzwOY1Zwb/Y9
Bh1UNV3yIH6eqZhtqbSukhZ+ggExmIWSVK3inECfiwshMIH4QfUlypxK0kpCMK5Q
fuCf9t4eKwB6L9AGMD7yE7w8DJaEgyiv7ySsSN3B1GUHJ5+5/yrIm9KA9eBBtDko
k60aOsjix5K/b6EPkEfzdxlDIJ/NfTDyaRyWQWPk1i+6H70sxsj1CpVoz6ACEpbo
ANuUEUfAK4dSBQ8o8saFwOnl7zmGQIszVeRI9yectZ/GEEsHHl/y6pKt2/0LTrny
DkhUDUzThCo+hPuGXjBt32+VaGY7/j3ykeHHPB7T/bUybWCeOZVRYLSJYkdOpS6W
5n7I0MK963+Kn9Cz0Bg2cpJl2SNQWBKJw6a4RMTWixycWqKv+qPrJPoGq5VTs2Tk
NYQfO2MuDqsud57cVsoLINR0xYhORyUjs95o4ulu8WogQ9eGqd21I6iPUxemSAgZ
81FTdeqXqIy7xmhlg24GYIZ+eHeZdkOmFu5Blj3jaxe34BpeUL3Sh1QJ6UZNNaxg
J7NJETksxqdULmkxtok+urafsHs+OabsihFo9gck54UhmQCjQZAxicDC5JfIvfiy
qWLqxXUrOfxAjSewkkPbZC1r6JszcfrXkWu11pSCUGREJcyC+aBIqENQVoqsGlVA
tYUx2KQQ0DpL0tILZjBTOnSohGR5QJ1eUFbna5mlCBhbH7VPM+mchUohq+74mL3i
+Q2d83gxWYOcj/exdk7QpAdFXuRU+zIuZuo/c/J56lajdxtaaKGzQulxpZQJQY9x
vwpQso2u7f6RcJBmNUEPQRMfwKttOQMElMb7JRsfnylr3MaJLOrS8Sp5kY47WPCd
cUcFfUEeAlggcgL5DApudfJWiQvwC9dqQsy/qJUl3lD6GbDTDgYL5flXbUHnGbhe
0K5oK2gDL3QNDmLtw+MI62JohtW5T0CcUaSC45O5dDKZ5Cric+092MmIisOchLZO
IXcAjbqg7l+CE4WGOSnCQP0WT7SqyG12V26wJpPjjVl+dbczv+Ci8epXf8HyCk/z
jy6lvgtiD/9gz70PBb1bRoNucHmwbXsSIOrAytguj0r7DA9OEi5Qyncgfdr6epaJ
oh53nS+6cyeYD6i1spYoPVELwCCiVNonetaF4YsLYuncEA9GcjeprdRgfYBn8EPy
AEbzZRuk+GdMk2pRAti6WWOVqAWPwR769v07p/14mHfO4nM0w8gOcxeQbYjs2mIf
MAuiTY9vmcNkM0xSZZXzbFQno5l+zodwp5BVbRwj6CJTr0Q/v9LQRl/ZpZF3ev1W
yKs+MJdlzyMAG6Q/ZjC3RDo984GjtFbbbXII8xsk+FB744VR8oP0rTKuDqGMB1J1
/NDXrsV4UTjR9DfbQ/o/tCpzdU/iDqsKR/7MbdECwnQlp67GzlvWtyvvvXo9fQKm
kXX86mT89puCj0FqSHUe65ied4A2jr1RJbueoF3SUOaBHAg7F6ygfXPjmOOtJgmE
FOX8+rwnaocvsfgwVMMUqhq5CfRlrjKd4WrMdcg6uHZ+1P0E02de6puPFMtMiaba
6Vc5PWCN79ezCYZgMfF+S+XC2vmbyIhOXahAQUfIh655vdBAQjZs4iy1juBh/BHC
9oFgUmpDx3FhiBItLwCtOXFA005u25BY7N6zoIcsA9GUR5TpbeXe5XjMPjRzqymY
8FVxVipzXyFfjvGicCx8SqL/1mkP/OqLvGnXcZGWqrto3R366/7f0HXr1qltBVmk
CIkN3iH0Vz9XCqvbBYZF1HtXL2i+Zetwia4YwGeUJxc9RIPYQkxb0le9C1yU2ayS
/BTlqtBFHoiirfG0qiufVH0dR9K4+6ZBQZ22V3LCMSyCelrC/nyFKQpsvTQbBjv3
M9D8RKGfFVV6B2C3uTDUeWXjYdr62iKRy1Q1q96Xsj0jE3X8dlsVY2vg4Z7DvvPK
ED+wBlupOywj4CZZSKFNPFkPhfAcY+OYmNGTiT94gKwnk82HTG2HieHhJ+Ipubji
2Y4rhDBNuKrWgjyl5oQlwrZariWbgoF+haesX7VRm7Po53OSd1F8QsLi5YT5LcF8
garzYsNX4p47vZywu+jUwC/TWbLcIaejxNehET1kI2PYWyDyexMRdfe98ujxqy8x
bnefZMBkrKnuROz4RBLXRt3Rf8U41+QdMOj6yKntlBNcMB3zQSk2an2nt7bY9znq
rMMhsRqTal4FxwnG13TzZkv6rccojnAB6aKnUPUk8fRt8WdQ46dHsHZfbV0u4vBD
VxxmyZDGknYni0Jj5gIWAYjy6+DQiXsB1mLq3pTXKimwh3FDY9pAhnKo8ydT6H1t
xAS6ny2fdJUtRhBz1oVZ7Fkpp09wVbjigK5KK/bQbcrR0BTb87aaaErpuEASwHe1
+mAmPUaZsp2iSe4gIGeBlNe3Kz4IDrGSNh8KOtY4CLOuANFWbgDj9S6i7mXX9qEJ
ge4zfVkMbPsduVWTKv/+4WV8Lq8q290/c6BNLfCPY9ohht0qH3y0f3iUGeEadlO/
dJW4xbMuxoKFoVgCP4Z27wdDBURPxLtYXTjbpPC89VEJaYVjlIS/A5URfYGslExW
d73sUhP7faJxmy+RHZpc8ST9Rj5f11qNN9OWIOU4Ynv9Zf+wysBprFZwX7ARIIvm
pojNu1doCPQIx9j3s5laFm+mu04hOx6zbRK/W1tnDn8pP59s/DQiV/wxLBwxr5hY
nr5Kq133f1IbcdMh25E9X0iBB8EFPMXLGBntJAareMpfVHC8q0pZ2f9YY6g3Qha7
ijSs+28BNgbXSE5nojjr+VF5ala2N4Zy2xMdT5aNcT+N8y7iSH6FaY9Zon7Mq429
GHhyhB7yYY+yIfyzSUH9raQDKpc9jk48g879Boh0XQF5aQTN7Ecgz8zoBNAVkaOp
68G/VSpdvJTS4hT/DwCnlqNmTx1ZC8mv71J5vYE3twAsUly6fAGy/wqzJPdPl70g
GnmLJpRJWpfhQCFjvc2BAIXC21cBTvNPZg937tM7BECiwwTVr2dH5ghyGiFwMns+
ZpezKG608plAH3YVwT8f0mjFbb9atcheTF+QyZgI1zD06bRbZhORY/KRomR1RlTD
dPIigRvG5ZkncowHUZpnOUO7AIfzYFupXyzwmGDwtjZgYyAKbFd+k1vx9qdMEFdX
zLYnChHAYPnOSiZqOLeBbn4bGXJdIgSaObG8H4xEWgKMqtdneI3yhGK9ffDCsWVa
m0A7Dsy4Meb9tpzcoKhbQyecBKYFGpaOhncVmw7DqDqrJkmpheZoGCG9HTdSIfsU
iFL3nl4oBfBqfbJ2A2ZFLHwUlt6lNt5H4M6SLtvkYZjxkUazD/WYqPaTwnddruPM
/mDPX7lH201kdkm1OrL/E3otoCEex7LJDo2iE8bP652OjstSpPzhruu06ZA/Gwdf
Ncc+/Voec2IDSZYs/X0fRXp0UtzIEZ0PO1nVZSRAhOQ8HX/KoszdhLdw3EA4DPQ5
RHab6ExpXRMAt+Pd5JEHI3ZUWPf9K7j/K1SeWRH6SfiwyqwYlWekDak8MTCpIgee
/6+1Ast7LklVnv/Fn9lCihvT6tAeHEQT75XQ1wxg21eUNNUL0mzbaZAqE/Ozk908
UE/0uHDnmtPfeliSttLhvTF9RJn/uwI8W5NzZQxP/wpXdijQmnsNIcP5MhmaqtA+
C3WuPokm7uM9Q3xMPMkeJ/EZ38uPSmLEiTa6qapwtrwIRoTyMfnNGuORM7aoW/Dy
aLenfgQnojF3DeMbGrMzhM07PkC4xZK9FJu0i7zH54E46wiRJhSyt52J1dJuyKTt
c23QyCnWVRCtnJrNYKFJZf9Ex/0pw03oxX40m/1WSNwZn+RbNxpUpp6qUyLcoNMB
WCCikzXybvUICWwGDL+Hx6l34gHa8KTp7w+OeRutg6UiT1JFn1k+5cY3LQd1kGRb
eouBYqG9qBN43qe8vcTduxQycHntDfIeQF9rKrnrMz+fQk85W6D3+ekiYyZeinGw
qkSXw6IJZB859Al0Silax1CWDgxOV+g/a2L8oum8HfP1BTbtnue1H32YoSIU+RIW
bpoBjULmen5aFpk6qT+ls+I6rTH4ZVUGIlalAaKiFJrwJrP1ikrn6r4LlJrlMJYy
M7bqOCoekdQAB9Nt57bkgHP6djGC9PqHl2qCKFHftiyTbf5QEIoIEj6ufb8Ef+oU
Ipw4Ipbb6oXNhK0LSAfdbfeewJUnD0bziimfpEsN1pX9yxKFwDkTTl1zANaLxefo
MeGWo0sNtMEXhOjQO5uBEM7zW1qg0GisyZxEUjXhyqS1Tzog8YeSVdajAC/nMfCc
4MBtGdL9yiqHZBA5ou34T+c95HF60WueaA71D2EVD7y+QHx7ed+KaSGVPvhNenPS
pnmJsqKrapbZVRL+7HDJCMvTVjeoL/A+gI8cSwdWXGeOil6HzjFLM4ESl3x3YZdj
HAt/9H0xMyGA/hRuRP1rE8p8uNORjCwDNj4M027CESxIDQJbfRIR9B1GUAT+4Oie
eHabEOCWMdCn4bFRKeQh2uhCIRIhGF5p/7xsJSznJVIIuvmMwkagvApVlQDDC99h
TPxXDp5zonxKTc6q9sXSGTupMMryJN7PqCqJvw73vKKXA9aqjhtxgbOBKuiHOSQy
nliw752tsVvA/Nmdw1OpAhtyJwcVihaKD5M1oVjHxlwHvyB9060So+XaAzPrC7a1
yF9+/gtmT3VO9/LvAMC4nl38p7wnmnbKzSK1VjCBGBE6IczdBJAXN79wOc95u6iQ
Mkg0cvI663RipQA1oLgN7qO0E7mWYN9izligkLUzorZnfgqxNPGTN6z1T4M5Kv2U
IuwonT7u/vFq0RfxS92CasKiHhZcfHR9+JBneDiK33BV7upjX0aD2a+/PLL8jhWN
/PN+jH1Vs82rdA/ypIKKuJkAfxaXz6YX3Onj0Nv0y8vF66Hdnu4sqodaG5EP9Ml4
WuwBS3b+747Kq9HjGzE8sOAboiqPqMUV8KRXx2KbNNYpRzwvfqB6lDPbw8PpNP55
wKD+2P1QoSe8NJXtvmYxAUh+Njp0GLay6M4YVutCWDsjEGUz07b/z7MeWg24WYGC
Y9yQYF3kbjxQGsNKKqaBBcWaYGU7BP9+7h836iGfTAuJaZdyfRwudWXX25XiKWhN
H7+pu5cs6cRhPEZFNUuDEcHBu6jh7I1gO6sBedgUWPaY4BLlXjRXXpDSKlYiFheI
83NjTFL/Rz9iL0rVjhgKxYUk5ylHF6egQvxrN4V+7QocqYznAfE9SqpW6ilxaOFH
o8na9lxuU7uE25ua4NC3wBb/B1zzS3ViwSc6O8NPoh5en5x8BgPqn24ARS2Tb+oM
Ynml2MDvInPn/IerIl2XSk/hPx/ksb17p3XIIlG2jNB9fgzLOQr7fME0ek2ayKnR
vgPiuQ1XV6gl32NLapud2LGSSHXRMezdxTPC0u0H/JPAwf7sQEEIcG+cinQyZms2
QfCQAEuwG59NxtG8w1Sbca00p20Duje2HLRN6+Qq4jWt3sCezcDQnJIgggR7FFsU
/viU3ymvO0UJjEGmnt4v81ZD2l8R4fcRbeLfrFXVL9QInhEVhIsVp5sQ2CQNRP4t
QCpCWS8e27H+2dW6zujsgoVl93kIJXTs4GPT8SOdpf1dcFWNArVUJlgirij2Hpe2
hHeyUkInVX+F1oUsZL8scWxmV4ZIuMbsF8n/WGNT4PgFyswQRY3bXb/yxjKyxJd+
0A+SyernDB+ezW+t58CMRsSsd6/MbDzi2RMlpJo3xPD8zJbc+RFLm1Z7Zr/cESD1
UJBVu2Tq6EU6qcyTjQCR9GMaeWWiAE7W0NtmUgd1klNAXFiJfw6ML3DyF0Twvzz7
C8rcyUrLKrNu0gnXWFMP58hO1VTM0QrPkBMwbUS3DFkScCNTVhIMW1cgK6zRdaCa
bnbcffXKPNlNGM8Kq3UqBw8cMob17NOotibHUxzuQq0UBuX9OuxAKrkgw8nUZeYo
P9r0gIeE6KfH+4lQLIawXyNYy68BgDC7Aeunbn8rhSNzcM/3jEUXOH68QlGemwJr
JbOPnWppOBP3IZ0BvPun2M+YJLUcfFUBP3vWtr5IH6CLQUdD62kWeFsN7JOjdrEb
y+E+l0/7BFbh5DpKTgA176cZwZTzTRDJkIAOkERuWzzdQnuqta4APtQ2//gj1Pe8
nPV3gy5HgDVrxshttKaLTVoT2gIwlKSykfVExGGYkh103nhRy4xJd4ctJb3FhCQr
2lV2/yoFl4BSSk8XgL7+8v/yPC0tJAkbsRS8iPrrPc54YL/dzzsgsN07fy6cNUn0
v65qRfON5eCmD/G/V3Sg8FJdXdi7kVeAob9lIPzJefGgq+tckGKAZNuTEO8T5vnG
kACqSgifLYdZSR5AC388XzXd5F/ygvaXBHJ7Y0QELveUTQCGavx2o6vNcIn14Akj
uvm6i0oJxI+zLH5xFKGSkXyX3OMpn1JQhoShk2DZgcktMXvzfBXnYyowVQu4x3R5
+5GPebYVxqpSEc1aBlH1TjNqyej4XtupPpHikjT+BN6/UVy7+mN263xmpdbNxySN
hMeq0H9G0KAMQDw5GlnsVjONIBbQd9tk07bEDbzun8AqAPZLOLFatk8o/JV8g9b3
/0d/FhYeW1o2JzPsYHzeQq3z6+bEh8rjcWkwoRfH6XwT1JIKna0vnRPbMVYGqe2n
Hcl42yyLXbTp20BwMw1jZ/qdKk6dCFSTWB3sqHi3YwNEw6b9DkIDbTeuN2f0PcFw
sEX7YTnbw9KcOhePb66L35fPl9WDh9Jh1vOaDb0uW3TltjthgmuvKwYdE+zboB4n
elbq3eOug/yDmE0F1BA+XY3tDBb3dnsZrUbHXQtv4x5iqcZlevPSnIi55JTxZAdV
Nz8a2YW5zUOr0o7HC6T2j86uH4iFmJMpGZ1F8mfvmHZIq004+OGBQT045IjMq8p8
cWjVWT5xWy5TPctJX8BcH9wDpi7dPU+OJXiijTtCuXuIZurXesESDXHbYisPKJkY
wtAtkEAkRxE6/+yHka41RLTOMjMvVY4zbMz/CIGktVOGI7fFa/VzKLddKLQ48YqU
rivdSZ2nOTtcsTchBGsX9zqVN4Jzm9nw6XYpY128cjOvED5poLy07oeoyDGzfKlU
ZG5hCpUYrWTo8uaO5ysQO4ACmxtyBqyf3CecXFeFpW8lYDILhroiSbqT8wlbCdQw
qh0EP2VxgNKaQXloEttDdLL4FNDss5AFBKZecze53dQNz/Eibk5J5x+xkxJeXZwL
+YSGt5TDQKZqXJ1BjdDhuDuJCMTM4GB/lhoKm7V32Vg4+HwHQTkkVjVA6B4TlHLf
Uxw93ps2ATcGXSEx8Be7aZEOJ54/+Ri8D5d+BmNByW45SdAEksJpk5JnpMdeE74U
iW/2D/SznXMokBMTLg/NDqyeofFx/SkNqLZi5aEcIjA4JHYl6Hg434rB1AT2j3aj
jSTvVnOdYRnhgYGUnFXS5AyaqTpKUtvWzmA+bhm+fB0tlVg0xqfwZkyX2AOGrR1+
RVRR73mqEbCl7jRPHeZwl66qeeLSRwZquEvuxGITFRiqXIYET/lH1IR1zOdIGgbQ
N+5vJ0ORfewdtEAq/AXN4o+BIWf0WmRCNbmlx2xwQFE//Oq8xLrR/L7NqYnSg0R/
OVcVwY2Db2g8EeBRzcAc6gKKYDIr9EHe5QthyRlh1koCc6ev/+bI+RgbyIb804b1
q1d0ww/NJiY0b4HyDBD32uBm19DDYwEwHVyCTxa+fULNNJDcaE2DNLE6yQvXLyr0
jn3F+BqEVMIeZyBGpVCsTc25EnMK3tBbZ58dhIb5Jq2xXTtvODQ0i7D6YVuFW8Pk
I9B/XmWB6UYIVLGNxd4tXIVrhdain1edYJa4NQtDRBTCNL/I0d3MCYFE6DWw/jB3
zyx6te/viBhIpq4q79a4ffDggPh3rEW228fWQnlMOymbxaAPzyzHkz9QEyzEk6BZ
0M7ofvyM+cC1g+EBM25uwz3m2Yz+53TTOC8v5NdZBIkJjb7MDL7DgjXh/4dOCMnU
8hcMEwTox3v8JnqJdEfEoFx9cPkjDyfyI7/xzb3m2ryfq8Ms0eIZhLhkUsSnp0pn
I7dZAFI5vfPlmKUlbcdYLLu+0S++0hktgkvVnIpTNXGZY3NsyDDNsG/zJVal3nLb
SwoplTXwGGgkj1akLJIMLaosHReurLAGhMpraNGrvgfVJkiRqvVMV8ECzLhV4yjs
WM1K3AAqUmFx5FhA15ggqwF0gNm6KPXfsdK8qxPqN/GDETqS3hYNg1fvy8yMV/SH
WcWSd6XcpO4Sa1m9Tr2u3D3VySOgKCO43zP6WPMkX42CKLeGkwTSqs3w6EM2RHUj
1yEsBQ5Pk/+u3ED1mKvgxcabkoz26PsROibzb7lI6ObEGoLyYaxS0TSMmlNcsx62
4udLoQ6ArGY8HcSUUNPQ6LGlL0hH790QqWIMwy5NPRLxbe5c/owdJg9KYfjZ+DG8
+RL1AHnc6ATPd8uhuOBBHSYD/rssQuWb11E4w1NHE4o1akfUbIE9mw+1y4dW6i6n
CPtslU8jY1v1c8gP8vJ6dRLZp2mOaMI/eUZCZi3yPzMHeU8urSzf3Sa3tGqks3/f
qleiM6YwFPHJdZsPWTV7CO3gdp/ez2kdq95j2/c5Bll60ek+p9rVrPItGHScAiYc
gb12Ku+mCbUUxWw/juaSJFVIiTZV33Zl/gVIqK8Zo7ubXmupCafkiw8zPbXEuKrq
kQaZAAqdsn35lnGsiiZgPfzQ2CIYNJlclZeipziLw0EajYD7WxUXOyFG2uhljU5p
vKN2Oer+FXEK0DvsvqdrT0pbld/cyR0Ic4ckdrXKA8WHL+AINNm4RcQNpH9nZyfy
joNU6a5WzkyTs1FScCoL1HBItmrVxXB2EQ0GRIld5OxTtdKov84OWJCWE1c3M1iR
TxRWgD52Y4mCboxI2Els7EXPov5ZimZS7cZsqI0fVV63fhWSnm0tKvzK4sVGLtyR
TLov4DO+N4ioaquHqQzZHrnVmu+uLydsz0B/CzrPT8vN+CdeK26de+9tHGCdDzwa
u/3thq7N1dAX3fOXJC/dA5XPm4uCrCtP2TaNeXNzphv1PGez6UE5Tcjc8BYnozb3
f97SXjdkLIvd+F3E0dZoZBg2J8rOEIvsulO+4d4lN+3Rc5EDtIqeHSfALtA0qWMN
JDwoAY9ECO2qNskqhzhSNusKOqQ0MhtE9yBYf2N1H3taKpEPIHxbMtKPVa2xiHFP
paKpStcFfahe4248/yU/iurZju7e9itn6jG3d2DmsOcHSa4Nog//Z5njYRlavRI4
H4K1Pz0pvIZ++hsYx82kjoFk4dVQQEnVZQ7XY2jeO4L9icll95T6BYv5Q3hpVUuN
bTcFMkemlZnOplXOmkqhCr2gaY8d1roKDOeTgnbeg5mEjg6Fa8wwq6DfNctumWES
edZdfKpxTc/WRzk+8EpXucmlYwTBZ7mV6mQEbUF2tIUkQeimAco71u+XJt6wt5Hj
yKYUoIJfSn3XQ8+lT25QPQwMkksGJdz2smCBQQlPLoPdW/qP3wz8ZkbKlVPDmPLH
EPN/sFCb8pysy5MrJWl0o6vAEPvEMqPTqjIIdKOkohaaDn9gcCxb0HE+H3/kz2bR
FFNFpnOXXNtV9LlE4ZEKFsOBCgiT+qjovVYSFgGxbIgyyLqnqGh/84zb76pZNhUD
CpR+DFqP2TXScAcQezkFiOuuwOJK45vzbCdq7BjhVWWfjbujWVy/qxRUCsKPjFkL
5GwY6612FbLdUP9PDnIKnxzUFsqPfhM39imOi4gRFXiv8NoxazthXSCtXJR4jo+R
1OeHw+KgOTElMdbYNcaKUn8GNH+hO7+bOYgcbiBh1POWPyAXW6oHzCuYkbW2I8j9
wMoYmL2b1rvQvffxGKa0m+aLx2mrKh7Z/VXt4wYyTy1n+OaufsHYTY6rquza+hwu
JXrZ+XbL4IrQMexGW8fYKEe8VoRXcoLYE5AT7gYemROUHIORtmmQC0XCamrD0WNF
QLjLwXTNKz3FjXpxftrzv9vzd1zvNWChfnwApaJMtc6AT9xprLS3rfNzNf/khsTq
iCX9I7OYlQnVEqz04S3cZTQigCGbK+krWklYH1oyMtEZcfbFcrcQ53U2pVA4fXPC
qp3ekqcl+xD3B1xxN29rrpAmytOe+MhuDjltEjX6f/dV+iPyGy0KN8Qy99iJB5I5
nHWMRpJP2apqz9fiKCPNj4sBdabXN61xmvZdFyPDBzfaBr5ppt+0O/BPphIz+geJ
qrO5RFgfNKDAbRkjYYUGJhj55trS/xWWs6H8nqxxPO3SyoGR4Fu5qEGpa4uMBjvN
bwHECN3md1FDftwc3xs8gy6IFB6WH301C2d83itToFiyVgHjOgnKNOd0fgtrHBTz
fmmajl6xFhlxHsvmGbVWHdLgaOnELds7Ax9S5DZYBSJGQ7uwdWgVszLW51T/gEAo
gKuNE/4y6TYdzsa70rwFeMERnnROUs5RK+ViackYVLbPpQAYdJMyyWBoX0a4Fe/G
xN7bgDdZehgXpt6G7aorvefIqlmEw4HNcdkh8NfR3k6FEHBWdFq3K9nrxfA7KPAk
pIMK0awnEi41ydbdni2vBQySNS3ryGQsfTsMkaGV5Z6bP1tuDETHLLFgwZ59MoYm
T2EGfwbs1fqdfEGG0Fz2cLb+YkeXxM1NdNwlE5to8hvGhU88LP5OrfOF5VVEKpQW
Y3H3RNwDYgvqGyxJI1Gtr7PpAaIprpwHZRl0YD22o1m+NA/YPGdCzk3VAOQJYNCm
RMkXGQGIw3B7Y32sm04B8kEGb90I6ZATLejMVB7HN3kSjfQLG8esEKpAT0lnyHUv
qShcyxJeoBUHPvWcFo9wByh+340+boHOLgwnv4uF7nabysiGBbuq5oOLbwlxGLhe
RfwG8CHOXRgJrOquWJ1DoKURoEEm7db0XrHrObji98ZCQFDF2tkUeO8daVgmECJ/
r8laKVQdwmagS9N6KY1pqyx8OxVGKAO0RMk5PhQVdIVXOVwc2iuZEwjHKn2Sylsn
b3goXbfyKw2RDdym/0NX4W1+kvg/cRp4I5izybImzs5oy2rR00Ea9Jjy4DuS0Ol0
pOfDXwD4HR4T6Kk38k05daEXljnY1FQNsOr7iYOE1xWhzHEC/HTgL3JURTnQghFR
6Ruz1j4ehw8LGBwYlySn2DOUytU7WI8utVNuVmzhnhmpBcudThsVkSBXez5GVk9D
Bdx1I9GcEiG9eZOEeyPR0Rh3hA2ARzq/p+P7FfiScwWVidnnJevt03fCibFKsHhS
pCjw64GZCpukyrB/i1+PYrRLlt4OUUNIk6UZyDxqXoq+cY/YfStwo6434sIit1Ui
bkzJ85pTN8apoEj/D6mV04+zNbUrAQ6LtVCY+is8qfQPgQS5eBYjnLTw1Gvy3oom
QGAkQfGQdZUKpdGCE2qyDNdAdnWZJrKgZgrEkor2Z6SBKyIycoVf+ZZBfkLOwknp
hgHBcyw1rMYLU+Hojy7IWlazeqxd1aoXm2PK20oLg68l6EalpLcOHAtOPe8WCW11
v8IJp4g2Jlz/XRIHxKKmIohE8Jou/2bj1u7uTXx4HYJOrlnH1+Anc0PKjgFDHywK
mQyGlIbMconGcHJVdVDNv4bRsP6DMYGr9SbWX8uYtDFowR6TrClR4mgOwpUozLp1
WT2/FI6ot5Dq7lci+YABW0oX5eS1QbijN7XYrhEqT2MiutfD9cyZYpPQE0sraUVf
KB2bQww26xTUSXzt/9/CHv8E+KdV9pbzFaFghCFMeGQgUVL9Eb2Jhw6RcOhYg+fM
PRYqjoJyim4M1q571cHfWeKBF9KdSY1VxkXTveVTkGAnhQpAKfMy8mpfN2qIHdRs
GsZj/t+em8eRTzcpo7srSyxdqMKj1wkcFZB/JY2am+0bPWJUoCLpjWSCPHyBsw31
Zf7fN7a+KE7WsuLjop9GN3vHSAJAn6qHLPn6StIQ02D7B6M5Kau6rNMQhTf64W+G
8fit/cYQLFWp1Ej+vSZghqfKpsdAv/r5vk6HRJxYbPId9PpvJAa0t+r5/TVsxE1p
1xHlKFanP/Q5bW9qWMSsXQu3dL/Fiw52OcGCToG1S/73o4Pq35xWuN5h8h31JIsG
B0efkgYDLqjwM6feXtVgAV30RChIcaQQsfYAG6asvBqBec8IWn6IVB1S0zpRyg5x
OI+oJajG2+Rsn/o99G6jEJ3pz1jmiXglfnoZ0dTDp7xBMHQWbevwet5ijgH8GGfG
Pt/dSviv/J9TiHgwdSXXXr0GaOQhv3B3QFExmwugSJbmcU+nEAk2fl8ZYBm1Rp/K
1qK39uRylS3RG1ifrx2DO9HeovBXExWzLxhjMUHPp4xbZpSLGwhCvGPsfmqAJ03A
qDvkSBZ+OZdPCAHm2qAyRzcVZl5+dF6KT07KaM48UxBWczlA3Vy2rgwKr3WHCx86
RVM/n4rSqrn0DN7gQchEA/nVHPHqbkSJ2HaDE525CHjFfVD5o8aIEyphThFbTxFN
NdoqyJKeQruTbJRJQwAxdMIxlZXYpOAGcjSAuGgeQD7fFBhpSXOxa//RyFjiFm5c
TskMFV+P8OulL598Ycv9ZyM6NI0FhZr9qS6LMpC2M77gyu5FkiDXEw1mpDvXqz0Z
0QVI2s/iX0btxCzcp/KtOA0t28UB6/mIP6izwhJ4WrdPLShZeg0Ga68MvwnXCG3H
Q3bxY2anIJ4OM90zbP4v1DIFuNEySICvETvwEb63wILvaRwEYRztckV8Qrnye5b/
QTj0I5QBsi/ljg9Bupv3r2+VJRV1v+UZBVzdTX1cdS21YajwjQyBG6eWBLziCaHX
2/kDXxZJFOz5zWWWavv7Yq3JJ7bVVHCBJ+f+Pi0WsMTwpxZ+sv7fg/8z37mOdS6k
MeTePvY95xKQgSmlWf2G8AuPRU7LgHw4qJ+NCirH+kVp92lS6qRqarifGzXmV654
LY82uAL1KPcVL6jQs3cM8zIUpNC5ZBczD7xygHXVLFK1i+oAWvHqYUdihyu9Je6u
0O3YqdOIKBN5Oq05MAJCznjfrLNf4vraqqQgJA1Nr4B9eRIIJh27uYqQu/uZ2jF8
GWvuP4Ok37Ymz6PaGXjPDWTvxCItSf6KDdlmZXiay1XjiIMOf4eV773PZPSDenVj
sEJoV42kM+iQ3F+h5TC2i/HgSYw6B1amks8Lsi0ofos9IwIwW3e9FNJuvD3AZzGl
SWYUmX4+EEyjjRhZa06i/Q0jkQpM+HPOIF/eB/D34GfioxH903H0UxD6KUiAj8aj
a6BrQwng6P38hKfBLgOap05UJ5hkYkWVo4Sd37gC9bx+gdn3YpVth9jkFfTQe/gt
jSMy/X91BEmLaeyD/HNk2/CV7lpsQF+yZbjzvWkZXLgN8LLIHiQvnWdZhqZe7MzK
ONAfkt5kPD3fnVtsv5/iYXpaJtdhr1iURhpGLBm6Nt3OD3EmSCtw6QD1qdZKlRe6
HTshBBrFsmEpq17hNcCSjDDnzZ30D2BuRUN79rEAo0noOJjDElgf73PBDqeYQjhF
rveLoDtfxuP4zqU89s6/PI6r3UTrNtpErIDwz/BmKBDEUNqhQO0Wktpau8qZX3+E
LGzu5a+d47gDh0DMS88YUz+HYf1YPe5QoFGki8y7hZ4G0+asaAU/r5yn6axQnNoN
+Xg0lT/aRnhFcKuMqe/CzpkHhkNdpXjxkrgxDImRKlUmawQoqV0TsVFZapz9S5bk
Mk2R2GTesSqGvXGRc+6vKOwuRZTraNjuGsKh0wNajRolHWCtbRx7V7TUKohsexEc
aUGUSHHE6s2kV3yEM7BARPtvnt/8HkUSV5K3yQ+U/+9etQXYG43b2nT9lpoVj+HL
7Bsd9nXEhtaaI/dQzbBT4qr3zshrNFofnes2lhLdy+LU02V2IYsce0/+JCqItSBK
JaHJSSIsdMIeYtsyfpZ9fwRPwiZoTVQT/UKCwO/ut4tsrRcFQEFBPdluEnBeDGn9
HhyJKutyLL70p0wXvmKnaZXUgMhNLSrKrme18pYwuZ1QwAb1+soVMPb0yQ5It3fZ
iS12bOtMWx/TEix4nUN2o0rOFLQonqoVOmfX/C9ScGfkcYgWuBO4JBSGKiuOW8vM
x4keNMHDnp1EgA/6NFuHGRxxMpI9r//b8u+WJyntDNhzZOodcVCZGNnNh9Z6pz/p
Sgr1mx1uJsIwDL2qdFYvrWQ3sAQ2r97+9jfxF7M1TiC7QA890V6LcdOH4vo+I4Eq
hRW4BFHGAA/uQP4TOZZ9cGmfgF+tO1JdL3ae8AOZjDY/qx0PuMCs+Jvi2H7Wptgj
eAxwEqvdXqlK5YC/8Q76rQKUJ0ZROw17zSY7kyszerj8Yy1kQ0Ej+3o07kAt1jWj
/8VdaSglnReY/+BgXJMboaGL7QKW0hg1ShRTR3h6ywhzaEmgY3y6lhJgY+P482O8
OngF1kr9c7Gy2UXvtlAm96JNuM6kx0N79fTNbu133ZlbU3Ga73vf4MnFWxuNQ3eR
SiRVK5cHlEFy6Alc8hEUI5x3VXM5jjvI5/HXGSFUkH7HYVPiVy4x79Ed7rikUYW5
V5A3pYzSTkZD03v1k+C70O8fm/O4GLsgqDXFMAeYAj4u2vzNZ3Rh2EbKWxKle4t/
XShpe78caR44xvVLrjoqB0OZxI/wnGrdXnSxU0GzmxCfFBgmCt4YnXHPKCsjj00J
W4SbVl5DebTi9dYWdN8SnWaMle4cpekFDtXrlSFF0RloEsh93MyCNCBzwvCNW4/p
MEhkT3AkSj8Vj7IYtsA3rNvSAxjNhTzyGiFqb533m7TBp0cAWYym0qfApSrrfVup
vHJmV3fgyEzYGJKwrpHqGrvz/1bAtUIFNNkc09KremwFOQn2x7JEW8ZbwURm4yZA
LFEL7lIST9Y8C2BmoAiVOxAuvWOJQ1skA8I0dFkKMgq4BlW9uZMprpC1EwHNWOj5
YsUXSRIRZcpXUg4yoRVVsBZj4H1tTPfR7BgPVG9h+7/McLDYsxK2MoOT0GEctL9T
6SaQmmEDjK/QBSpm8vgcoNStnm396STvJuipdf8gN/hWIps0OE61Ow1xXWV6RTCk
3bchnKv+bw+CZhfsKiNAtlyTeSrO3xLj+5pMMTzlGTTSVrFWIIupdgYchdtudYph
A2BY6X2oMZdQPCHAtrWV1QPDzsoZffHz4adjDGRSYU7xw5QRtBSjpDMQ9uvei4MA
N5LAhhtXEW7HdwE6rlOdZ2mYSYSpaOHXKz94xAHWOIbEapKCMGOnuSCiQL0ddbXc
7e5+LiZcW/HAUn7EPQInq2WXurIE+wbydYoX9QreSo2lw1nqMgYZhB1/LPi6LfwK
FhWXDIrL4ZEmFusI+lK3ETlSFPnRiy3jRxC185WTkZRdbAQL400wtQGD/fyrXdMz
lWXIwIHKxCanRZq5mLwD3LRSqH8E6dXdanGIM+ETbbYrZP3Xm/XcKrKP4ihSbyPt
ObqUXho1OKQViZ3u3fSWlgLRN3x2SC1teN7MbyC8ybpQqgrZSVoiMMDr34rdlQY1
zKu/FzXKQJIn3BGGMAGhtWPJVEN0vC8HdQiV2ccfbIO1/3Rni/Ri4Wb+J3Gyp4j5
P0LcJDcJCmB8hYZ3lAnm8PVtaD88o0SgGwhoAjoJRbFIiozk5+pZ6ESSzTK8jsnF
HlUz2Wy3FE+yCuLr6cLka91DaBOnvU1ndJcQvwV839PZx4VQjMMpNbVpt9SpJewb
adKf5qUClMqKi5xHKcni+aU8HgkOAdoNWPKhYdCigGJ5zSyPnHf45m24q1dSjwLj
RMclzImB8BK0lW/eXaK8vnimDgheJ8qQSp4W/BYkLwfpLM9Pmg13R8HjSl6Nms3B
rUuQaeFAaUUIiOc15RxFpVxlUSR0MHpHzaJkxGTqymMFMQfuhHDcOYoXehebQpbj
aMeA5zaLZuIVSPal6f7BrqjnAYX9DTL8ndrgM9krZHwQ7njtPx/hh6G5fH8yXthP
6w1O4t3ehQQqYgmlN+Hbr4o2RPY0TE+1UdMqQ8LV3T0MGvb72STtOE81CDwjrgKR
zvuaMbsTbRQ4odFxbGscPDMcajOlYtrTbrR+rVWSp9pVE3R+3mnMELkdryBgmwlL
k9mNgrCaMxmVLVa+S/XcnbdcE6+4O6ftf/QwRy9FA54En3pFUv/vrEutq8nuF6kD
VWrcB7iCKubDrHSHV78UZ/vPHvZCFvS9i7fWgDJqIH5kj5WYSuNuUHlW0ddt98CA
r184faYKHEZvgoJBdvMQ2Ri7P+0gif8XYhNJTmIz+aH6lL/I7KWVoGmzvqw8ygTg
z0v7iMJl9Yc7TaUwTTbEZjor+Z66R6ILthYqFdmRps5m92KnnMm0r9P8ZhbdCxSI
ZIEdrIRivfqG13KdRqn6jOrn78ElpPCsNLkiJAB9EsUonYjO+RL70sT2DwdZgCES
OqepgYGDrCwgQ924YnpJMZRSoOsQN2vrLkkjWbSB6Tn8MhCakpSUkbAZ1ESm2LU7
ll1Xe5bJ+XipOltkSMpa9jOrI+fdy5++ldI8/P3HztJeLGoRAoeziaZ/UFpCz+hV
Nrl2SQX92qxBDyVSX7JDwe6JGmUTLErkOmDutlRNfTwl/UDs/bfwj0A7vpv283OS
U9dUWYI1A0zpdTirvRVWq6pLKAYS8I/GDGK7HOj4U9/Vb2P/3Z0Oau0/69R3XRoR
cX/9WvYr4cTmTLI89CZd7TK9xOdavWSU5DVEJmArmwgmQTb3L/41CpfKkdusTQ3d
jKKVauuDOULMwwsgSXU/cm35ZT1KiWFHZKOpCYR8jQTthRBKuVaUvB7b3a2x5vZh
MNwi5qfRe98Cuix9ako7ZO+ZJTNmA1r2j8oLKzBUpuuR2Mx85M2o6h4kqSo9vRxZ
8b5yyE8Cid8n9hlsFfm4tjinF2ldeubbvgTNd/DdPmM2s8PuLfiQOaBwxh3ksMyE
qkVoFRiaGnyH37Cx5dc+HQnvC3SvkhBsr+VCROTkIoMddsh8ozxwFfYYZlab9pU9
n6L2BAkJdKmpKaeY/yIJLnJwGf7Glqv+V42nJPySxXlTHrdV7/fChiXY+xgWpvzb
beyLJsLJdWrq5uap8hvsaP9uPelpGn2bc4vuHq5bErLhy68RBeXLYYmtTii33/Mf
ncB+SeYBzu0RJuqqnKhoXCRnLeeH+Ax6WmbUYyJlD1//hqLZ4kMzMis0D7UY/8T2
cpHVQaGRLmydxxzF/l0l9XQbzda/4OwVNtPfZqV75pVm/n9BQR//ZM15UCEUvnhU
ppWHeicgIZahnJ1k2Hp1/t05HkvbhqpiKgvcPpEDDqosNda+RHqRpdTKNybz6V7t
2mFMxAOr5sJ/5CUKDTM8lYPJyH85O5yy9Xf8ggIZxXfzoRzJEg6O55Hkl2dNFpRF
syt3uPjQ54ywd8CCv5hlglydQfqdETiuyh1L02LFwFHNz829VqOR4THI/5g9IsWK
GrIXqH5wjCiQzW2EiXPaZOPj1R/3P8LZWeDsIVBMiTYkjekhiBO4lZ8HyFuAJWYe
qDJz3T8ViAB7qDQigjrYNTrK1ZWA/fTddoMRJjtLv1zXr6Z5UrnL8R/l1GL2m/0S
8vu7jDQudKqID7fI8MB4GIGCDMWkN2xM93+1sGX7UxJulw/sikEL6v+lldrwO7VA
6IN4bLdIPxFXqaUKfdsz0Xim3HwkbF7isQf4f6kpVlrAgyRsStFz3drVYyXXvEgX
6VcxNJgHywNThadhD/ARw1lZnodeC4iiNuLpav8r5IY0l32Nkj7LMAZcVIQZuMxB
inWNpCp7EAqR0pShNu39JPFQGCBzZPTO1dE2pL+ke41m8HaGMP2hOAFG2hN80wop
bCJj/7xtamw+B/9GgHWFcXOiMOJgHTj51fteXfEnR/tHryvyERtMvMhO57syD5qi
kekm4NDtHiJCiliURmyX6H8VvsiQJBBL9BaQBMFFXz1YfFcKXhkhfEoaRgeUXnLP
fan5vOjQGQGzkVumBqd9In6V3UwsvuNHHU24783A6Bd4QjqEBAls2chLIyvY9Nrk
FflXqRsY9PQ9sisDr80I7bnTo6oxfOwemsQ1GeaTrsTPDtFI0N91khlVUs2gCfm0
pwDR5U4u552wy6ZD9oSoWNv2GbpOXzh68PR3Xqn6H/sq3PZO3sql4ZWR5OGVzzFh
QY6KDhsmUiv3A3D7aYtehdEJYku0U6SQrFbv6NRQMpa1a5UpHpXDOaGdRT/YyjJq
NpXg4UuU4yLcbAG837tudSjFQx1OACW/s2Ns2VpxNtBFvLGVtbX34kxd/S/GFJuw
wWtjrOKq6E9qRMzo0qE7WrzNE7173UuI6eRtffJNJi2TDGV/Xhhz/+X30hvQ3tf7
TwuDdoRVhEMX2z6CF04iBmGjsC+9ar6/x+bkANnd47eZ7V4Iab8ht6Gafn0cl1pX
lzgyVQbMTFGGtCtwEGUIYYHE6b9yyDaHOpKLmOjKdVWLU6v8RkrxbKznBijmRk7w
E+cpMGVliPd6nxdu6+/KUUTvCsyvSSO6iE/7JW86d4WUxMI+G8vCgT692qgheSZ1
4q1LVP5WQoHBZCavQfg+cP+79RAUBl7XgtHRFLxOzjQ3r4ApVWbn31wErHiJRg4y
5tjl7jb7iAFHeLMP4LLLvXb4beZgfFF/CFXHTKrJ73Li6WxA7XrC2q/4j3U/PUCO
jd/nfvTrQpch7qDQbX/O0EHaz0rAgGnL30DyXs8deP+gqIxooP+/166q3Pq7WsZA
VvoopGvXMmO2wpcZzgV6m6i8KOFWHRY9G8l559h+Xnez+3dxn77iOI15DtfgJDMl
KVdJOYyHMuXxBuiT72D4BgQ7aseY6iAwTFI+lbnLwUlr37EjDfEGwaYFr3MPmrYv
RUs3p5m+4AGSpLMlMhPY/dyk91jfvy+Evb21UQBmN25nGjEiOw/f8ZB79G3zDwTt
5TiSmGVNQZ2TuP/Jmpt3sNi8few9kWF/NcDy3J3K7F+YyKSSleapLY12Br+ouD0T
rJw/dhz76hObUD9Tv0TT3rjKM01auKDGBiZDxioPlCnJxvWY2SWIsBey1FezBojZ
Tm2Ko6/0RXzeIRsOkYkPGr3mgtMrzcs95ssjiZVf8MFW3gEzyp4ocJa8Ndxreh7A
QA56wmz8GBA37YBdJOzXxG9BW6aCVPkTIUlISbdRQiTufdpRPKMOmaNK27Y4CxnQ
O0+MfZP9QRnVrMKYeD4mnC2sV+MEKtDNRmaj/wCNFAt2Dv1I0CPMm0AS/4nw6u43
NLWGHm2mhnWPeIOlBhS6LOddczg534+jNPiHN8lVCSqdcViFeDxKactEx49gVTZ5
zN1VvE6dpJ4f4I6pQqHeNMVv35XYsfknaNXuS8PM2C7IiQLp0MHbta0C+7+/H4Lb
rk2JA1vplUCN4RqHyDOI00fMUyVpVn/uKj0QJgnVf+Gk3f3FKtMXeCED8tDltRn+
C0HCCPx8Bd1fMfmRvM7nvvcck955ljnWHD1vvf3FeAlYUQNg/Bz1RBbpYvQgEZU9
6zIzUdKsabDSpKEyzLk+dY5ubROlF98OhMjjgqs/zFrl/GxCh4meS8jznLSEa5zd
DMM1UKrGP1QK8zkMYL6l0qISQgHoEhWtLcfnCHy0xFvRA9Dtzvkyht1bgHIV81VQ
KGSxgQCPCBzC1Eb+adNmPNUyeAtbDV/EXT+SZPtwcgD2wI9kx0idSg3GRgcdtNvq
Q+5zTDel01pVlY4WoJBQWIWSUQUOuhu5VLrf145o3QDixgSKSZPA1PP8nRtGvKlS
aMMCRZL/NajIbUkj12jMAPzGjehoq+/26rQtI1DkxDrOmBdoOTcpB7hBB4zGjcRp
fIP3FQ3xVjuQts/Vu8PpY0Tkq9OtILObUHZbtv65bqIkj2XhnHgqCb6KN0/peD7e
j5GPjwLN5Yxv/+DRzssk3Q63mH/d16T498fFgNnXcysP11bgm1BLu1giErtoJH5o
U+aObbVhVrUJYPcjlDY3xeHnEhhnM9NGr6qYOmhAjSNFkm8cn9kYxpda1pBaotoy
WrtA4+vJInKXFgw2EcHz5QP/T5n+KCDpmKhtZU5jKB3nmtUgFS2WVR9YCKbwnAGj
I6Z6K/AIU3cSa1MN/SMD+J1kTZyo+fa6WonDTUsa3sgnjYrwb5AJQObcFXYC2X72
Vf8p5amguwbho1dWfjbbc52YfDB30h69Y/UBYs5dwxNeJNGDqZ9bsGpopmNwBMLP
RRVAj82Kafl0zDmBgNF3WSTLy+xA6yq0BQ/eCYA3siHZGXxdG5aX8iW6dQGpXEqq
zxAh/wtEtwXp/ZANhtapYOX/fP+ZG6nmc0osM+Lr76l2NFCx9PHSJcvjm4Y8RISV
RrTxAm5jwyS9aAtYJah7lblsS82HohCnn0cmdsHgTsJaeiGmaTMH67gVwqc2cgWF
WdqQKGlxu3OeKJr6vcMZllXz02HVkaQ9GzsdQtILpwxW3+SaFXFxZ4DKHPMOnvKT
QzLQ+FTuYfQbv1jjkdHNKc4OYkwh3fRHXN2w1obXX572tIJELwj9XsMmPC1HktGc
odpL2ljSE71aYkWYesVXtYcRk0KQFPBaPp8gkZABN+2dsgZZBQy7sOaN5yfiEmoX
UKe2blD3gTu1TlzRYj8J9q3pqEEJss9vagU78VheSDF+dnQLak3wzUald+ZZU2rO
ZAfNZvGRIEA0Uk9T5zT1pBFmtLotgOx4h10ERPvsh4Y/RXiB7yXl9Pu7x7CNV35d
0g05PHRM8y5fhoCfW0ilD7duoOYZJxj+F8PZoyENGXWkt1WU9Mc7u5O66QKJoG4r
hbGWVLJzTMxNRd3y8IpxOtLq0tR8zv7p0hja7Ng/hOFS03NVDVeN5tPGWvZEAs00
UNBezRDbglqizHKYpCrQJNDxFc8s/l8Du6s5/OSi2MFjY26zOvVQ4or4y2jdMekH
bvCfie9hPeQxEzPtTDX1N8yPEPWWB3aaxwQ9rCeEgoj5myzMV53o3IahLT0xFpYO
UPjLoBn6UfjHWgIblBEkVhNtUf9m0T+pz8N6KCoWPW5LOkJHaF/c62Us4KGPYF6t
kWsVb1mGi0poj1ONQLaF4vy1QcU47JYVvYOOKcWdOS8Ummynmy7ELRGDjh0VhoBa
kzDx/6y0XvkPzmu5Y3VBER00In0hWEcJ4A60pM5GeYPLqAp5eNTIZBnrGebtDeUh
Lz0tvhrkwz/zscgldRGnbsw1MNnci0BpxqdcRaIsAAjZqzRfPpISItC6+6fNyfxf
WKTuiE513XgKOnX0aEghELmV51Iw7IXuJcPxETvd5sr7+0O6EGW13MeIVHuOb9/o
ofd787vS0hQUNIDEEI3Xu+tROXYGdZ1Vq138B7lgpLczZ9o6kHdJSybdcnaUlsfo
xHUVSSECTGjI689ZyJryz8vBcla4euEbeSjUPrSbV85J2m/f2iZMm9U5uNXiuH8i
QesZvQekMM2kJ65QpC1NYNbyVnr5QC5KoGR/PiAm9a77v7yLUUwHYQR9zFzy8pdZ
349c2PpUIayLmogo9JZGeP3Ox5g3lbdvrkqJZsw3RYoFUrJgFXwxh1BMHm3PSWcS
hFGnbOAUjdF540VQSIsjMSbAcV8H9HiOoPTvU1IB/P0MdLAMiTSa8WQIxK9bPZJP
UQOTZyqTR6O12smot9GToslapwrB/GG4EjvRokJkc1QToW6PxnJ2LQhixqIDwDsB
dzS7p/b3ROAaOQAF41kxXghfjBCFshLwoKFPKuhjZVAZ+jPMVss9mQc/oh/eQ+Ht
9VXpDyPmkexzE11r5OfSXvgIKCmhhz0dgA+iPheiRP9oY74OjCzri/ioAAprApwG
FfxegFvNfk+Xx6fNTGorxeAzMh5W656IA6bgBJ4w8jk8JfxtsaO2pewRKN6V1/MJ
LkREmVk+cNv05ESKVw+xLd/invsmuApBNiWut7YYBZeUVBrwlb5sAOoIaCpYA4HU
vH393tNqUNNhI2tsXuk6pJek+hXbK7WOd3GdEiZ6x2oeqxdiMMTpvypgbCHcIYNs
aZsOoGFdTrsULW6WS7YpXMRebO9lt8jFDDGKTgtfPGvkL3l7c8ylKkKc/wW2w1Ae
NfZfQA/YRAZFPm6T1qnHBgawZHKoBvyfYUtq9TwfjhZfZkOz0/OJgWpVxMYB+aH2
2A/JHrutrIFT+uFT2wQJvGrRDOTu58YuIdAWlEsN+Mai0i2xiY0soaL2MAjUaBEX
8NWkdsglD1IuUDrw9TUIItfQCUupSbXK63KmMAUSBHlquD4mHjaw6TtQF81VI0yd
jU+QlNqxsbiTs6GKKBo0sJcwfb3ORqzANIg45sN0APU102VFt2UIubBRIC6RRHBk
PXCdk3hBLrBYI+gA6uvTA3qXx/rPRQNYTV93kpSyyIjboINJjewftrsExsRiaa4w
nIl0IzrOGcryZXlOnY6S9s0K6bSJHM+4niLxRxWycP1hTXdXL6RmX1afD4TvEP5q
8iglDcNzSueEApmuHbi9hiGmkG+eWovsRCQhusQSc7WImrHDs7xQegc+9AQeTX4u
G7hkHh4iO/nFt5fLAXGtBsOFr9NsFLY8eyanTwn2OxqDyt3jALQqVwcpW5AQw26a
A49yvEG2nzXyQ51agZF2pSThORvKOVz1VO78mkLWz0Ka2eDbYKRmffRq2l40/gWI
xvsW+XYONa0oES983xqhmDpwuJI5gwhmdKlACMjvZSvoNNUatlmX4U9q45laLSvD
4dfkZtCCeD5IAh9R8FXWneJWdlb8uFNjNU69nyqqgeWh42g5Ip+6I757I2zlcdoY
umtTBBtEPDGf1jeDB8lGxNeqIYcQvJx6dgQXrMmSumY4GOWiNCHwnCMqsGDYi3/x
ElVQJ7bqUds9B1ibVoA67wiMRabdtKFFRg1X1ZNn1Z3S90vHxST3TVG1rPx49oGJ
zGSnyKXi6LQgp8+jPxD/GzNzYORy7w2fVDGCx7PNFlAeJAP8ZmCXK0nM3JI32lFX
mlcAlp+H5OKEs1ToRN9gsVFhm3fvtTP2D52jOhUlMMh0ijFMKczP5V+Z1xovm80A
qzicxVaiNaMfpQCa0+EuK7e4B8QWEOm4eQ8+FRa/ftgru+if+bytvr9Nk7hHu8Gn
DzIGtr/RqeKCOmS7LJiRamXYoQJr9e+KIphmZ+1Zj4A6Jr/oiwyNPcNgSaZVKPeg
15F8A/4zrjj6AbhR6iK6M1PufvRkaJGSjwiUSB3OS3nN5fJ1srXBUG4qlRdY2CWw
ABTNQ5l8s/wd0zMoBb41YY8WYwZ+U4hj3Hj8cpAz74NkQo0QqSZP8LoKy/6rUObh
S2g/YylIYPnqnqVtyrIPQbebEYrevdKp9vSZ0Vlsk4lpjRmfCx24vqOvDLS5Wk2r
0f948AI8ltxn4ZmiI/OeoMB/54VEjZne7Gm1BFyHbLFw9hKohBuBZTNx7+WDH0WX
GNSwKNHzyCzLK+j3O+S5K+KspSOKGRVWAfxJjL/6orgNkL7K/LlpAgu/YPhTfHVm
A61lAvVu8Lvr+IXekYSlaPu5UUEMNdMaHhnrBKGdYW1cmiCN+8CdgwCrCcO/hxO2
c2P649xPojtI+Ed3EbBABnYurIXRkUPbmdAwjVG3KPTjTXbKiUJXzC0ZVJTuNE03
obbA8twSwB4TKB6Om8lp1tw9wUnYXxND7CDaKhFRH+lljxya38BvKKgrSzOoxcsp
UOKDJN1Fz8KPe/UDdIvau6DTvg+S31E1dFapFLL9JMXiuA/xNqXbaVVXvsiRUfpR
1kpPLUZKtty6fmQ0XQ55uRQuPpt+scWBvbF+y/ntVjcuJhCYHZyxStnyXjiNf76l
V7beX1Ct742n6+NoAyKzA0CWf2aDeXYShVrsx4GLY1YSrFN7YhbAxmE8CHnP4dwh
cJk+YzRTd7P/xA1eUTqLC8NtqVMlyOhvOPfVVpTe0AzGfChYyk62Ro7NSorB/iax
FQ8XXL7JP/GyF9TzVIgYwA8cp5N7XgM5e5naNRx/GVt5CEwCU553ptDjJyrn0gnU
DjivMUkkmvTdkalHHzbHPjztc5cAK/VcUVBs8V0fAcchq37A+gDBPOWrA7jP+nZD
+EhfzoohgP93Yf9AYTZ/pJs1tW+zfUn+eBvGUju6hUy9zpU76x7wb8BYPKS8ODRA
x/ZpZyPnaxvfFsfaQdYTMlZNXsLTruwY530accp5prhrtLeSGsXvSbDgoR5U2LTJ
f6UvAi3d3Lyb3/b6ug5iCq42kkg0IAGyzRZhlmS0xbhCmMIBf1Xs7sJzILfSlc9d
K5EEmnbp41qfPoZj4ascLkXJIMSKXrIuLuucWHYNFcYbolbnWIEVzhkBQPnsfBVR
4ag0kam3A7OT+nfrNVAKWmAGVdWDd1M0BNSIDkhdIgWlpN9SlXok2VMJHArddpS1
GApF/g02ObKwtRC+y7u/vyzgk2r0xUUO/aC6VRSyACcFm9tn4c7b0laTj4Qvsfvo
+F3JoJ8l9HywKLO7NpPxxaNexqUmhYagEUFzu+sTZTbR0k7Br6dhZPv9TmTsO10A
qHYa+p+r5IY9vfkXwHfaKcQhZR96zZoFTLnWBN/SC7UP/BquibEMMDt7fBzbk71X
U8GsrSsDjtGRawVu/8PgpZLF9CB/2c0dMcWtCWpWE8Ru86ANRH7jmbg0P53RenFa
vWiHWGWcJ4BSTRqn8v3JZc1pg3kOceJLQiNRewbPNP0ZP4UWRk/PRhQtB8Sy8B9B
zj+LRcHCtrlalNelObBfJdTbVRSyH8qt475v4BUDjQKxFzTFyQEfriPhVKn2u8hb
CRXnO8bGsC+ZDKqWx3uHlIQWdSwRk8PLvBU70+r424ekhQlK7uHHWzCB0riZQ2UQ
LPz+54u5hKpz3tLojt0/4/niQOuPVbsxtEDCz+HZfl7CqPrtz5GfgJKHwah93sWH
Tswy6mu4EWQOSP0S7a/tn63PfBUhGZxd6y4u7V4L9sCHf0Db99f60Rvb3a2G+kG8
ZFk9FvH6s3H6Sh7aYLEC/pEK/zuAhi5PCQKO2/+qqXyOYAulP59KKKXC2VrTYcAZ
Zet0GvZg5Aw2tp5YNsYyT08olQOwMpTAA430divpris7U0iB2zx0LkRhfCWbeH4Y
q4yoTCxP7KyyqJCbApPhqwKCD+91oWGGv35aRzRLh6+nm3vVX7ERsXWtWyAMTBkz
teZMB5BwwE13XuIbVivnTHwy2g0U262AfojMRSRg+KjbU5pjanCF83rzZlbV/lKH
44FMQnwmNET2WonStK0qH6pxyVQxeYGn+skt0s+ocD1vIFIW5VZynKK+FP1CR9mP
nVcUsszscRMiARLjuGiWlRHJliODLLLO6iZXrwE8wfVO9VScwnhQu1IokdsSFPFT
WnUUfow91r4LjBzxgwFart2elO4fhNzhlLJ5AVGplZ957QIeKIIKVK4nj54h4aDE
`protect end_protected