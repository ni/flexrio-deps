`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpuhRkSkIxIZEedbxXTuCWkFmvvqGLMboY0l+btheJGv+Q
W6qZwT6tMv4md50i092Mag0Ri7ihFc11DV5EUOS0ohZIvjB2P0DhLT/6l/OOtUUi
AoqRp1EGNejmvvmxYtgnAZRVQRC0IJaPaoMW+ePobwvRQnXmRhzL2yUwT0uyV/yt
tN1o6zPGNTcL0D1jj8QPECduho3lbpclebyx5Bue5d2ELlDNfibrsLj0H8zPvAul
FRY+12i6YTMU/JZ8/YoM4j1oKgaLBo/nPJAeGrk9upm0cjN2EF/+445Z9NHIt7Df
eTz97ieD9gLZFJ48qXJDRLnjAh7mphLoH+TRBJSQ23Odn2i1GsS0kwek+CU2MYhv
b5LANUjSRpLejmwQXNCx0bTCrO1JXxfWcdrxBdgSZaXZGnQut+aDrRO09q/bCb+p
OO6nKe/CI64J9t9rsIYv5vMabcucZd0u/Jst9ERuhkq/fwwOXLrN0X1caEHN/Klk
nZgayVJbLB3WnZWQk3XxTeQmUehgXYaO5Zm7mPZPEHy8l6BYXkrpVvQ0DUtl/Jth
D8Dm7jsoEPwY6pFaRzH1ROuLSG8UMTG6oO5+FeaBNGN1hY56GBunHgU8tfOysCRx
A7icM0OVB72aup3eycaz+7/gOHa04V8jEZ1zZ3pLDzwONXXXHaL+FN6+uywfWDcp
YdECq4LT5OuSSlbSoPPLPZgGS5kE1D4W0hZUWvUUZktjYz7g3PMmPSL9bxVaa+Cf
0bMU8OvY/SBJmHzcKAj0DtfTtcMBLYgPO67JBbl8ifbjkehrkqR9481B0G3f8xdO
45TxPRr8+jqorIVpZTfmZNfJKKCYCcp9kvSlPNTBGm9OxFYLYhz8khcXkT22yd1V
2TCLpsCEIex40dSOkrICjbcVkp3+dOwYSx1zM50G1qHSo5W7zPXYjYH18YhXINrQ
dOq56Eq7fb4GvAK85IBDCuKalRJ3VCbj/DHRjs24A0vMgzNwmyP7KPbxzZn/thLf
haG9mtpXceL74a78FiBCy85C8hgNGSOEd145+w0eMHjlENlWWFvYV4Arweq0bFmI
GQH+37ZCYsUqbg51oOPNCgNGjkBrdDUkkppkxPUXnfUNQgPyGTSNexvpgxgMIQUD
yMD06Bmw0qTe+K4l2Sae29dzAfMyStFpWpUVfe4mR1XBajpXeyVQfFm3RB4ZOc2k
Sngu0XQ+sxjhHbml+GM+nBOIX64ZB1zifVIX0AzOI+NHGwx4kkEYHrUUd9xJeOFv
0vtHAauJDQ2PDmaw2RGEOnEyrN0XucD8N/s/xiNqy7xze5PqozDOq5JTIR75S2Re
B2HIBaX0FH0L9uq4QsKso3GLGry/XEeLJs1vvO5MVU08AW/kus2L4VtDV07M6noA
IQ6GRM3x4o8TPplhOwvXLp10+LYzOuuM+amBrkW8XQNAOQ6tt428ggM7Dm2XUd3m
AR+5zB0NihOodK3iwEXQ0+6TjVN+TwWpY8rePce2gGMHtxvNy7Fnwk29icuetPhj
0pIUJYLfyVlJI7keXeNDdxOo0EgImevZCQpwyHRBgxtQEQONTD+/n62UOlK5yyuM
LnoYxBsFf3O5n8s1cCW+/EF0LPdgNwvMqa65Yd40zqkJRizeJKna0AnHz2/dh4lR
eUw4hmBbFeBSei4hFojRQ9H9bH9vza8VKD+ikSwhtkbukr18LJ79twV2kZH8jrUA
HkhHbaoht4BVXY/uTkMG1yGO/4z4G+tgLrZ8cufbB8K5qjR4U4iW5xz3o81MrouW
2kqoIqpbElTzucwj8ha9eTQaDqUCxiWPC0UicJt/r7CmbUUQ5x8aQKAUT3aViZIn
oJTe/pjKM/fMd7CE7DH1lM7P1v/QmjM/3kQ/4tPU1RrxJKraUfuA5Nx2uM+ihHFG
vp2pXOMBrEI3OF2dc45fs0a/mBQb7xElugMvf9DvJpUCK3ZQkIVxyxqMOrxVSeOj
dzzjULl3EfgIyuFG5ReZFpp1duN9hCTDhT0okwgsG0ow4uYhQE7TH4WzApWHl+yn
NmfayLCpMVRVuJxiz8sJ/QaXXcN7mmpezyzQK7d+Zt1qIbM1jDBU/c8J9SXa5fbO
+Te6d8BkJsp4t2EkTodS7lac5eTgxqhli+jy8MhdhH3DlGjr+deQJb+OK3Ms23TA
whrLlxxrJTv/2LvE+0NCc4xGX3KSM4r9HGuUeH3lSQA1sAyoXbqeW91CrFe3ajdM
FUHQ7RZw++Dj4qH/3dJh9cGjspsVzbR91CT4QJCEfZcZS/oDD0kBXCP35Kentcht
H3hglh5ldqu07pYqDFcV7x9tmSG1IVqUtR29qvTUU1U7Ey7SoTEaXhZ9eT1WxVaL
KRnyZIMeZrNoL/XJ5YIKrK9E3H6kr++OlJCL33v9Hdg1wbErgIHasRFR1o64mEoo
s2SAoBexiAWTmFzH+rLK7oZp/lTXEDiAyQ2DHNFsN1c0i2qKJ0tu4+X3JrrK2YVq
GnGL8uZ3gKwyQH/bDwtqyQft3mfb5ER1ShrCNmwNUxdbkGU6RqLqowR6HyHEykGY
Hhmklx+to3uttRk9oj8UijuQ/C6AbmtD2lk7yjiN0rjJTReib+CKIIyvQG8UvlqL
8NoH8YJA9N6wRumHx4hV/SeelVM9q6hoKTodsdk8+gLZhgxlAoeu9vAGkIS6fPfv
10qLByEky7ffYYtQXUcExPzAKddySljCRhKkuKZNHvj7LnuSinCDpXLHzJVpGHJG
p4u5i+dT9FAhexKa4qbFXmB1U0kILtoMNF/g1tJVwawokkouN1WY12Cvt7/t9m4x
u6B7Af3k0eQCgm/PO8H+gvFtr6VD7bTnUT+2ftW+Cro7kIe+mcxqdRR9AVnG7BUj
wDOYSXswYk6mCMs9cF3e4MmhJnHAGHImKkLXJksz4UmmV+Bgd/6uU/aZweYC0PbY
0cV9Mm65dOZTmWgLXEq8V+P/KWN/fPLKx7gZutzP8gomJLjJEAEWXOlVOYKUWNDA
NZZsifXiOCHiforNMpj3i84kEdCLxOFhTCMHSFnVvQwMc18+qTHGJClAkidkC1xq
E6JXYWHMqtTF3awiH1YXNfsFIIUPOaP1FlIUfChNW/LQuX+0BNQLBfmGWMcRkHWu
3tBcIyHkISQdez3We50zguGb/nHxm8de3KeeH/Vtp5kwDOOScq2kFDhopFB+5KSy
gJi/Gu0ZPoHl5FDdyZTLTN1HqJp++cd+lTHEjWSWO/i8Edzj6cNFiJOQ1CBqfubd
EHfJ2PFE5lAXb0r0bn1EJssBLUjLuSjLW4oawnp3tDrlHL6zMGO8Nh86uHsFFsvA
yPFaTLYbwV0YuiLxcYfghDoCPCzc9uXmm8C7rNSwZcgEtK5s1Szwrc/gjL2eFhNW
S+NZ6PUtlffWG4fhenAIHuT1pIWeyzC6ma5k3ffZ+xQyNRLN3/2jlcTaHYg8IU0R
7q9olvIaqD1BJfAmkbzwMRNZnTUuI+Trrr7z2KPIJUuvPoWBszt3y22/34aFB97j
/zUGDpnx42BEOorUdg0Rxnjw0dtWdDkfEgZ0nv9OhPB0Ja3m7b1rpeX++7aCvJtL
2lQdtNkgQBcASVOx9qdf6hPXMRmr2UMukFzAeLLrDC7zl5qkYok8Eaphvly79RXB
ur1uBvSGCtkrzdILX+DWuNOzHk8xqByZNV1qL8teReQZn6pnB33LONVwSizS5Kh8
qbhmGt0Mnj/Ay98oc2/a9/hZGA/HLNTBqHLkYqr62twGGbv+/vdR7rq9CeHgj61R
hwGj8eP8SyI3hDCtapXUXHnTvVcE0bkADKvEE3CV4+Ph+eK5tteUsjAiVHG9vY/k
I6ifTv7i7NGoVzBoi8KtedZZZwbUaGGBfQEVZvfrxMFFA7W+lh3ioBLvTWmt++fh
9mpZRbLwvg4k2YKyw94UlpCGgGJSbAHfd1c4B0KqHrhxMMi0fnDGjfgYFTQwmNWF
nAJwWx0vt8COSN020LMlje+UXdN+25CDZ31IXSreupfbmeu++a2+JQ5v+mkn9UhB
r5PppjDLqMBs5QwZ149L82QZ29VQKNtp8GaZwqStVHacgONreZrczbVUq9NOtoG0
ZP7p48gEvPEj+aZoKBOQWrAOPOg646BNwyK6vPaABXF6e54ADn+4vAaMgpDpwHvQ
LRhYJNzvW9f5s82eOPRaautgKaQCw4vYxADLswfnTcmfqM8G3NSE5HRnJXU6ntfC
2kHCstFNDsiq/XxfAtZZmt8fgX51NneqyL9YmMgzINgzEV/IsV/3CHQpsrtomzMq
MLAWr7vZdplXiz1oaMjcw/adY1ithaZO2mc1Bu8/D4Hd5xYc/M/2uy6GvdfXVMT5
pWPDdFG1Gs4HXPdVVO4n8G7n9iT7LIFCiAlGbkpMhEWClzdN4KUWHTEeDc8EhTyP
ZQJf/vypAOM2Ty8aLQo2QN2ur5Xr5u8a3XstVkwzUhRRwxEIZVIhLLss/XvO3yyZ
WhjKy5iLVNgD4ee4gyutDpRL3GB8jnbi72q1n+TtbMIxq3OahJQVdcX3aMaxhsGD
i655k7G44IfnCsb8Pvz2NDOPwCG2aTQMgsQdfIX0M/KNlbgsnXq7OMSNRjHxTTGV
E02bzljs5NjduWWYnawGluWblPpts1SdDOmLE8iiPIaHbravtEkeSSn7407iKUND
rSp2wInAlJn623LI5IaG8ime3kMLOoTR5G1w5uNbFLq/8l6ztjZpF4KrkRY1sCac
2WjnLsXbsbdbUy98BlJSLiKafsJyOpk39ewlPGPCNNaukOcBIaiwLf+Now+pShZR
wCkuy1lI6ON+h1LEKcDomRXXdlX9BA5jQH3mYzXZQHtfgK/tVASrqbNM+j4OiI14
IQrHlMomyBoEY7V3sF8GJH/X+XNcciVCaQMUDHDN25va/tyOK0ICC8sY3ClbibZL
dEdaH0RA08lM2jo0c1LAdQkiqNgIadHLt1IpwnvyWMkxXxG7E+jGfBIPeId2eU8+
wYn8j1TMtAzZLmCwlQuckmUAU5WRHS3oKuLeGPhmcERbNLyutGjozBo1rtzKWabx
OShrlJKdPRxJVNtL7V/DJv6pXG6j3NGJpa62MmMfIAikvBg1TyWqUdk8b+LBM/E6
eoljO2HXgO7QuUSfwI+gd+KZU8PAcsMdTPNgalHpL4OSe19W7kz0ZUz+hUpOoKOe
BYZPFMDSng+2hERMWXFQuU6fLkwu8QpKI0LSyBAw0uPDFurw2GqON+zohR9fyw9B
nO0ou82mu/9cL0zjcqDL/a684kmCCB5mfnY4sWfgklGdgkne0+POWydyoInEKeC+
H8n1ZEXuD51R6is9M0kGdiZ25mLAOr3b9bUjY6+OYvO6nRVjmxlD6CMFISsb+HFL
dYWx2nKaebS8Ip9f31tHHkgBWUEaN7RDeg4r/6jp48EQ0Z4kA6RV9V0HB9MpCWt9
pXmZDpJ1ic5n8KMWcoE01tTqCJ+u2qfA3uQijOdq/hSuUjAGnIneGsYdxOtts4+4
DdBOXbqmbONNjnlAGpWLxQiWJ6Q0n7ggpYFZXDy333f1hY2K41tOsLj642Sl1+Nj
vMULukX8eg++8SoPP/hQL1Op5JB6I1SUsygAVuS106KazxbL3F1Du7veZy9PQil8
/tAOAIWokW34JyjhlQcCwio8TV9HkyO//jejjjbyh+Jpe8xMK2XZ3e1PjBmWPj1v
`protect end_protected