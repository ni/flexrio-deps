`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzkZGdUrjzQR9gfRaWjj8jjIw7tUyZhisk6EDDoSkXbk9
4KuPQR5mCkiRfz3UIhipt+XyNds9TnWH4yB3lDTDV+QhwsqsjXEUZ0oF82NSRxqo
aikx4iGrBvyaOU43YzT3deLFbAUdBCUfXGjh95G93El/EBVT4CjTGktRgWtZ/xHt
LF5I3milXrP6M1Z6nrRQRMxAyZ7PCvZymeYeI1rg5HRnbccqWZZ3y0ZnM8gtF+6T
th9j7EOpunZU4CmI2ysa6ZFSkYCrgUbYKCSmzV0nOcJDvwVt4gg0F8T/xYV8Ya8a
Vv+X/Eeehbhdedk/KPw30VKOdW0dDshLSrVN/1NEXoQRI6IA0Iwq+RTGLQdoXqLr
uia2XIFyEZD6oIJxq25tRLQAVFV/+2y+XlOXiukTSQlns8gJa0hGBv45I2NMPuea
za34aF4wAC5RCN2ZGaY5Muyp/WN7Ih6WgFQocB3iTYBBn0np/SeBp5r6lgSRYk3H
LG//FGKe7T5YNfEDAJdvGebyqQWpPYjFWImnq8H6s8PnmxcjMkol/dY9bkgFUurw
R29PVUcaXJrAiyiNIToEOo2oCA2VLFxeiIAK1B15nY2FQ2PgEv3ClozXak5Utush
C4loRg3R17sO5OTUKjoDxMDTtqvQ4SSCZ6mBno247k9c45oCcKrMkXKqilCwjItq
ZOFjKA20biCZoj8DbMzXB1Op1O09o49RKm7L1WkM0FgqUXX2czeB7CWxcwqdqEoP
zF2hjy9azecoYrft6savd1vO9rOXC6h/af3jShBceU8pL4Ysob234lQAa4+aYOqg
AvSMqnEbzOaKlvd2xo5O5A7cgmAFCAPbMVuolNjL4cTQyndoBqL4AWb1Yo9yg8JI
jTcDvZKmA1rdaMnhWrJx578U4wU5K4T4PMQ9+HgQwNNSny/ivGIiNFuZutSlcsRC
rb7N2VRN5PQa9vMom1Rlv9dBhDndAS8RkKDmuEmh8uxdpyMSwczjo/+wefYL1mCZ
WTYHnAnTWTvRQBMlOiiVVERrK6Oc20uYZBa538LkYsaUJ09+/5O1PNuSXnnR9y3Z
ktCV2aqQ3wxUQdGkJzRmFs2jT0xLirNAyJPfl4ONPvWzoKVgR4uDDc9tnKWg6aGf
T3ysiAf/kDSQgzFxUk8Dk8qhROv0dtFmRJ+kHPTKBsHHMS4rYYhnV0o2Apsg7Wng
hcir2LNtomcikhQw8cHjXDoqOD16QUCYAlUiWvTcT2OoaIWM/xVfew2TFQL5bHRU
H/I11B04xYdUiXxO/FB9setwcKWxevm20Fi8cskgoZbX+niL8e+uitvtNLxuRGzz
YwVbsFEvXIenhxoh9KxFrjawG9Y/vuxc5VOvoOMG7mw/jNwcMi2JfUCM4pE6vKc/
nlc27yB8mwhxET7ONuJ3Vh6DfOPhoMujgUVDF3UTvXAVYExnvqo1HB4JF3e2TeRv
KGMrAXnBOlP9s4laBhMfzsg4f86KtDhTrD0Oz5qbHqO+6fCpufW4M/wicJY6s7rf
V4Ek5eggtXEQOi4FyPA5aGwSjYW9qWHAVowN7i52FVz//NN8S4r5q8R1NpvoU/lk
D4rJt3BpSFcFgKtLsTAG+9jF5onSPkn9XoVydmM4NkCl/0mypxkflCIQyU2VwH6I
BXtii+KQ+uERtzumQedE3avIx5YXUdql6iwn6ZJDUII9/Ab6aJsDomfLBeqjlBiW
x6EEddQVSj0EN8obUX/ycPc9PuPOpgo6+jx8ieGEyjQaqFIiYjAUDfLlj/dNSF51
EDZrV+bGcSYfozGv2sOZAXcC9qa52eAE/uYovbbA/MGV+fMtER96ZDC7XTeIwa0I
28/QQyAx06eLgkpyNKqrxEmChcuGBFKlLjwd4u9pvnB3PQDIdvzwXk7n29pWuRE2
1HqJdORv1UzoJgSW0FV9w9N0NKfPo1cXsAwP487lnJetAuwJFpXG9VeLT0RYlBML
g0n3HHtws3djLmw6LILZ+CM7FuJKfM99wAzXII9OOKd7b3si2mQG45R70nHEtWsn
B9BSUw8QWuNZGJaLpel41JRw0Qk/cK71PxN/nK6SrcvqN5KNhJHal+oQBOT0MlAt
YweTd4MmtIex+keZa4ZL6rI9S5ZcM4AtW67dBbEkO+LNbdMnIGNBiUtmjwBkMkOm
OBurt0Zv47IegJjbabeRYQlSCycCN0Pm9vjpAXeCPymYikLEkoNUptJnUVPqtbpl
OJmB5GONZ0brom2BrpFDoWqmLNKn1k4AjjowhDOlCWUhOD+uzNaDwcQzMs98d3kO
gFwT0nykiYdyys3NY3uBFZbIGh9Y3BHj/jl5caLdoIPHiCgQIv4Au7sswO3pE6tI
sT3HnfwCtj73Pv0mUrsjhhK1EylKil4Aw2GXf4qhHb7ioCwEF5ElK1ORQox6rq1k
2355H+hYzMx0FD4WwNMMubLZ00t3gKShphuof9BIS3p65RTFUvfAewRPiA/f+A8y
pdYMG9OAS5LCBFBAea7toVF++0mJZEv8u/ZYKyci+zrd8+OCzK+Zi9NtyqSxH+2k
4CoN6h2gFDPlC6dyiDmBvSmoRDioLTl5Z+reFkbuKOmMIOxMrnfAo2t3ITX2CLjv
dA3J78ayikrvSp089eBITMJj4HnP3Qdas+9RmyON8rKLgrwMn3klk6sIQ3qdq2m7
ymOJ7vfpb/buw1a+4FmJYwUkAJSjsiHjB6vIjKOGv/vcuOcxLzbKVZ3KQ0ImkJ9E
Ni/MsDIz7C04uTR4gJ6YytAQujUJrFWv+7hH2RNl1gXji+IkCMtc30sFeo/VGvZh
zgIzw99AgTIsaXeZ6SV4MAAqbM7wfD33jDpxQ4Tl5j8ZaDNMt6ISXqrY8e7hDiU9
hSZO9K7ye1TYKvzBd6Ifp1WhYYapVsK0HomMJ3VMtPkB1MLMRiULppneds8PPotE
o7vYZOqcAehe+EaEaA/r0em0qGtO4U8MSpmM39TcG2tr/AS8A03vnN23pqmVUAWn
Zn8Tlkm7q+x3yXzeMcml1b+oH6UVMwRr7OSqWA/FrND/Bof9BywE4wNEvBaH7XpR
X5/q0/NLgj9cPkgi6ESQpF93YdEC28F676GDu05jGEcloc6oO57IlzXlwyfRkrF+
0DfnClrigER/7QNi/VFB2XkBrD8VmWXHDKJNDjU9cRAiwvh35s56E0xuGqAO15hc
xc5VfHbKlf7iSf9wwd+WYcpdYLZ8oxxbFrW4GgXbcRQ2GimJeqWDmNnCCduazebK
opkUjzeMPtKDANge7fPgutf2USCoUdCYpJM0EQUEnSctSkGK71AFtG3pjUf4Enom
DT4uxC+Pd2Rzxv1gYqgASi2J3tx8WyKnT/HbCltnHAWsYoEFMv4W6sbQey0Bt2rn
CAda+esrXF9bKFcAg8lH90iNl5qn4wYWgsvZzF+y/yRFzMl9Gn8mTb7hdoNwHX/T
a5aZVjlYJjQye9rCisZrxDq754I1tk2TGf4Iqd8UWE+7Cle4Svrzu2m0ZUfwo/lc
NtEo8XCAU7LfsWwn5pRqNFZEjFAZLvaNIW4ldHPatRmtSxIhLAe7Z+urKaXI34dX
js8nLiSeqQ6hiLo0bye0GS9lLnTW9ojgC/6kJkDo9sg7rOuTCn/xCkvRoLWSMC8N
a4DOnQpm4RcoOyw2Y6xjhcqqrrgM/Knu+zcA1VGmedLEsY/YK//ql0Lhf3QBi7mm
KdOHk+E+KdIIrZJyI6vYkGI4LRT5qJJ6FEpmGAti8mKP7C5Os4roDxLI8Hm5Awt8
OR4F0EB6x9Y7L5RzEnPsyCIG59qMo29AA2c8g2iIL/Si5Ob9Ct9XbB18qA1Cp5CZ
TAsNeAv+KRJLy8fH4+PPhM/SG9fZYFr33XfVxOxF0uKSKQ0kdvqpbKvkToFe+Do8
g+JbxdjLPJGdHvQjRlezH8d1GOh6Q0L70K1HBbBGgY5u0QjApBkwE2vhw81TYzJc
LR36XZ4pYK+SrrcFyUuNAr4yPhD+Ei3M0Y8aeBD9ec4rArRUYk9VD4FemMK2ENey
UbB+hRDSci9T8QbsiR+9Pn1OW20yNS7A0XWca/W6/anApOZv3SCcGYLy2kD86NOU
IVfwUnhflQvc9Wa1DcarZjGOA7iljhOdOXymzv9T+HEA2jvSl0MHQx3viFNQ2Avd
gxXMUl0inu+1f9Xc9c9RWllD/fUMXftOR+sS4BTG94i8giJFP2yuw3BOX9LXoFEg
nM1jQJ+2ualc6EATIAsjsNExQ6/SSt7tgmvwDyl1tV3ID+NYwIDK7RsWdWRHG3Oi
8YtCbAyi0Z/zPWxo5/ajKcwWCFeDS1uoM9URna6xss2Kgw65hgoVoVIFwCxzQheK
xUmtRe7Hz7YeX/DCizugyTFbAwqJ7iM5InXEK/ncxoU5LoDtvE9c3+PMtGST9nDi
SY4bJMojrf22urrbUjTc/91TNtNBxFRg3Ko8RiUbmTU6HUBzlrdOgihLl8qN6mbL
ARcKHCJscJCCKiNFZMHPjSjEBrtE8YmUr55gxgMdRnjtQ9Y8fJUV3xHdHIW3KCNk
mERekhTHP2F4Y6Hylu2s0Q4vvzRZZsGhEvWoGD7XQ/cCqgS4rmM+IeC7SJk747ep
XizDiw8DZlYQBm5IoxtvGl9Ih8WwTJznaHOM4pYUANsx03a3CyLgqAaTomXyDSc3
KFkKNaXPY6hWNfQMX4s6nfXAwWfGS9bKGG17As/gRnSYy9jrix3vhd3W27N+olvG
HSQxi9zXMgNONWkaR/l+QtyjmKkfPcfDViZKckaER2OjeBKWMKDmnOoGuOlddDoN
BnyfpFHbWgXNDi87Jb6v73tGmrCPsZ7OoxhCWrJpEl/AW5sl96+Kkwiw7ca/SczH
yASY6puYhpCWsDMIQiFAcBos1Y4PllY6CYDTAokbrWRVvWuESrfQERdF681ec3fL
gUVaB+B7FxuaZOfMIy2aBdPIWfZIddygcfMyAXzZrh1owTq6o1VWcyWsmi6DcHn8
aEUakwZFygzLfI0oGyc3I+qmpHL1Jm+YkHbj1ZuY0sqm5tjD4e/d6HCswUZ4mpNJ
UmQepTkNgFrdN9m6EWr7drJhZ4b0g8JEhnvLTHS5ap9PJpUcy5HjcepXNHLZAekD
oSFI4k3ixLjD4cWHw1p2OXKOCfcmQPDcqXSKmBb+ViQEy+1Tso5/EQfj4EnSipDP
hhxW5fOKL52NcZwghfK1Irl+Whc2NHwt2/5YNmlMYc20NMc1Gv1jigI4Lc+QZMAl
zFL9g5ww30PSOZ7zDXWNrzlXHNelZMJ1z3vY1dspjJLVlXWMqAmq/tk3cgAfV9sx
N4OsGhXtzeND2fksWoVKKCfwz9ioC0Ie7u8XVKf3iOzNeI1zkctddEBps3Avf4+M
KGL9mz5i+w7BusAaBb9QNlDG4jvgXVoFXUJWcAQ8sWFAC4Em2z9menC2vDZ++9kF
VzpMruhrPdi41StSaflPEmqy+g9m6f3htNIR++jCwbwTskQuNff4zMUaJYEDXCwz
ee8Edb4FLQDDy17tQGiQrdMMY/w92/ivC8aSTE0jcczWVyTgdcOAiTCA86NoTEwu
LaNVzjvrXSFaj4kSWThnkyDxYB3njzySjw9sAzboVhH+JKP7pIv5V4ulQf69Bq1+
FT+9TntSgWHtrhncngalcianSKiKc5f3AWfQ1aAH/V6tb0KuSajgDgWaGwMaT6ol
h/+aY7+cQSXxAdlavA0XanBA4zS4FjhKf0lhKfGCWg53fwMtBWGACY4BOve7rsOv
weTDlSNpnXSw39+zHVrBHYdcvG41HWDDEtKQ9mtbPjhMDym7B+r7oPNK+Nlw7HfJ
B8NPcZvkZyE5HwWukOR7s+qugEUNP1nLwUWJDXvWnvtwrNuJV2M1qf4CZQjss0TT
7p0bzluTvJWe09d1zOjicjsoTDv1Z/V7qbtMDzYBBXrymMMxoSWLRd9jGXyTniP3
XwWvUqyXAUjFlGhavhzqxkp3cwh/2lbdwsEp74jNJKsQqjG86AjV+/LKsGIaVsT+
dd4DbA43QJEKhCKTH8mXNi8EpQHrW7xQD1y/NMp0MNi7J+tKPXOJ/kLE5+5o7xXC
SEQPX8CVmXzq4t3mh8t8HzJRgb/NSjkZJvRtU+2vM1ljD8NnVP/nTQvgJkAPAfhC
oLf8Sy2YoFRYKTS9PLeDwk363qwISgaMFuleLBQ4J0ig3FyICorRDfsqZ0+AFX+k
2RYDsZpTnlHxhWdJWuclEQh1avxIomWKkldOXtDQ8cwOTAUN4A1/18Su4Zm0hX8M
hCbzd21JAIaywz+7iR4hSSMyHD4JYOC1GvE95B7DaAoy4STYV4NGW/q7VSkQGQds
7Y0SLSlyDWzzSAYGJCXUMVw6xAt6aV3tWQIPSSdTVudORKiQSqmayb2zFsUOUBmW
BI4cH2sxiPLkDo34vCzLAELV+COcUwrC4kK9ycvrqavnlrbSsD3J8UcDQfi1+13G
0noDbLKX1cBbz6ostp7YgQg7TIc3gZZg2XocGMGL6AceFUNq8JIDAq9YaV7WPPk2
vcG+ET1XbgqM02Ow+awGhSW0Ssq/Bf2vWbwg/Ro3RrA48y5+rVxnSWPc/FJkMI14
76f3R+lHxofaoDNzXUNDZQyFEWmTw7Uz9aX7JmCy7tX7uhig6mvgw16+LtnZ3F4M
A78O+tyUbHH2+3xAo5GpHVOSEAbCygHAfl+wLsVXpijr98eusYheW/rXwcggTdb7
y1qzXQDxsNtMwPb7bMl4hdFgE8LnYUkASQoE8/e5Bsq5ZSq4FzOKTak4abIqmQfM
wS0Ec4APQdjpI/QPk2KEXFZah8BTHBVhW2e1h57H8EH/DS7yJ8f+TD8OtnteMeHJ
weqKdup2jP1um69nrJSDW8dfe8bAprbb/d1Uv943GcKo10MJ6s/kYIpCW5KVflgc
+IXdmuqfq+iYGdbmPxer9wknC2Hl5q6bvlmLR8bZS98d9F0M5MzrnNHeB7UtjlTN
a0iD5PQ3AwT2ggUE6PNS5VfJRPWtHsw0hu0DzmwDaNtRTmPFh9pskVtOmrdA0OQ+
NMZNI0XIteuZTBtNKrvWDqAYn6zaDbKKmGnHwFDRNbrnF6fnZ4WhpExO1AcVDbmX
Kkf/sJbNSVNvrjzlPORbYYSRDaye3RfN7D4V0qe/rx6es/SJOYPKzgKVZJ+5toKA
mTNnfgFVzRAJaLw4f+8vYC/A8evao44RJ1srFjMxQ2eHAGp++rFjS+ibnoQySIJs
trXNzYItRihKZuWcsoArtlf1q9w3oKXl9/25nktBgST/qqX47IuOCVPcFHJC0z5S
V5PdWrkkPAIwkA06oWChgzRhPoWBlRqsQ2fOzlgO3AMemB3NLrC2tfSfTEhivtIc
QE1w71eF+V2utFUZO/fdJvTBoOnKlRvN5bLbOQ/kaNSwEL2BjB8OMItL6idrQ44M
uwjbuEBBwoZ3AK2cr85Dcj1+6clTxmsAyGGbciV8VVcmTAq6xdNLGH16gqElG23Q
rzCFULZX+ve+CdkGZZItuUEcB0iFv6ovwNQuV8S2LK/055dU0VDp5NvnxyG4XGvx
BPlBk2WShWFJgt0Rq0OB5Llq+hL3T0iVP9uf0s+krmr7MH1Q8RneaACViNqt0MTy
+Qhi1WsUX1TFvJ56z+Zafc5DF3VJgJ7gK/k8XP3YBMsTXHom9HQ1Dkqk2BN/otu1
B5tBKmsGmq8bvKMaRu+2KeUyQKg+SAu+8VC55OSaT3/OxXbk+GJKLc4L1S1VGwW0
6uGYMFlijAfyNgV3TuWnHi7JBfqViGsr1/43/elOl/N4vcmMB63rOCg2qxrZhHdu
Y76SUqT5J5+F3GhbHaYU+8TYrWQQkI6lrrIddfCc5eRzGusk8A/9qz6v0GIHhzrD
EFFTRAo6wk+9nj9rAxeYMru+Em6+dqFo7qrWiupVA9s00+FBSrcFkTweYfrxKkP3
Uy2Ie8qK28f4jcnrCTkq+nxPnJ1bg9dDa1i4FE/cjz1mYc9AibOZFu+sDs4BD1tm
+JcQAlruuiiG7XniF9aVCYdolPbA1Bd9mUCiLvExShtgiX2EfECaWVXxK8FjmXRQ
uGZXzu0tLoZmZskkeahG2QDO/uSiVy21qvf36+uAHWVvcvYhmhW2ya9D7GopP2qp
X2Pi54rfC/PeOFk+u0R8qPxfdUxD010txK+5dZ+L/yUGhrV95z8HEBerSJEyJfBB
1noD2DSzoW42zQYXllRdoX5rOzdGXog9w8G7XTERfHMzsi+Ftw6QaXONjAx+5U0D
jzvM/pDVch5BwplO7wwJ+L2KvJlJmroF+her01M77QuuqieTEmzP6SdP8XpqrQnp
NHJlSByLLH8hVSqgBz8mGO+fJ21hP9ywUJhLFwkcPvYDiQvAIECcecoiMrtaEgs1
q7bmHQldI2qHvYsILPq5QpA72+09tjJVpnUmxHptVhSFcbfiuegbqdtQ4W8tB9l1
Y34u3OuRtKED4C581RfGtV9r2+BP+awXscvL3fAw/br6+si3cXzafV4mAQfl7aFm
ayGqipxyYOeTj3eGWZaQSxTylexVc3NIg6u1bwLj+RJ/7r6HZ/H4zZS44pg75BlU
mp/IET/PiZeulPOw1a4HnSr8seckUOUW1ARth4ttneHAJZG39nqN/BNdS5vkTrLW
A+F+TgwY1y5BwE5d8ja9NqQTgeBbztxwaK49O3eVZIlipXCGyrgsU6+vVPOLpC8b
+p0xdm7grWpx1K0IfZ9DmO+9yxupYwcLCmzTJ4W/9jRi5Tt8QtsAvIllML8xM8m8
Jza5ccp40HTgIrSkDXRvKprjf3cEuFHa1lTWsMnyw165jkfFQAJeq6VJqVTjsI+i
TN/knAjQ5Kbd6tjMoQuMu6EYMmmM101uUM9bPqGsx62Q+1iH4zGuR/0OSlDeT9ks
0rc+/jINZf455gTQlMrrO8g8y/DEOeKCKURaLoGohpTgxG2yUS4jHMwDU6td8V9Z
o/H0/md3VYCkZ1tqX8vB09E3JpmdiOhaWgJbEFgESzca0V647wRaJLRtTV9AavMq
4UMNwmF2Nb9ny0d9F4xgDIGTc5rL3rA6XcUINd4DyYflxP981OEa34CZHwXJaddh
iPgHneFMW71ophxJ2LZS6XvpD/iGy2BugFDBa/di2+oRZLmrclU3xwez9A2RDB1a
3UWx3FDpAeHalHzQ+0ulLnHt2o11Hq/ZpTbONyCZdmmaHx1oMdm4q3xYbNqMbgf3
e8CPWOHvcA67uCDWv5czwzikAbt0CPNgeZ83WvNqDbrVDLMqOBKMqrW1HqWBdekd
S15RoGxng58Bch44sqgZNvbiPjn2cIdYzJqgmFnZyAUn5k4nGhiI7UOeVignm7dL
6eRE0e851D2KqpjP3fU+LlnuNmVGfaxHKvQWI1MN/BC4MofOMOCVoINh96wdE7oA
2nUZWThwq8c+7WhwQ/x8ViJY2e8SFhFFEyNk7A0sNKLJUP+HcR/E7RcctLPEFTg5
q7j/AvfZ1INabaIvRq2MQ9aWMCZ11/524vpKUHc5Kb7nMPxOREsCPvxV6ZTDi+gz
96Dwkd8oVzR46ZtfvGs3lYQbl1vXDS2hGOG1LtPEFRhQ9Nqa+x2RrniZHBe28Qa1
lWN+w1K4SRJ7LjuGXapELCvlMwQNNnq+BJrzKoVN0kxcBnAg+ZtItIJf9ni8JniI
WR9vQi9rsQd/c8JULqRAiZQlLGJAYp5WMN/CdSdoURv+zC8d0qjcNMP7DYjTTaIm
pIKqDm74RHFukCqhslXsvZLmpsZ0bJ821oVpAqAD6xjeu0Bjzz81Ju6Zgc0Dg7Yp
BoipUVDqFEZf5BdOndI+d5OfrE6vZ2rSNkffvVMJNHu8oYWC4LAQdVRxU6zmsb0S
RCPrKyav+NkkA9n9WsZnV7O1Gq0mtjT//u2K5bHNGjQmT1S5cxyqAw50fe5cQoic
QTamwaWItAFCmiX+IGIZsXgoHO2+BmAc1JBijzrLHMBUAxboXpACBFbKPvfaS+Hs
jTcY+r/s5gUtHQUx+KyLRTa/qgECbgaEuNOoCVru/stNBOREBph324weSYbU2kqS
gY37EkYLLyP7BzPMPwI31FzPHLc+7Ika2NRUyOr2LFIfYnSq84LVYNdG8kWFRzsO
qddtYWRMrNN4CVTU/ejqALR14T8hO+qQq0lfEgLQDun3ICF/6pMP7as7XPfE6xgp
pWE7WL/yOKd6G/3kW7rWdAf6AsqwprAJ8ex1wviGEO9KJF7xJsJTCeoL85NGJPHz
SxTmc+drI7qGQC3f9RkNTCA1MuOJLGSKCrDoaEKUTDUNeFwxP3gWcverluSramgD
pJKptOxD/6rASdh8WDgfulqMD+dPIQYqKTTczD41CM1f+2yDbEpBI/ZME2SM9HcH
tFX17uj/gxeOeVwQ9s4WUmXM0F3ix1A82fo4pwE8kwD3CpEhpxmFy2+nUDJMSkXB
sLf5u/qv2F/7ndZxRDwCejSmBQcFt86YckinJvHVNhBfrhlKMLZDRKtJuig0E8YT
7Ese7g8aFvVcH1THwS5eYb+f231Q1YMUhuF4ZkegfXKiQ5OeTqpb53bLLfChLpN9
HDvIOQFz7RuemLyK32PlQpFrzFwCcawoTDWG31c4tiuGhNFtoqEVfzKoFW2jCPZ8
P8S849jp8xrCG6akTQNXR5jMOvSdyGX5BHWvgWWezqFkJg97aje+GbSi7UkqMTuZ
RoZhFH5UyNC73n63xU3sAPUc6wX35j8ykKR0vpIVhJIOm9QI8OpIAeM6xWjMDWyp
dIoTNe4gSgLO95ZCmGOxmteMqWuWY7N0nPqRUMdHdbHfPRj9PwXv3fNYS6Thvg4t
E67k7ZrKc0NHltW+/+Tkv+vOSZEJ7p5sEA0HKEhv9ipDiuAHg7mJoc4ixlxWv//V
zwF+DYXAqkbR6EDg2Tv/0wde88c/CTXZhG6MIH6zTsr0vbHRsbr//OaYz9yyDUiz
wAC553PC5Ofgb1PxOFD+tWMwjAiqGyN8Hre6j5BJzAy/Eiff3zlT/6RZYPvqqeAN
pxFtliterkFNf+GSgq7NyacYkphW9rs8QSY3pMwUwtDDoxkvg6zB+w9gNe6rj5S3
Lzuxrx5YA1H7w2zPPGrfDuKaXlzNpOjsCxOjRjWPpO5K6VefZJ/bGJnWY1nMOzxy
if3YfhUTt1F9E5guxuIDyfCxJqoAhRglq7ET5IYqBZXWPHIq1CALPCFzCCBFLYn2
xryo1T+6fymXLtRpFydZrRzdwoMmb3vvofNEwrCSJauZRkj234AvlbLhGjgPzZmY
uL4aLUfyQ0laRldtC/SjQsOyHypp50QTrdMp8RfKEOgAbQ6pCBDFTAooEp2R0QRP
9O6FcGS920VYmfSXB4Vm5+1KzSXvQJQ12kzKlco8BQyC3YxZDJkPqHFuXzFFD/38
l4i3KwOGRBpKip6kS2I3Hkftk9PQeIhg0JentYAIn736NgF6an9IWVH9nagEvQWB
xKMKp26FEoIIGhPKBo1hWUuKM/re+F/3YczBwAy/uKJsTj7G41v4URfG/d/xc9sn
wy8UcJSJs5GWJRHCHXAPbeuXfqrPQ+jznPJCQJWsJbu88k9RYHL1c065kHCxD7qe
IkCefrxBQZeDSDY626YPR2zVzT1sbBY4SsnIrrZvPjqW8YTSiJa2Agp473ZjT+It
q3wdrnqWgrctoQ5Ok/Mk1hDDesFXmAsP9hlQBNA96e4D0d+lUD3LLDIzK49X9jpF
f1PVxv6NXVHIQw3zU4Rh2WD7p4iPPbBntiIwRInzy27SJXs1ekatpbIyVdO3ctzk
DyKQMW2sbkrvXnIFahdJRovri/YcguZS4aR5C8EGYqprencvpeRQyusi+oA2zdg0
p07L3VbOiwFxEgP0mVsoTdhz0oTgXJFx5HpNjjmOg/b5onC6RRejzDlqtq9TcIk8
Rio3dZSqX8yJj4uVz+nntwHDOTzxW/xmF8ZxRaOXBqe11qSofPGr1k1373ewwDcG
K1ngijfTc7409W+742dFxS9PGNvFbKv4+6HXfQFmE5NM+4R7R5C0VXEtYIURUS4z
gjpZj42iQ38G0wNxOGiOF9LLZ7nc0A8Vrwzm9CGq+UoM/88UgryqHT5zkMSI4P4K
EhV+0gVcrAiQ4QUlRXFSImzqHbK/bw/buGY57jdYWhRGifqRBjhaiWRTh0lYIFSw
prXHrSixnfCe09JPx6NJnDOh8SNi9JW7p82Nvl/l2BwD/8xL6LSopzOBxXwP89sA
YzIyOOZVzo0MZZoy+jmSE8fHcOst8oZBmcpONOEv4E65C27JUCA9GHCgnsxM9b4t
4gxOVFSgRMSsYLEcxd50pD+mK6NXH2mZ+5dmHDl78v5FXkI+E5wA5a/U7ZETg+GA
h+IOTlMsazTYONdP3xMMjKSrhikdK2dhNTjNHlhF8Gl4yhe5sVeGRt8j0yj5jQs2
DHS9K3bE40Ycp0Xsg2jK+Yol4josnXMMPpRgpt+lX2fzJ30nF7kkYqNJN/HmmtEu
bVIJtnn7QUL11VeZlE6tg2nAdFoTDwIQStJB3/8E/4qNqT92DC6vCm/jLSVxZhAZ
cvLrhpkAOxOsKbpqwkBUZEgeviv9qgNY0vqNlXh1cr0awt2z/Jq7WLtmO3NiSPRA
q8/maUCuCYw6b7c5v7br1tLK8qqsBRkwP3pRRqcRBeXsSiaDxzTTCuQ7wIpPakqx
XZ2fefOzbAxJnG/J1N9yWsCi5jBMrBvEDGokN7BFxooYuwfw0dKikSPDYoacgLvE
PETRV/ihpGfsgMdPk3uUeWVhCU0ah25hHy4nxal1+8wUbaVM1wXaa9E6VGAa9GnH
UNIOWJqHtndJZypJhO20CANXRepNPMiCqP7MZBUvM/lQNIqRZ6q2OJEHKjyDCUCt
PP5LWMkZFKSnGBZt6YR266d06IYWOA5cfFEVr1Nnpd3vTKAVKuWh4DhUsKgVKjE2
rhMTYM++rXL4bIEgjDUKtGu/j54eInGeekBcWWCehkbogzycF+oCd1dzqF2tzyV9
4PK3795FcfdESFu4y6EmlRMogeJ6eild6Qo69SncSXA25zu96JsMmbFS0l0mnKci
6HK9JYJyVCixqo61K2OnAkie9LZbVnBfVu9UM2ussq9GnS7mNoIikH+x05e/zsuk
9Syc0cZtV5HdQFzL2EhzfrMOBtmFnS/BYwphSMy/2Yv2XojygdyNzSI/7gVImgxy
LUe/wrlm+ZSUGl5FUWcqD78o0lOOfzoqbMGMCrAzARRB6VjFEH9519gN16ofJm5I
+IKSMA2xp5aCmpTNiLby45qfYYcNOmvKxnc6Je5m83Z2zBo2sg7p5TtGUtfPQ0LC
DfU+MYyjaHkj7x2tYdZnAnI4MfsFG47C9Wu25F9SJGS99t/uJCRB4pa8Yr+OVpWw
ehUIA4TQQA2WOhSx1psjgMFZh9uncxANHMdbFFj0Y78uAAs7vodZhojZLA1MokcB
/iKQ12NRzkQ5r6LjBF0YYyjlVvZePaBp9QD2i2BnkQLZzMmNz0k1weTqM2C6Egaq
W0ilVygvSs7cB6uABic1S/3aU/fT3C3gKW357l3UISzsRDWdfU497CurA4YrZfUB
Sgb7O1071rOko3QrrFiHCTuoBTEHZQmzFwndbz9pHj0NJ+5ei2XFYsm0zvEF7Hbu
tHq4uLGJ5CEGdsUIC6OP3hrGyowZGquNQiKZCwwZ9LqJ7/CnpCIJnZoNVixLoQCT
6bTNNTugzfzk20pM7+NJlHs9Jx2/XV4GK0u1jp4H4kOwVUimAzk/l6UAGZXyyXlF
KfjZGHrT8O02uFBt5PI2gFnYCLlNKdG8KtP7AftnidGZ24hoBvU+/+0EKG/kqh4g
ISjnD+iMlIr8bizPCkRqHW1pYciSyYppWYM8xUXQcDUZCnD3b9LC5B4c2Bf0NTFI
Rinn2iq70KvkE9YpTyAXYh6yryQhKrd5lOnxQElMSNfnGD42uk4JwGpZSGE9I077
uOK1pctmWpBr3ewDKTREi/ZM8l73mdi3QV3SJlx7S+CFwW4Y5+P98tGfFBxQWGY/
h/76L4EPoPRu2Wyy6J1oQfEdO3THIzuvR0QEV2Ti2/ioPGSVIFpDHabFJQkGlsih
2ecqjhA4ms0p+OYzfxiVGi+E4qBVHgtVwf436wv4nvJAhp2gmMfGVQqolDeA4P/u
U5S0n1TTBsMPdQDIoQDhH7V6ktNCJ0kiRq7w6DpxpQYofSIn9Zq/DbLQDLSfS+lv
dEJJaPFQEcqS2y6cmXQpa9b8TwDXpfkpteiMKfsS+SJtboGimp20ZIHo5hysbF2m
dPOqo5MfONPSCROOdKcW4Fof1JIcqFTu9ycxJ+KlAdgNiVv7rjOIDRplCFj+PEGc
hQ/3C6SmRUcH4+Q8oKTt/W+LxiUr73MdMd2lZxIde02b8qThB1h9Usx8ZqMYigDJ
P36FwDIpXuqg7cvuPro/t30ddW49ZSlrQOYavtUb4nWBwaRtX7hVyEZ+fa0faYUj
bu931twrd5zrGntCrHkCJhAoOWC9ag93oHJz0u7/wzimGHHeuDfuTcpsZXBUW29T
blh3pNyuK1Cd3hXRXkWrNfGjGK6xqsnvSzdGVLQLSvs3AXjrgqq3oc9FJsou2G0H
pSglYtm/R8E3/x79I+oKWDGlFpid2JmaVBinE2GxyxezURBvCoGeRI4/KvIuCOtO
rpKU2kdhSN5Ps6E3JRM+GmjoGQxNyoIb0AFOnsqtUJoh/f6bl0fffBJsgLx8q765
HepK85IQhKTtE+STRAnKmdzsHx3sAJ+wz1tSv1RWV8wD+QVyQi7rFXbNaBcxC+gz
Wt7wne1kt9BZUHRs0LWQD6RRnkIine21dBiMeH2qW7L6t2LdJLSRcCcIli1ZC7zO
1xLA4RoK9i5wOn0izo4K9Od9vLHt05Ym8cQTZu0DNekP8vnanTUhsGDybPtENmLS
IV5gTjitbn2UywTQV0LFKPIhTcpcnbe+QoqptVq04HEfDeSbTTZESNX7SN8VtAwP
CZSYuLh8S+JcE/HrOrT1/006aRDtzX4j7iPVEiz4vLpPEC+EVdtgU8Vp3CQLRd33
RswCim9dmzXliKzRz9yTfAqWDrtipVhBALTMzcPXpYX3H9ueoe56tmpwabbT6A2N
1dBLp9im5G7Xe9Ff9LJ8U5w2l2NAwT4a99jJmTm+Rf+OIuXetH0dV9P8Qkyg0/u/
b/Xnx9jERvI36kHOiIKjd0nW4ILYkknknM82QqsOskObziZsL/h1kuz9X+F/USED
TPBDCE/9YheYSVuaD1dlzBsR2Hpu2Mj0+jmfF//uweTfjGg4XRO1JbaGJ4FwMOj8
rne9RZp+S9pdLlAtjZyxJHh7Ks8KsCutJfYCMJ9Bwc1LkRbUSl8rWQ9sBuVaWqQt
AbSw7vBwkxSfHeSxEOU6I12DY+LrdyqfMmVR8wrCySSy11fBYrUjOM19Y3fVuWlK
jxR5qN9svUjNTjlTtu67De8z+o0d+qsZL4RSrBAzJkI48L2xahDcQZXdCNc9gXdk
dn/ZrtGHotc+0+Vwc9+dj77WWRG7zp/b2DyfoGIycxojHq/cv2QEJfJj9IYEi4JX
f9aX5r9cTBQui1o5y0TQscSEaKoZ0wNR8I/hLEfP9ZnSFIAwrqiGRo6R57Nejup8
gcJR+Ttq9nsTUY7C+atuBEQShyPqP8aMNjDoh6W+92orG9RvTPhHyfAtCovUUHzI
cEZAZ4Hxee36eeL6Gt40iELW1c2dpT3EuyDlqXMcz3KV0tImN6GIcxILjneRgc1e
X0kJ53wtNp08Wb9+oqtx2A+rzdjWEHXc05iaVbX49FaFdZO2M+pPTbl46upKyopF
SM0xSOYvtywWXLGsJ2Og6wUGvtFqhYKTk/eGOI7rden9hkBPmond+LRubFi7pLKA
OcaUfxjg2BDO2UcbCOEfVB7CfYVPqbTEabaYLDv/1Lf9oFRuvOI4HwSYe0sYTCcv
kOcdmurZDZfLW0gwP3QDV/VKV98MpheJm0HHKHY+A5X9x2w/Bq3Zg48nd5vli2pq
hQwFzrp3eJ79vYn478NudzMVk/fQMGmdePsmFHmJsSX1jU6yqlBo9Up0H6QEcaW+
TjJjGlRZviZ9oaHSihGkGbZV/sUlaIjvZa/ez0nzoCg6YQDYf5mYxDXPqcvkk+Mm
1V0F2OPvMOxkVpn2oQqr3KZmS8Fx0OCA6CX2UjNk3cOJQV0cY7+nD+yEUGqOgLbd
IbDmjum0cOXMrFR4fQE0MzsmNvRCiQgg57VbtC2MaOnZ3CGMUtSdV1iCffbIofsn
WvCI4U2dMh5Qe95rWkc9XPeGn8r9aZabyPE4OFu5smUqb03IN8snWVAPOy+4diw/
0rN+nqE0TJwkgveGj4A+Y9ZeFP6TOfWnWTdthMYzFXAe9CGv3Hfu4E1g48/ImOcL
wJSm+zV7AACwoRBWWDrPjmEl3NQi8UfIMHO8rJDyPB3FQve50gfPsqOrbwjCHFO5
YiK3S5+uRvDRFtWSwQtAqbvHGQCJGhOc3ieMb2yd03P/3Iusy8y939H5sjMx17SW
e+HP7DpCLQzv6ccCBrQh3hE1v8rQZkhrfDgepJo7vIJTUohytVKefI//I4kmG905
hS3yPjudj6z8jrUjqGdSSyoub4vLYp3MuXfmVpMs+TXTV+IsH614EmWt1U5jqqTz
JEDqhwO8CQUlk8DYEnPrBUnsfoj7dHaOt9T/N8X9TM0xmhatHVAv9ong/SppuiLz
NtDcVm4OlOc5LcA44h+K5+MnRlTVkeusKoZlafTiJje2l4QKb4rHVDvV0+Ar4ZtR
nkNytWdzGyEK2ud8sntul15MSfKJG8SlgYoOP+uN/lh5tZDj6qHyvTB7RzlOCTW3
zX478DHv3cqtnObCa4jaR36rUt6grhEsdrnYmpN39DsWp5J85UAvQoV42ft+vEdV
fnVx4Entbd1Kabp/LflLljy6+sB3r5vP9OGQjhLg9Jz2y0UXYxm7PsbwOBh5487K
8oM0CDVoVuZpzE3Wn6vthk/b4wWrDlTTYboYQ4sEJ2Fx1iosEnXNgOPOsZT3ll/3
goVu0KpLxdfIyEWw7ZguMTPYqRwkKnltpvF0TdPiK4vO+nAf4yx9l7CObkFZ5GU8
JgCp/hh31bSxV50rBFfhuLjqwVMlQx+2XpLMpupjNSBTx9CxYHhjyLrv+MYgbDrQ
hrhfYhf7DyOwt9fz6a1A/ZeLcoihR7poo/P4AiLKSdMZIzGvQUUk4RErpPvkdX0v
Cg6R9re28vB2462cGJywmfTTjWZ4yg+u+Y21YYVl/a5bFp3ti0R/k/ja+41IOXLt
a3+zRV6iRdOUbFvovciIzqcijMReGHxfi+mpn4H6DH2Vl1t9Tc2Y8gfIInEWbYeu
39FRGU3Moj2B4Qe7xDSjuSSNjoAi/Lx05/xa0z8rT2dpiQfiuGDNep3yW7IzNuTB
NufnZVCHrsh3wDsGjAt9XSvSjANatOlArprnXpY4obYVPlgt+sicRaZFHSo91OhZ
TZ50kneCdZpnHy8g4t+AvjZr2ZHdiBPLe6oL5P/BVw4LhsJbP7/K0Fg9eHaiUavT
mUvod+YqgDe2hsWvyZPEtgp1OPrCGjklaBoh5M21nO+nZSZx2CHEyKIFCrqgX+53
A/VNh6jHVItTKWH2zB/CwcFeYCBJQpPdRAQsiTV7Dd9fl0ThF/hOxV3VVhNai02P
Zs3hg3zunFTtasm39YBtq8Cx3ZYpmALRRtAj803ctcWrVeMor1mepddKWGzmDPMn
1S91cpR/GaUGeh7gND9hs1sCEokRGyxsbq4T5pn64zOjvzIfu7HqHLkwA2wOv5/P
EZQWsXX6t8AnX6zblfReaxKa/ewORb12Q1D+YOHzQ8Mzkvj2fW4mDNYdB+avZFJt
6CTdLwb9H8xyRs4m833s2F/x4rvoWMuBVUUQHA/Ev8j4K5V7npF0CTt+pHm47cz5
sXiUS9CfJjU/LvGLJQPNFtkViiAzoryjo6lpbNZTPutTUxL7W6YlvoeDPI/tAIOp
LoGRDjNJerWm+Wp8DrsYlKEsicPAcjG2DnLVviUG0ohuZI8e4WI1uPw/jtg2iio2
D2EuhS6H9b0l2q27q8nTX2LMJAG0D+1NtTDViDpF1iCZD2jKahLbYm/IuT2u5nFW
VuwtGWzyM93n3oNZA8zRJzkKyNkAuvqDmIGmFTvjT33nLOsDJ/6F30L4PL/R56qk
veZHiITeIQjMktNX2XWfQzudbY3x3muXlr5qB1MMDJ+zckSRsTB660a9PAmxqYyE
+GcuR3xcmLp9CphPsL+7CZ46iDo7yyVY3GjyDZMotcJJ8g6snB0OSQhW4NXLP96q
3mnJkQTVF3DH1730wa9AQyZ9Nrx2yIaUqWXRmtbi/RHq4N1Hnn+nNwvHJQc5AeJQ
NVgWPouhUnKOxBF2JDnaN49CWxEchtbCe1AARAdOpPyqD7cqBkVQ1JZtMzLddHgt
jIqkgWwz4QspfuvstGNohMUtzhsgDGRJp7UGfs4+LnlIwvFvqt5pJRazMiKXRzlO
UCMiavTfsWzgPAQ/MhWeoY98RGczQrJ+L3saAKupXwIcSqho/umB2WjlvfKI250V
xbGFtgE6S1DMJEP9V+jKDMVRiQ0Lvj8+RcWSNpEqRvIJicDIrNTSQloY5GHwKjBe
UPK3Weye/tJWSHPmAMrT3yb3FfLXfcJGJKR/5KtWUJ1wnIoy0glayG8gXP0kXMup
zF2nbxzdo92pBYbThoLiytZAaJls/DErcejAncrp2PF3e/QncnEqFyhnjxxJE2GF
iwdrMwWTXQmP3+xkEhVp5Fs0ODl6SxjKY9HNEbAfD9nX1+6ppudnA+wU+SZRuWRx
qIDg3fcgx9uCJXjyAwOcUsn4Zs+R/lA3ZbuwbcVBKoPWz4mjbIBmNorthAaz0ExQ
6787S3c2+vi1Fua7V4ln9k51h/vsIEFYjG0ja4MGrO2KrcuihF2y3Dlqwtjbdln3
1B6cSiF7EFf5NN9pKhlNX1ldT2z6ij/0xHzaY5DzaG2xuRaZrRHzdmq0cw6Jl4Sk
sjv2nj9s0clXkxesV54a+6J+5VCPkcy16U6zk5q8dszDP3CmEeWaHz8HP9uOaZdC
HmRUeenLanZjQF3hO5mWGwSu8jjgjW3s4iTAdowITDTBPU0SelHmuAhEXGnWadT0
WwgRdieO8IwhvA35FC9aePGgCgTx7fCX6GNYC3mzxfAOcx/ubrwFJkfx+6XymtO0
bQnPh5jA5g1SIWI/mL9dNvlBT8xDTbgYe5mno9nwSue/EQKDL6OoXjP1ITgyjpZV
CSHKOXtrQw6wCATCbeYiBZK8Aq1pFGBARkU11hk84UPFC1yiwI4RwK9CFM4UhtQH
juCRiOZvfY5uLNIejggtuvf1iuDNy3mKoP0CNOqGLX4bom9T3W3wXdfTAH7F8BP3
0IDhlDXHtiZMKOwMB9TWZyEcYs9IKhssYh5mOfV6RpafznKys5lHeRUnH+2c3cmY
lnOGbtLoKHKgIP2cstoqZ644FalHEmFoXzxAx9rb8y4J/PeEjv9/pK90DACbyiRM
f7pUQ/3Vu9hNmNYtNeYJQcORK/lC+CsbNaKxSoMl6MsB7VgeL+MGVmuk+UQ4SGaG
HcJJ997izyQ7zoBwPsTH7s/CTVBi2OFFJrQ2J5BfoVd6pgXFXBR9HTiSCiyDe5Vc
0cm+ZzAx6I1++pyeW7fRdiZPf8QWFmUaezwdhMUY8g0yVLSsUgBQOLiuj8bPD0f9
XDWaJob7TLPEXapMKyYlCrr9SzMTa2iTobg4Guq2x9JPG8D0vBKIk1C9Hv7BGUSF
/c3m8uf2shMDV6HFDqn3iQGMy+gt6jEXyUqDTtbD4yq5b+24py0fp/uRqRRdcXph
Qd7an3tmxoJupFcex/FTGAgZzB/YB+qC0h5O9o21RaNPScUBO6ym0Z/0qYLEvBWP
UyLsTip9aNuxZbe+TpR/Qm/OlhDBNEbWuGYQUziBWDDI+klAGlE3g2Qbw0Lo9ebY
eWKWFs5twIdWrUP/e/61/RO0s2m2Tzz5yVhLtdKOCXF0B0zeILNYOSZE5LbeqvIL
CFLiCXGEWdyWWVweGQhcq2sKDtgjHkz8uMAjG7Tt6fSUgF3e1WCKkmJeM7fxoCtQ
XlI6E63l+larZmAl+5xEjLbp4foaJiPxgsTypMg3eEy9XJYgTqI008pkT9kxOrTs
TtkZJzOpIbJ4pmIGzjDuOt3HlxGeHboGOVQLf/B9L1ggPuD4dLjImq/AE8sZyzt8
TMxYVhIL+GIM37uv3533NHXwhD5cBkp4Pfq05y0SjDVLS2EG+JZoivef/xhuJWhs
gj/s3/trJF2bcRYYNofU467+ou0VWGbzI1PhefxrmwjVZhkstYhdD6L7NLXnWrPV
ZXNIoi2kuUzV/1Fah6ZSvY43AIE8n9TULIs8Be8srrgK/+Uy2zxBRk/MCZBjij1V
TArxOsnkK52NGyxoYcDyBhNEndb6wWoyCQPgmBj+jllp6hqMzMWYeSqwtnNQvidT
ydLPn/UhdVwAEUw8F530DiazfmTyrkqHP4vSfFsEpnXdkOpYhLWKqLMOg+zzxrKj
N/l3myGeYAn391w7KCU+7CgqUNJgPexHiYkdvIwSqxzHqH7V3KYZ2DReony2PbIh
dxK9KretSBJd2nSN3xw2fu/e39HmXjw+jJWYIN3yspisZ4DiAOjeeHkcw+XjZ4ck
pBcMMXzHHxJJDFnQd0OqYe1t2yLT5FydJuDPhdLYPkeyo3PjUdz3ROAcTkxRssQh
/HSqJUQcm4Afj6ymrs1ijgHDcf8JqzmN9BIWyTrrx49HbdSnA3pb4cpRari1cbqF
qyZ7lR7LbWiplbUsMAu2sQcAvyCM1sSrO6mMJCGIfwZ9vfMX1Y3ApkRbZofAIESY
GQYZFu/eIImcKp8F1GSIcMBesTTWHCk7/TONcXAglYyeNub2AWVaBfSaNJqH+ROk
8hX87EW/pJC9HUus3HCat3+pWPpZFIpI//hRwlaAzL6wXxNmZkjcp+FBu/SOVpFh
DIo8ncDM6TaiAHqp0YOOSrkuBBVXswHBsu1jdFxCD10S0ab7tgPVUrzxCADLv5HJ
8FzKiQiGpvtWIEnmAcukWPHoTdjtDcjiBxJNjP2fZX4ZzuXU+wfmuI82Q3LyM5HT
ZCPWnfJFPemf0OhiSvEl7iBFzChBGVvYNFfchX4yJNvHwicDFbIbLuqg/kiIUFOC
nrLpERnth2cdJfj778lYrtzFwx7p/3k9f+xShWRfRqFJdiV0AsF9K2eoALs4wCxN
sLhcL6PSbydkV7DnrlCoZ2b6PSa8S/Y8NlRBxBAG4w9DkH5gdPT3p6krx47o/3iQ
fCtYRoAKIrsMrxnJAVyd5tt1tudiYzxLf839B8teXMpeMrM+80egZjXMMwidDPPX
/s/pJrM0BzQLGlVqDBYePRIBgCZZJeWo+mRzBflogsqD1ejvuKsp51z8LguuWlKe
9+GSslgep6sM/JI6CN9HtJ8oqo6nd3jeQqcwpGArCjBMuRvgRVDSuPrIehDSBErz
vXiqlrSn030pQXHECWQkGFXdw47/x8jhXeFEy/l25JvPYb+hHFZ9kQJQeYN9CCGt
5gZbkv4r36E1Ig7k9QexBNGaZ9AmYd16YENm6Jh9TP99hGRgiTFlExB55zcAM3IK
FqOPn50IsLXgZ1KLP58T3bOMbUckREfwxsNYUR+wyAqbVH/oAVMunlrV1JS6s4mb
F2fTWyLcgrg1G7lBR1c4rMV3aIiML8u7gzaYaAgKpuWCw2hNWFGtM25gpCEobruP
foNLQoJSPU94WK6lTVMPIgh9x34pX02KApioTEZajblzoqRgfqeE88GbU1moK9aB
DGi2b8I3sm2gMgeIrG95OMFns16+zYtx/ISEwsvWjCgG+5M6U1AnkZCLXE7oo1F4
NikY0p2vrY40bJwGb8eAFRfdg8KnkwF2IIRTI/aaKFyRnoaCmcLtoXEQUFlwBG0m
02gaIkku6GjnOnZC/vfsGEyg4x/XuQmbk+l5MQTRSm4DIghfe9j0JGeyhuQ5HYR2
yN2ocwAm5PPTEpKX4tprdJp7LHgcALl/huR8NOupFXf76vn9cc+wvS/HDh5s2HQI
7mycPhXWP/q4in/nZl2DXVEOaBIZcyJunct1epN3Jc49U81+n2Ry3EJFbfHVRLtC
wMJlGabh1ZZwFXcJupbFDJcYo1PBs7+5lj3lMm8AeKhKxy95k3+NcCVq9Zh7Kwwr
0ZZVKVJaryOPruBl/zDY7UOFVTDjC9E3ia5PpgcIp9utwnX1NBIvNfvbt1y4JU/E
PLJG/9uIat2nJ59DTf2l5eKVcoZJlOC8PHYGaaMwpHoKToavdn9TEa+YqnharyNR
0+jZ9eEXa4651RE0u7dMDbuZ9xTn238zOPu7aWbTPx9ARidDglhHWphfxveopjpt
+fQbQWqzyvDt4AepArLOGLokhDw48QwdwbxLx9EFx+MaKhZl7BZk0befsmLqywir
GrB4tTkkssJZmSCYGJ9ncwLAt7KNKywcfd/6J332VlWvdY2j7QvAPFHVtx1UmBEb
Vc+heMQVmQki800CICqRTfFcAj6GiJuW5WTczj3lMWzucloInUL7SE+MmVkWUXVq
De5nut6bRhc3PqSsPDrJP44tUVSSQt0oAwl+t/XBy7reuNiUOtDyWNaMij4czNJp
KAi6sZH0SKt3GYvYjHl68oMJSNSEgmIilJx3eV3Ozlku3jaRq+yduc4U5zfiu4Wz
6A9azvO9ZzLLjufMK/rhICESfl9Z7iAXA257TAn2XBxYjFB7+efWAdzsEtlwYQYF
3jP633PKJcz/JIx+IX118Vigb7Mj1rJKjeui+r+RZV3WN0936ulo+5IWCuyLoXkS
XagO4KH+JmV1EyobbPSB0rPpigNHyKZt+zhzrlRQy0kJ+u4LLaP9ID5nY9SdNuTa
EkeA1v1yRT6KlVaFmFiuptW6ZBm++WsEKYEQtbEsq0NDT0RJRVZeEAq4FkXIWJ9Q
zPqZdqfL8ZBmceRW34DodVeBWUOkGyt2FKJAoO78AQbCzp9f5PouJme9fitSwx8+
LM0ihF/+iP2Vz8h4y7vyOLcCTpk0FYvw2XMQqNwBJ0VrQ52FPLVnqmBigNx+I/AR
yccC79sPRDXr1fPRsLwpxGdWeqx3/tSwCzzgnSoByKXyPnWsiRafNp5hcCuSyqtn
K1GDT4XsJ8bsTOjI6oTIVBCfKTclaq7R1yUDSerABaBZf1olg5R0iOlGqaeo4jqV
211/qqA3yHHOuqEoBk0R3845/Jgqzsrd+f4C991wc1nCAgKHTCiWhGeHNHqVmxv6
vxKtPq8pasuymvAisKS/618u2bB4q/25ZrkmFPy8ZH8jH3IMoSznyhWrEeH204Wy
+nxe+voxAYlVWKlFAcUK0wWnDBniGb2cAVE+cKWeOwjijpTqRwIopTvpBWnqwkd/
rAJejx/JAJNvApGDDwW0q/53FcIgT2aQUz+Mjyr1uZmp+WSSiEZDE79CdiH/K716
NnyrftmBzo5aE3czmFqE+MLqsBOqqqLnXvh2ykbfM+86KdBP0kNDbRjxIiWtpOdu
BlFhKgp3LFhwzBkyTGQ0SvmusuCGUhBKdTSsRpsp1n/q0lnfYOkgsePhpu0drmWY
N2kfoE9Hhty/TBzw9UM1FfE1lecj0sm/+YZRADjvRrW/ZgK4Pqv8s1+galDv5/EZ
2KKu+nWR8zABD5mEd7x9fpbHe6WuhAevaDC6Yuz0BFbyIMrIfjdP3W+SzwSQMOKV
BoeHpJzOO7BGUh2+PAF37bj5ig+5YGdAEW05xsVhk53zssRNtTlTFdDhBJGjiyIn
CcBR6hp1xkOgO3nlDUXVGiqktvMfGpNhfdgx4kGTyH1l9B9a8yWF/Y5JUBBgaRcQ
uK4mvP61bn4n6qH0A3JE7DAWFqiQJOuANIsCBYAL4j4+xK80stjl/GEhLv3MJbTK
5UPq91GRjPClTE1ke89bKltgzUL09VGajlwlxL2EDOOh6B18EzhKH8K1LUbl4DQg
tvnzvJYfoaE0pAxgu+5SNT4zL6yujI4z9j4x7jd+b3yaCXd3P3+OJehvviUe26DF
kQlnPzsgKySWd0eS4OuwdNP+yzDmqn67RahodDnqkMEpACunF4t6m5L8raxWnYOa
t+rUcxpkjrF31vvgQ7U2eb0NTwIcGNYYbWM9355bvmAHJM5QJPiEUOQau1/mya6X
gqQ9s+AY7MTbtbVS5EIrnpmKS6fSGUDy7gNMPlwYEuU21JMowZHUXlDvrpcVjmNp
554v8F7b6+8geiE/LZIcEFG+uduVcPEf6AcLZ4ILsmvZuW/UUggKFrgTNHsmVGY0
PjWcQMR2V7VTBPc1a0fopxJMyxv6NdHzRzn/JiNjwCYi6ywJ7bpePMnxokX1nYWm
eyJ1pPw5BfYvOTR/mXCILnvsAS2iNK3kTWkW7IbXrGAHD/IQOVM/m1glCdw5JZGJ
u4e8HQ96AMTgvQiisS8y4ly4E3gEifGXcdtkvBSWuOc0lKsiOIsu+HIwmwET7J9f
c2lK992UywME7jy3NiiGymeZjCcQlyAoqyy7/ExIrlM0A31fPa+K2lvPAyi+kCJG
SvQN9/aeo/eGNvSwwcxeMDO0K3tzF4KNoiM38llpRD98OFjqr9/YGHnDkbVpPm7O
jCf9m5NRABJscDtqGi68PlT/+TfFuSJ/VFlABCcehPIEbSzPa5/WhwfNtnmw7DHm
/H1Xcbl6F4oDwyuMOi/gXNu0sJl1ULXrMXM0oaehMgmxZGIM0u5q2n+y+JqyjNxH
/joWWcz+8EAPqGo8699w+5fiK6Vwj8XUuC4G5vzZzdAe3p75h6/oo3HOxGHKkchz
N/IsMKthDbdz6Px4yfXlfJdaZ5Hk1NAeQLZjG0kx/rXjXrzvHIOLZEvI2xohek52
znan+LByPsaBOJhHVCdylBL84RzELyNYy3tNkmgPR0ne8vU16gJnRQmsC0QWu0n5
Qt3T3a+QA2VMz10pPJB7S1M4fWvkxVnI2BD8MX5UgVOUOwCS6nRIsa7nr1kz5SZJ
5VYOctcZxpsCGDY6j1XnAUAGLV0nJqZwoirXR6DS0eYuw+yFKuJXw49okMxrh3Cn
hrt+C/9wA0hROWf4edCa6dg7J3/A8uI1DV0nZvrryfutXrhWHIM3m+biE4gk6hPp
Pmmq8o0rJoEbVaejbcVXJCC66br65wCrGAyI/XnGUcAkUl4FOLWL+4L+ByemggQ0
XMvxMNZPsSFMoj53YIzYwU6tZ/jet2bMvd/Jzjd9ZTVDRi2hFKPSavpvLaTFdCn/
iySH/ltVmkbihjXo5ZSnWSoM3hsi10fmPGnTDLWfU5TuU7V39MyTgUaxOTZAc7ji
rcyDMIjLkHVYvRGy7I7h8TLwGCxAtOQKBw8gIpC+nTdEK8LTlDt9qm9FqLLyt8fN
uE7RrL1GMQa9lqqboDQ++SfinoK/L01ZdrlVP7J4bdb+8ir58doqLrHDmXPapzSk
O1YgjEjDHzKb49TqSJ1hZ7E5TQLDB8YLz+VQr8JZe4YLzEXcbXUKpBvp/1fVoNFV
H4Kvayntd02xrbJX5igwnCOVS/LssWi6T3CWPteU+4VE+WZHkNltQLAS30yC0gVZ
Y0d0CIXxh0w7di+PKmajOUPcp33rtJG06a+j4nrz59xYTn3obukWdFGvD4EinFZW
5mGV9MSaFpn1C4TRrRtNnUZy+eJZQ8omoPcKavmKk4XYzHouys9eUHDj07yHZf6M
RfkAwRFqA3iy4v3Y7GO0f8R08tiReWflrnZB0Q8wKOtJj0On7KgI6r1rNkE9vCWw
dvZyGB5JcLs0RUUx15Hj6GnHioliE2YvpAUTWHxOyyYCnFktooaFiZrd6GAPyOmZ
NbCLxY+k2wZhqTuPRyb25KGiVb6gk31pVnuvDfO86UrWfBLJCk1UzpJCsp+yg0T+
UqzVNtVnwYj4/QUtzUWq4rKF6qoNePLxOV2O/oLS6KoISQ6RVNpRK06lutm6VjXT
aJkOQBMN2yyjpznNqJsaDrYYg+4hBJOEy1go+/OE8m2JbmmNHZkwt3T5FeyGpcS1
brA8a1tkby2OJl6LOQqEm26yBV0KggJSGIzq/7TVWhwysmFFZ3lLaAwO4+fkdbZg
hr0+j8HrPyYN6Pv1WmwjJ5VVaXTn8g56ylzdR1OoOMmCqhCuA8Fwltcb8Vs55L33
ZdYFT84PXlxWUpxMXxR9bcleioq+5q96hWhprNf1J/jaxiwlvKMsZnWuFx7DD8l0
vuN5qKc2cPztL9KLckKsgSYH/IZTnPMQ6CtedilX1Di8GDFH5c9Lu/O23ze01g37
ot3fNo9a07Rby4VYJfbOTuqWfLBYdKpUNtHuMlxoV0dj+WW+bI6qm8bb2sXyimL4
iLpGoz4x8UmMKeC6ot+OKwmcYDMy1uU0CjFL973qYArOKF0zBOGDX9xyxaFETWg/
e1hhzSdn76QAMVYtZRRUBxgFkam8IDoQKbOqTF86r79YZCAqSc6ZKYGwuVp+freX
ImchTWFGBa5snyvDEmHEAS5Z2cUwY6jOXDsw8HKGSdgW4c6ruf4NlrIs1nGUg4x+
EmeTl3Q1gLCmuE5dztKG69mBOEqiZOGhd2VqKb4eafHYEsb4pIcEN6/t2U185wtR
Xqcc2GIZfr/U8rhML4i7j2QaWIfYVZUKBDXubMOrpP4yP7lDuvuCa09OrPy0WmFW
IuYY2T5n4PazEZ0Hdq0RqYrMtQObyYDWCFDeDyZ1zdVGrK6nwRek9VjwASa3oIjp
fP251/g3avKaWYEBgoHR+Nx5vOV6ZJYYdVNSxZ4w37ogD807yO6GciL+N30ioiY+
N1bMAbV8lVS5IJaCcKAFhwQA+Gxa3Qc/Gq+PjKnn4FJE5nAtc+N73LMUH5xlbkCE
kI9nR3K/sMIh6S2V+n6SnVgUt2bCxOFFiFB2JQn1LIXUXRnHnqsu70DBTCABeX2D
YcaNbsUbD/32QNvk4uCBNyao28ttUsHYqkz/ULwhlRNPjdCBFEJ071nSjBTAYCLi
25qbZKXNhkrBMfUfjwu9xiJmuWo6syqmkxkU2aNDIFdKU3fwI5Lmbq3dcm1z6qk8
11jwnLUpw8j7CMvxRdU2CCjo3ul4ffIZe+ojNoECA7JcKOYISQx+cx4UNEGRcOf9
+EYpGtf+ctbxKLKIJzmFA7MCL66/MBKzWC+ZGhGtRrBolK/aNrjg9hOMy3qmSAnS
pN5wByu3tuOZ15//h8gZEkSv8wE2K+cNeisw7tA5jeyW6JAsZsuZIOkI5yoiV3Bz
++M8cGZJmcIugfEdMCKZZ8DdlGP7pFDzujS+U+wQJdB2N/bPeni+bNZICluuffZ2
lJKZNWUV7n+AMhrW+5xQwlDYCuAMxtnp1nMmRQVB/qIAlNbY/XfNIeHjArT3HHcZ
KoQbEqmca0cemqfhc7i05CTNJIJLQ6RHdsmZxQUeTy0dha3LSYK930gAXplPMcpo
jIVfxvb2+ExZrzlB5G8NZw==
`protect end_protected