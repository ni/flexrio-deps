`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSRuV1hXAfiAdaOKVh1NVL5q
S+x8Ec/svb27vi6ssDf682GfstDLM6dU/QRrOzLXNd1fhscQcx9HarMRg5TWSL2P
KldDw6jyX5jU7PP+0g+A6R0frAJdtbXUL5+mVPcbqwgdpgsG/ROGVrk+1Iyq05ld
lIO3TgeqAnBeoJJqHkYb1S8ZC7gOypArKcK13pZqg28w6rVCnA6mgwp4XPYbwV6H
oeNXvAptYbcnBNhbZ3km1iE+ask2lOsaCJBBmtFYdNBEd5iSGAcOE8qVipj7cbHO
UFHIVjOgNOQGWI81eWlbjcCc/aJq76WGVvUjHZ38SObQCMCKbvIvFjbvNVyjNel9
6lJ12MKVBo2GhFl9hwMxaFkJug3en3J2JkZcR3zXPHVIAWUKpgRGTElmXpxWF2aL
gnU9XhOmd3Q0nLnxgipEFYIoCYuf03mfnUN5G0dz68wDPbOppkl9ZX/Fzl0rh4s9
4S8nHE4Aa0j3c+m+WLDwc4Yc921ykVMuVH3BczTaQhhzltKNeuqHx12qWGJ91vsC
HsyjzqR+nsrDGCcq1XcUfxsO+qG4LfXfKJtdv6YbXKFx3RU1DoZ7iZbf64K6vODX
kfp+TlG7w57x6j5FnaYbArlIJUkiBG5twV/SNLoTScV8VK91PvkrHWXyZQ8BrKhp
7DRzG093718tWXym0S9gmbg2GnOJlAH4Hgo3c3imoUgwTk+ZIHeBKbQfZdN/CTXi
xVdg6mwk/CBrEx0Y9foJmW7u/kRTuhx9Lxyuy1VcMAKX0iz+I3YTYuzkw0TurXIo
qsVANyBpBftX98np+P5VcJbT7xqd0vF+h59cV4120+djl1bMnUlb8ANgn9xMdWvv
qsohLtPaka5QLyRAfMPYkq4m13Ali6eUEb48rk3ccz67K2eCEyUHGPJWetTMKfRG
mkWC+2Zr1QZUMbkceza5287Qm2mcYcsMYS5s9/W2nYmFIbGXf4VgdVzv8YNDHDJ8
F0YLSy7/BEx8ibZ4Ibtm5lu9BZoSKhmmxHGmPdRP4IT6nFxSxQep0m9hyjYn/qBF
sU9mtfAI78m+Hc3o5xAUbu7Vuj6QL7xh4heMK0+O5faGogiz4HPNhKvaj+YWPkcy
R5TUZSqSHTYMfsQlfFsB7zJq/uUy4J4+rpnY/sXeb7taMXnUbJ0nC9t348MGQki+
nAXvfu5pwdewKbtS8bFU7L2MNtX9u6vl9xdmq3iK7hXzPW6Ak1/J2cmswGTxNBt6
Czz8k6RRSd74vAZlLikPgL/xLyQMdk4id3pnQFJ5NTG3XYi+4S2T0nGZu9GvSces
BLPkUihSqZPI3kUbf4gFpCD3VKOyegfSsMf5oyYy5nr/DR2yD/K0TsObQrwztjdM
iLy1zuc2BLJhcepmiYtC9j4uOx3a+iyBOtzRT5BYkyWNPwy34ly3+6PlOfsO4GK/
CFfvq1Tgh+XXKV2i3/oDCKiQD7C5dAn2qNiZuTbysehwAhBQjehtj74USI5ZCV/o
C59YJnNT3ioZmfKngB39UEEGg0eFlKxRh46ASZLXERvnzTi/6g0yaeEBxUmqxxhI
6UhaC2Tq4L6D6st9AVQnAS5ESytk1k0BLPFZ08wvpFLgvdBrKauu1e3bgumtRE0A
QKwvRmueoyjHpfMScQQP4uOeaiV5w5mHaZqljBPC4NIgFefeZNdRBxnoBidadFiT
ufY/CV5TLSiFZAwZcqzHk9AB6vfDvXeTGWdxMvZTKQPt+apcShKG0dfUtPhHX96b
NJanH9Sj709oonxn9j+5v8fTYzgeis7wml1tnGmTftNiXs2eaI2w+g1tSsg1Z9HW
qjJR5ECw8G/mrhwXS8NyoM3RFmKVnVyst04o5Kot6u93RNapcydU7T/6f3EVqiZB
tayh8fzxSZ5D9u+tatmZgi2X2u5Fytu4hswP18hhJboKWBOb54nWxpUQl5v9V+xN
0cSl8zYNOUl/GHym6u7ohtJvSRs4YhK0nZHtr1W/wAccThZNR9o0uRgdS3TqFNgP
BKXryHyTk5sX8DqIRQ9ENVLKiQ/QShXhEU5RV/FR64kddiVeuty82j0b/mwBBjCw
E/HbL2jnGcW+lJdCR0OL6/AdCD3F0lUF25HsZxpaNOeaQkSpq61NEfp/dO/xUN6b
sv2NMDRj76K56lURWickPjiJ9Um1oXMHOICcQaSiNxUGr+XtkcJEssO1NKPkQciD
pjJJrwnNXeeRBTAStfHi8VH0qPN7Cl6++1ijwh/DYLUaM/Zvut80qsLdwf0Quz/d
bVDZgTaXyEU+BmzI6In48I+G5vHy3n51HvjGy/h6q3eJz22z/sVyyYZUG+SXostH
vRRM+LBEgAmjScbTHXM7c0ltDcpZuE06/hnNuVHGT9C+SfjsrCY3UP9DCX3KEwMa
CtWNWDf6AcqQnYQ43apNAu9V+934JLn+uIlji6j4j8s6Js4x4n/IUxSQwJBpvpXk
ctqAKzfHihOvZ0/PQG1fobw3rD2qmKnjZHAHmS4eh1N36HR/hFLhJgfl/XQTJyaA
tpycBfYZ3QO9e7fqpzpXPCEZND1/D0seUD436oHHblk23yBIjdmMswPkRPwRlvc+
xaEDY2xsMh8cbWRvrugBM8ujwReETVg/9MCQpQVOWpPk2YvgEAPvSdkhZcWTgUhN
eJyLagWKGT9N1T/zlx6XnZxb23GbsWaj96nyeoJIVbArQzlh2rEd0Ul1BxVsajm9
OUmpadwLF6EVzx4ZDwtFOuhRl6+9HK1Np2Ty2nibA36zefspTbNnUYqm5Vl5AqPz
QT5CVkfwS2JBwIQ9TMVoW/MQWfoPL1CBiC1OGxwqyMKDTZcnp1n8W7W9hj2UKZ0d
Am9+WgiXtp4T4JjNfOWRdT3fKBbxKkJcTrfh2kZkd4uHAbtbMJwwOxUhoY90EXGG
ZgZUF6uC8TijNYANrvUnX/BwnGcbZ5uvBVDmnsTmt5RIx+2XjDaF0yc/hmbwamOt
NDMcGT2pdP7/jD58IhBasaxxMXPUFNAVGIkRzP8whVEu2JpVCHJce5rQ4VHth99T
RgrefrEaluktjNJo7Ic31SU8MqRWmoJol5as1FDUiCQFryxrajKFC6ZlOuKGM4Qn
S8xPBXfVTVzoTkpNBTqiEQx+HMf3ByxjzEVMH1+y8I18QosYBd8mip8qTPmEl0PK
/85xRPaXxl8b0O32JVZleZz7Ibr5h/Uc67dkIidtApbGLrqnXRT/JiHN2AeII0u0
yY/VKZ0UK+zVAJOUPB5V/4UOQb97Io5OAi4jS03AN51jtaso1hPedL0pj9DBeBel
ShskgI3CgzIAAWHWRlNw+kqjRdbJqryLR600z9qrj83oi3PeiDn9W0kUYy9mej7M
09idhxHNecdfdPsASSFN3U7eFnyUd9L+jfnu+N0a21b3oRBnMl6pfpS5G+KJmRVm
kw5RH5CbD2+vjErL4P1XNc+GhI5VRSvtABZhBdOjzZaylOJ5U1N3XiDio9e0jiBD
cvDpF8RJELsQoPr68FHt94jLfRRSRmbgUukp0iDASut5X3/eCLtVPy/wBjfTC9mn
w5H+C4ANYnPdspUi/OiZKAXo4jNBSz/Wh3VYdzjIoXqZ4MbPplD+pfpcGal0Wgcz
K/pfGBPE/fWwkkMXwhT7zZCpFgVUAJ6CJNkrfhLatRucbY1af7r5+O+IC7CbHRTd
F0I8ynR7BHVUAhlNLr01stet2i/H16B6LFhvSDxGnWFBrJ+D+QV2HTxKj2v2qK5B
1ilU0kYQSUVUMr8GkGv6sDMrtcmyfM4Q+hy/VPD3fjeA4xQWLA6mcZoblCcVE5dP
saC/Ehs1cIvq183WlI7QYIx0fkHk5CFCjuvo/tscCujlzA1jH4sRYMpx+momQ9Cg
MO7KBJ/IAavvog0bZqDtd2qxjpSugnItSnqSN86wfbYJ3FPk6gPjhNyZJ2e1pXwZ
DfpHTO0VM9BIAglgU7PKAFFAHurPg0//6BE/69YHpZn1gqfFaKOON0uEY1Qj4zQN
wedfypH4oGM7UOgwukKPOTAnFJ9sEiFMsawGfh+SfqtCZtI84hUbJJ+eIDNmCXzZ
+JQjFPVjQsa3wuZZrAGsxBBxb4+pM1fTcwLz4+8ThMTovO+SBF68gNHZGgsywgkx
yDHiv7rIBheqSuyb3SDbVIuHwEegRPsE+v0hRAc/1HE1OXhzgzzQqOxoA+cYmghe
9aU7D3GgoZCq1oJSqqpgGiaibTU8IzHRuzdRnAeU/n/hoWuk6bEjiUYXoA27oRmT
OweB/L40VRzm4b3LeaQv6QFKFqmLbgEe7wzjVgbjfi8dYxNkgpaJfSFn8cGCkvVS
WfMyDDmZ6Z38phdZtHqJzqBjsA8kMwfPell03YQl9xFyiQD7e0ziJ2qsDst+20lM
Bo4ORUlw+gI+6+f+QpUPZtkzJ/a3Ax9miVCG9cCOnsFvPRSGc7u2YhzvDjqvVu7o
0uo2RV7hOoF0s8k1sRmfi6n0PvdM9J47paqW2cTT3I3hrWsImL3AButcp0O4gFlc
9X5M3zVi/Fdu2bY099bnz0eBIqmCnYo4CuK9jvS8RK/+UJYjV+cnUZrfv6LekwzI
JX73zIkiszemVyU2UpSV+HsBOu2iJNgJJ/YMcThIDfpEI/8wohqQGZ2LcbHXTyay
qvExKyV4kdFb3MIKZm3W4vxbY3RMggaPI/yHw2Ya202fd9nyLYdfW1VObJ3+k+pu
oJBsAizd1lMr5DsJnb9g8MFce7c5D5ay6iOgJvMTriULu51z8h6SQBSwOBSMr+iW
KTnLrK0Jp82aqdBRS+N85mU2RQzJ9FdAom0EUH2ErCM0JgsFEx1fi+hufTPM/VmL
pC67jYTUpa6lfhEc8E44WF5goh9xHCaoI5uVSs+PfuzEC+NpS4YuuWrJGAalEs5H
3dQ/6hOWQ58Z4AJ4Yb7N8aO16cWaEfT5yNB7pJtUjlZ9UToqfbt86fJUJZY+Nelc
crqzRrqn8GIYWhIQzuqkQULoAJ89f210CjmIlOuh903oMB0M5E18Hxlm5NcDXf/H
8V33/xiIqgx0IJUWvBOzMy/lkfNpueESLZ979bxzUjZArWwXr5U2zUp0zFdyBINZ
1GiUo700/4hlihKDCAdl+zwa2i47ejp6Y85pIV5PGOyWX9/AjTeJ0eLco5Z2hPYn
GpszJ6uJZauBZJwUBz/hAxNQfywNa88CsmMyLqDmSJciYY/VEnf5ZSl8/E7CxUS4
u7p6Y5LD4T7hVYU5fdGICi4s2MKcRgpvaT306LncMb1aVVk4O8YbUCywDz4iiGvt
dEZNmBv2aCFqDIsMj7HTDGrn1XUGKtavGlKj18rGQSyU4tuNuuhIARZeckOeLVfH
9nNhWoYbrN2D9QlaJUL2Owc+id/SaO1yhIAExXa2CTljwLxaz+klce2JvJjlnUUV
oi/oJAZYYwMVGP8uueFwJ8ZzoPuvKxmtrcp9CkZfEGLrMFd5Y0HRVYh8KsBT79+0
Jg82vd50rXaTouiNgdcxaTj7LTISUkVt9zYPpG0XvMU8NSrvvxe6LE7GLbVibBMW
9YgFUqyux3gmKSqWtaOTBNWzECPmzKoQ+zsyUo19c5tWz0xrHGvTpSj1dfNoHZSu
q/JL28CNJ+pNIQKh7Vth5ZRnDiZhhhq8kYM+XQegBulzCJtkIMiXJ+iq61lO8Iur
zheP7s4Hi8CCPJpzRBEAidbnHOUNfrODF8BOoYeWe1BRxcu0YVau2kh8GgYxSaP4
UuXAT05ChI/FGdkYkW7630C2aZFWinpIy/5gYiRT/BIsmlQwza0eNO1uoKILPRoL
2Bk/+H7NASzfL6N+wJV4QyVgrOEuDppPfF3mUwCDSrvLTCZObo2E0tbwtI+gronA
sCnpYTsrPLI3TNfO+/68kuf/g6KLHy2tClhdC8V+HO3DfCCPN8ufWRdh6d4PH33J
Ldkv5tY5imO67W1iwJpRrM3hbngyHirgKnzODlcWeofyQAYxDyB542EfOKhNZkuy
MrR8vIcSRn43V6qNMsTNrD1Q4RVQFVxqXOQlw9qgxw7oy7xhC41qNy75gXAp1LDE
XvcdmEDr/HTd0vspziVZoTE7ciADwYh8nMr9u+TMPuxnUc/Nxb6KTxyOuzaKbseP
7CiHVpcE/ranWhsGmGcAteYdkXbtUHBCONN1G46wMQLKCTl1PekJPJUd9ttvLBaQ
yXs19lzyT+VJJ7PVyUpr7Q45jNjrnV2w+iJR5j41sADcXt4DUTrx10J/z7LOV3/D
sC56DhMmtcXJ9vmcwAzVhG/+RddScGyoNsP8/9mrYaBWcmdexIJo3Hmm0W1nwe1u
qg//Bjh47cWIKLBqfnLyUN5xmplpxGS1GvDAAOeHs2hXRf5Yr7k/kJixCBCjJ4Vh
MrkB9cIQK/p28Fi4tANZ0YkIX8FUMw8FuEGkJ7nmJZgPLFIv3ZnxgMm1yCzswLyx
ve386M/G4HRHtdLLIMekUI4j90mTObdkhyrMKqA4R3aBK786aeW203ufelxZlUX5
Z9CX1REHAV0zw9Q/AKMbb7czKoFLddu/kf5B+fXpd/jh9mi6tnHfb23PNIPTAhZG
Z0SLYf/ZPM+R1/VS9Mtrl7r7wBsj7wJO2cpRzSYfr7COcqeG60xKpo/7VrTAfNEk
TEuEec2V14680hEIkUog0IrkDSz0l4e6k9W5UQj/IlF+zEdp68gGNOdJ8yGKmNwQ
kOE0RJAVp6LfKgqS2vs9wvAtKCTGT85j9fsuYEfjn5yz+3Yd/0Wzc9+Ce/Ze6Bcz
bUOQbrU5IA078ZztD7tjOFMBZjo3TlN/Sp2QMQzuMl0Aky8jbU/6c27D4bICd152
R/CZx4xPbavKz3gRGpWXQil0xOKuUv2hQpnIslggZVfT1S2eseikVgn0Pg2jpTR9
LyMWgVFlcIFJWB0BbpZ7iVHOE17J2eZ/dxi1SjOidIACV822Qa7kjBM3upXznVgw
F1SBoL1tAiMBmOfPLCSX2qvbvoGVZWl+RYSaIO0oOrnRlh0gbh1hQdF/0WPUEROZ
iDin8I57xhenuWNoY8x7qtk2asfLM41jE3UFPssqT4TH843+FoeDcOa2HcqwnQ5B
WuTvRTzGVTvjmxBom5c4MP8LU/028d5XOqngjhIS08SJxfiYuR01TmM+q/tG8jtP
AP4pjHV6c1Jqm3H0zJdckhP560PKnAe94rVuuJnAUTUDTLIi85SWXNNR5dvUmuU2
OM1nzWMvqSTHzWBkUesz/ManVspaZANnv9loAnHDu9oxsjMi8rCUtKwPtcdjGamX
0y1u21TOneL/ovA31zMpelmZD3lTOYgnlOFr1GRvaNTLmChKOalmG9keFMtTd0SZ
Zmiz/1Z76GgfGf66M6bDHviqAn7mPWKo0mIh8MkeMluKK0aQpaVydiH9l6ZE7cg/
0yR1KCer7eOFO9v/KHP28IHeg9QXl/O4ashw8pHRYWWohBEzSVWF1AH8I/z/1TVp
OGnRXJIEv5lk5vBO3fsiidl4mThDMW+/A5idRsEvKCdQKClcMAgC+/glBWQdraUX
Z9pSp2UWC+HI2wJlOAJUw5UNtJjjZ46HeZiucPzWnWPIxbNQEvdsFyaHgWUnXVER
B+32pTvVndoPVhmpmJYFBvE5RuLKbCAjZOY9koFJ6W4yac5Ifeo3PedCZ1CVlIoq
Jey7CpfyxjoqlAehmXSKNAiPki5eol/Q9oAccqfCm/qlvAEqP4YEH7r+mQDVFEhV
EAJhhb8erIF2nnKXUOIWW9Lb7zDe6P+FUDvYKsquFy3zVtGWVZzwx/j4d3zRD5OG
nGGG3atZN1RbSbWoyHdgxTdSCx4qNCik1uAJ/FGVp1x54mngK0sSI7qikzj7eTIi
0JJMblTLmVEwDladOutanO9FhTe3SKZr9DtYPR5tkI2v/p4sJLXDjOw7WBFiSdTD
Th+E9FZBEI7YSGXa4X4fG6JFXYawwlK+SrOckUbGsx+bmzj8jGRS1lzRn4/FDTdB
tEJ5vo6zMdW+f3u5RDV8t293AMBdqq4IcsWQ+uPivHDIVEqiOMGCwfwPczU+HQbQ
ZKXz7ST+DpsMDw1PetRRjy0KTvd39EQW9LggrKtG8WX/N8+pZzCT7Ohx0i7lF8Lo
zS+XCqbgEFZpFWHvIui/na2hvZrcWcPqCNA5fSwWYLB/M1mF5Yw8pdZKHNOixCTL
4+Fvus2RCM3BDBFuScv68/9MhpTXqVn2Cau59zJn9plA5QvhaZlK+FpJ1mca9GEQ
aC4yZFY5jY1dBHxpUOievAfNuBoWPO2+PXJNtDYYUpZvHSXNnpZ+kupbdoX2L1FI
8OBx0NhrXp5QA9r1cnYgNwTfM65/Z8tYUbsxqxfQx55fhOBFZL7bhzTPdfsGlekf
3zLSuOUDN0ts7+2uahpGCjCLNwFVGSpSmaH+rICTKAbFrfbrM9pcxo5c9c0Ts2oc
PiqNDfTdA6IQ/KLkA1gy1HZ1pQH86A9frOWvzQl1d1y2nYukPzmRvejiTSi+zFVd
4yy1RMeVWQBx7gWP5AouIW9JiPtyN/xMz69Kmm+aesWftq1w6JNKFiY7c7X62MdS
B0rE66EUn0JdJEb9k5mlp72OTAMqYbMVfLoal5mmsPSPdnfFirjcAsaWX2THxqW+
CVWhH54j3pslDkurHQ7hop0fGaTVKMQ3f7aTrX+ZkGr4jwctlt/A/nJKYyeovYzW
aP18YNPZAOejI70baDzfzuIF94RmYOwC36DJa8/Z+DP7udMLIjblhF518E8V7Ttw
85eZ/GCBcmPPvVNEodKylnt4TsxQxY++bJGBrPP242yRaCive4LDUI8K+bLuITLf
Uvy1lDXvkngHuiczDtER8TKYSxm1lSCVjl5YSOwntuGxfVMofYj+nZqhDNUHn7rx
+Y45IVaqgmEmZisKoEolzw5REKS0K/EQVPQJkuUuSP3ADK1RP6ew5ixSiD0QbJIG
uax0cR06m42BbeS44H/nmgeHzR61UC65CzLVCmJhUEhivtbuiM4DkTfhdvEjoRuY
aM+9ZfwuKmYXX+QduV4GkwGc0SRP0dX77p5wbjBbq5UwueZOVF0qbqB3DmOJQeIn
Jls5aSJqJsucEJPxFODKDlbaf4ZZQWPTmFe8eGrZ3QBtdnnICQFNVMHaiJLd6gym
bOLwK8e/bsL7rbJqnJ6XVQVVsoafKsDRwPfFBJBwApGcphvy+YWD1RWceKTUeY9c
XmjhRHmiqQ034Xl5Wq2lzkl8yyHu3SUmsfKZiBBpiL3J0BH3johj53aGrOSXEUkV
xVgP/uwaKylTlmN2p9AYpFTpshl6onIlKd9zHYG/sUa27aeidfREQ+phmEfJnXk/
elNx76mj/570XC7Ki07rWMZOFr4lJyX9lQn868QAx7YRpNeyKN5enCWzUEhv7RzS
`protect end_protected