`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvLeHJZWLoBW/PL2KDatzW9RzdkEiM1L4HzMrs1+vBftl
8bu5LHI79nVN0RuUID4ScIdD3/SGDP8JIzazL1xdR7sMSwMW70ihUPaH2u+3x8ct
nom9lGRe7MKzZppXRtpMcQu4upv66j5XIzt3O7VFQYbQ3WamA9h/tY9XplqBHPwO
DF6gRM5cUC0FNSwIb1nkhTgYz4Xc2OrRNQc5dBNIdDHGrMH0EkkMLWWxlM7/2+Fn
Yi+WLCUvestDQPWjSFdClc5ih9AS/3+BWzHHXWeeWCzJ+9ImTA1G6aryokKp0dnW
/XrAN1EljtJXTps36SHC8SAGdXtZzS2ep7/I7JAdcrU115xUqtx9ZwbXdF+CgTZb
e2M5QDlEqCTzTh1a7F7i2lz+KjtK02vOJapOd8T7SQ89ch3Ab9GqZuJEyXK0wi80
udMde92aJaq3c1cPC6DWGieciaV+dOd5OhXDcx5a0mW8HvvE+Mk81J0ulQVsZcVN
ZIFAj34oM/mLR3U0ohEJVbYxrgm/rNGVsD1lLm7rHiOzbtg/eCQCkDqulofTPsbp
mYt0BJaJnne6am3NfkelXGm/YsPFtfkRJuSyjJwNq/13b83rth3Pao1ATl4GyDPd
oMFKVnal+xf/kKwDIwS6oTILv6pfq//AsZTeqf8wKGAC/GtRJHyHFOdcFEy+5ANU
adsPe/pJI5eoquve8hvAaGIOk4dfsd7ZwPuSHy6Qc1Kpyw/hXnjdoxScJNtJSTkz
vN4iM9P81CG7Msl66LNhi4Cv3ernyIRW31HELZMV7GO7f12SBixWo56uNHvc2+jq
O+94JcrNQn3eX6bCJUmBp6U9cfONnNNSHmUPoeCuCRGANtCLWDCViAMNuLPLZ6dG
S6gLxqWCoWgZJdlTUKzyWn0wSyzS7Ob0UhJX4WQ62jpc38SvhXiJw28K0qLkboo/
VQ4NIJhgtoky2b8stTobaz7A8GWN3lp77b5jyX4DA/5Cc5n9UuQeqgR0ncBRwCvJ
vOLCqdjbOUrGIJJzWv2izGz3bUU7NBfEXS8Jo/U3wGPPQmH5Ii6seD5eJE2ee8yz
2eVIFBfY4Z2EImbcdkNhkr/wWTI5phiD+rp09WPrhytfNZYD+RqNTh1uWMIGUWP4
bZA5ohHAZRA8E0W0TAAxaRP3F6ULY4CFWUWUCU1TFYgcfZgdBpwS6gg0i/tiHwq+
sEjA/zyl0YzZmrh1nU8u/AOqhMPGdvOf5h+S0NUmaKLT2eMumtxWSDW6SNov+4qd
JJdbrXnUmaxOX1BF9hBRx0guJD336SEt2NLtPRTmDhS8dX0nnHocvCuqT8tANsFg
x5J2yURO7vQ9ilYbiCDPNOvFihoT3EIoH4Ra22t9SP7CBY2NBNmTKW0XiHEPI0RY
gjTuevG6xauIJGFQQsm/u7gRcJLDhw6oDo4va2IB0nXQPObG3xljh8Q68nG00Rc1
/Qw11Um30t+t9wbIpJ6+ATm1UCRDjV5m1nvcSQNeFVqgOb/W54K3x2YpaOi1KAt6
4SSTigBFOZ7BUIrN1hBTt2/45+XEDt7T6SDP6Kc6ibhfMQEJG23CXlQhV2/XGWpV
9tOXRJErkOqkgYtrePzvMcU49FEHfb3tJgdMJSYKohvp2ThKRuzhbKtwvjyH4nmZ
yrFf3TjhDxU8qQ31vVl7U/0iYzBa7pBc2QrJj9jlH6VzweXxa4RA1FKaZLZuELab
vx1AEQydRKrsCYUh9VAeDROXiu1boTcUqzI4P58qLwi/h2WtXy19bH0pl0x9K75r
jv0d7i0TCr+eTCZNzgh7dr9Ji3eIHha7R6VeTUtX8CKPwXwrruBqdtC0H1xzqbXc
An45uewg24E87JSiui0N35aW9ZQmx/pd4fbTLItH9rm6t+ZiLcoOj1GlNdZpIXxh
Kc+RPegJwUWOfpNnhP+Ptx73Yg6bi6JGand9w9gSyFdlnbthBfns6fsJ2Z5uXAJG
BA2WQI6EmVm0kDbHW1VHvNgC4rY1vYPgfQ+HNFkssnHmjmgH2KOy8eWvL7iw8VcM
gUcpLyUQWO+WSAQ2PYhwpdgE6TW4UbuEdg7dcyuUeF2VmpepYMa5BqJ+aAQHYTKj
ojeRChWEk8b7PZC/yY+wIVPbWCAfZK8G3fmWm5y1HsbcC3A9YHwX2dG9Ye4CCB/z
t/Cb+jqsrXp5XM7h7LTEP6UD/XY51jjkP+hBPXuDKAC6W84ChATTpBBLV39qcN4V
X1QEbZqt8SGZTT+YpyKjHRQwJklcnEqTVvNmcKOubTWr0L6fKXGKNji3d4ruHIDL
PM4VH9UCNmjSp3a8Yf4M2wyPRS/KbDxdpTTMseIiOkce/LNrH150tVPFWTiyPjiI
vVt0m3EUHejIbUQ1sAfEpyUjYjCe4kL3ofK/vHT1348WrxLpEY33OdIZQdLHD5Lm
Wz+XQfuerW7ssHlZbBSwpiMpKQMEuT4jiZ0KfzXQnLAu8niOTVtnYhDLOoAUI8OK
RZkPx8ZbmZ0P42w04trQoqEkKpjQYvtg2bdAIhENLjUNBYVf6wbzSFgwNucApHwr
Sfp6W3DDs2R1i+sbPARLUouVs9rsNaWW5t7ZJuX4+E11I9UHIWrefwRUzYykSfAi
UpBvFqBGefYG2/HwNCc4Iw8x5mqRr5mM1N6jvUCwZLXO4Sqv58YTtYl/iMpyDlNB
MQVvK1cp5Rt5GMMnyXH+WK2i9fgjmZrCfT1R/sp8P6hwmIA6F2madsk6FMORR0AB
q5q5JgFUoxHFyILfdbiQc5VkWkVM/Cnu2oGOQkL6zGJN0LIzO4TKpAWccJyZCeOf
FeAE43hbYlLT6e0Z7tkFl3vQ0DXaElIo7U850OQ8nNISlt1RsL2p1YdysL/54aat
+pfWpneLbxnczDsYtygjOiPgYkk2IPu/CpC1hAwrov0+Gze/inSMs0SdVuxgcZTJ
Olxjm9/7jRIMVpPg2oPJ6Mp0t/qeqBkK6l1jdqEHn9AmR/w9+NaPwPREDvNiPZrI
aadHHfnWwIeq+YCJB0lqlEcFCqqdKS5yRj+CxeylBda7mr1CR17RIkRyj/enPW0p
5HPlhtzjG9M/g/AOxhoWvPaJHYAau1erzltN9yCNy3ui7OWg71xSLvgi+EuXQpqY
rSOZnlPqJHzR5SvXrITfhQK/FRn1FjRsO0Xf/gTfw+VPvMCAmHBLdJkydzpHFiqE
FzIsraxpmhvhg3tPX5p2ER57zbAKCADz8CC3UWTNtvXGXVuyCUEBW/vW16B4bd+w
/tl8U8kGp7gm1LV1Gc8iRXG1abkzO6BOvtiPwC7GLQorSIfHYYCkt+++jUPYrS2b
NRAipCpat3B194tZC/35SLCjJl3xb4f/1ARmjKgplElsJ9Svy6CTtJOwL+h/I0No
swy1jrj3hTpC1hn/1ZFcUJRs9pOKm6wqddzTT7jaFZPhtgfskciCOPk+vXtxI6Ap
+TpbvcKiDAPW28gCUpHa1CvBwZqQ5Qk0v5mIopZO7OGf8rLC4NF8jrsR+vROGCv/
xL3G0PuoaRa0aH2nmtUA9oOka/BvQ/0i+trW4LEj62QvYIiNjZwrRs46RpbinzVt
MqWzXTKcwKq8Q7yejCL2IiYhMzS9QyaeehhqU2M4WJdtD8feR7S+GCo7CtpzU2+h
5s5U/AO/zVDXF5Jfx2p2qziaMhe7yfOg9Q8yJs2elaO12ZidHKZ9WS0Zggz1GlsX
QHnHnKphyysRiUrWdV/R6PbEcS94I/AU5K6SlwzotnnCTCJTuF3pLFFInJwgrBLe
8PLfyalwtw9BMzEZpVHIP4tt+DP1hPluTo8PRP5YONyStOUb/Dr73+45FsWXuB78
/T8BGHI9QIMEsO3lJdnn2A6F6KIFTUpKgUTVYq55gvSSYSOefhbHOe337su/zwZa
XWFxh11TxFyqAvZlrNVOZ4z9amyVRoCuRZ5R2TmznpIYVmb+XJDUAM5wtxXks8TO
6Be+PKWj4b68KOw5nP/bRdfHBTtni3s0uk39QTMSqDwycclU3tGVoyXE7aFD+wbq
EfH4WDVgbG8GamU/pwFHrb9DxoFtQLMrOIgUDHI9Em/rnlJDKjHkNQlO5/FF0qTo
beSJp1CEQl1gpqSdkG6Ext3xwTPe0WrycT/AoPEcb14TztUnWyhfW38roEnaNdYn
e7fTNh6J/SjkpX8upScO58tVR+Xk0XKhq5aSuJ9f7Z2gIA4BP9tW7SutwjiyIApL
ZD50uJvtV/2DUG3W0WxzNJpIjjwGTyvsTQZzTJD6tDpX/KdJxhrciP4uAR1AZ7HS
tjgG/jPx1TlefTKEhd6bjU5RLJMIQneLInbF9z8yzAEqEu5CBGejWq2B6D0wOR9Q
R1iHKd2YTsCsj9HHQG+FwfJ7LcnVAX9CftvSiZaaezSpr1a5qR1p0Qsc/6oiTQXV
zkgBWrs66FOdkCi/XZHFulnj/EHf7/6TirEJnYLub1nFSahzSAynXIM8DwCncSTD
ZFNbztnjC6c8JKpKmP20LQvD+eNMcsfDamjEaLdkJBzS4CDpp/ydSyS2v7gr5fuv
Qb3SKcZQHd13zTvYxHKd4HikyTe7RlcIu1kUrQVWGe+/LUwsVlssMUzFk6q3Gy/B
Y7+smxiM7Qahs3WpcG2kmSUxXIizEBdBCO3NbfbUq699GozfV0ZVdzbee4nnTsiz
W3SvqNuKlpllhIeZUy1O1JPrM2JXwVnLhTosLg2QkJdk6NGugsN+1nAtpVgvtGXo
WRT3f6bX88eYK/Hs3uawpKgcz2rX30ZNbxN5ppN+5nUlhNrk2EnfcIgT1pAg9pUC
mK9HEzBudg/SctE4QsWEY5FlYTML4bgYXP9rdsvW+slQMiJJHVHmtlfK/EP7Ei4O
oEL+NOYxMyc8PwN7yNXux+nfMZOwElY32V6hEzYNRyyRWww3KGjfDbTlxPFyNVi0
x1bMgm7dmytiFNPeoaTo35HiPcrjCn3T+fMeaZomApN5w78wJBh0EWWRqhgk3ZoJ
87D8p5Oh/QLzAt2o5LWHlUmOHCIx7LBVol/Gvbici5Or6qPveBrfllyd2rl+cX4D
UDf9TwWed46Ed4dHvlFLHJUBxPBGjDxI7mKlMoEUzihfkK8m5PPkh2W87MYuYmE4
BvdxD97DvIAF0M+SluoipiGWMAsLQGuFzoImVJo3xRh9PyWbHjpAiO8n1tO7YLaU
nkuCfeT1ihbc5u53YlEzrg8HQqYgBWinuTM9pMAuwkogF7y7+DrAUp35J/YBEeIV
vKQUiLkIhnOZCRJ6ebH7wxHt3eKmRlewDkOH3B7zM+HIf4Iu0it++F3FqJMMAPr3
ZthvVgf5rwk1ptwf9oASU59nGD4YRozQbtJ+8UxKZYA8eaVvXFoluHQt2wRJ87MV
INI2cNHMiQXtY8GT/fz1LdFkusWwAKIwzJqe/6LRfXZiGKQjS2VaQTHinG68DWZ+
317UEq6xFad9yHFj6jyqdCVU19cUUZ8WxOd7SMqRAV+lHBGycIZHK4pvdU5X7ByH
tt/muUEv0QZQIoQyrS4uCTz7DWqRNlU4XaP6k8F3okinJ5QCwcWY7LBWJobUxx9j
LQFhqOCUNAvlM5OZ2Uk/yp5lN8sX+4lVzQJeRV+mE0cWsMn75OkEfO3UbHPrNdIs
OJQx/wzKdGfRKgnZRHtsu6AenfCDDcU3UOQPPXEf/s3aBYYSjlcgUkpsEu6R7i9L
Gll2PR2TtqyVsk27A0mwwR5Q3qvB41Tyn0PjLPrc0XLl4Fuaa7aaFCY+11cY1Xm4
/YOxf0UkuGREfIPGFX/HCmKIHpxk+x/yxVxt/bBFCeFv4brsNioeN6UCNJ8fakaz
+wz8+L0Lb/AVoSD1Q/+BNbY2QHqDkQ3JbvL8fcZ4CnT3o6dCFCOsSt5Cao+4n5T7
Hhzq0FOBLOIKqioyJWIq3MNRw5ld1ep2HOcKOrmVh18NEaUJcrjwhUDyI5lZ+f0W
smjz0eCtC++bMBqAoevLPJz5rOeMNsbfVoBcThmDwt6JOtFhbXpm5EH/GJPuONw0
0Mi62TTt/Pc4QhgIup1NouhXC4iOrK4BQpjZKUwwEqP23o071Yw4DUYxYHuoqn70
pq47CTMCIk1k7BVRbCYqtf3f04xbFTrs7CfbSa8ugD1CuulRXaCt7eFcttjDaJD1
jTt4wwS4wCfFWte81wQdaJe0jCAQIlEbAYXeHL5x55zsEE/NNWmudOYrkCfZ9vk6
q1cOY6bdE4K6UIEfhA+FDgm18twsqJ/B+bmzUeVtGGYC0/k0CkiMAkCzjqO9t5Yg
QQCU+XXG3LE4kwwE8sK2zWbM7iyJe1dNWDg8WsfbVcOT/n8xzfgkFPu63WIwhVZF
o85Ddnz4rIaijmU7gO6ymKlp82h/D4ENOhcVB7B2+5aouRQfuwS4JoN+hJBLzqc6
HIUEKNbrbkNNxCGB4eNxsr/Itgh4SJgNHEINQZJH5ZvBNVqW2Nl7TQC0DjrmTFSy
ibHufgGMT+DRx+1H4wqJYwA4k6VSGAoG1t7SdJsBOLgpGv//5Yk5eAa14Z+AbXqP
/uaIQbDNE7lhIOxEbHlR1oNh/3fScm5uC8D6rpDtA9Y9dRwyRNw0g47dMUnZU5nc
0QoSOp/Jd4NSxgz8VOWIkcPxbs62MAIgUJAWLhHFS1U4P8Vfom3Km3g1rZCxMFsD
Rh0Lp/denZT5kFFAlzv+Seteexx89OWUMcomdFqPCihyBC2XNH/SSXzppBwo0e7z
O8j1s2d+ABeyjmSiDvKok/8vmF+5DT2jI0FnOb3Vr1KpI8yYJFpfPFWf/HrbqHID
Vje6qDXMGVgSsThDNAFUeV0GagLfUlC4v38IPsgatOAzYMBgcpTskMDgcjmQxyl3
gBPj4rrxSjkMQVWOzySnKvdpsEoh811STuHccsSmV6taoV7FfQ7oaUQdhw2HOx1n
qhbL2UxaxOtfd9lfH6raz75XzDNxRmQpvSMMJjwHNLKfx0ez79zYgFKH9OTyLUj/
pIYEzXr6A3gHknAmkbjV/eIuykr16+7m9PIK6QfVWpacT8IZnL8eMgxHhji38ebR
LHRZB9YsgW3B05b3WsUaNxDOYYm8qTqlhY8wsml1Dgzh2idv8VzjUes/MDwk9NBM
VQ26xXVAHjD+fFbTjpJf3RF7VrVuCW1SAmu0vND8ITflkPeax1udsndJ08XEdqbi
prXd6tNVViMUuMyNxN28jNoiuE7GvECa6o4jrU4rNQdXY1zWWZURwmtyHCzVgKnW
IksuN30qJc3QYiFzwW+B7gp1LAVKzNKTTU2HdY3iAf3ZokvgOWGSTcQ93bpW7VZi
kOh5A/s331SZlwocMt0mo4Lj+4tW4pEIv3Wdo3M/7kp5ME1auvAcuDOqwEIeUhih
fLEFMSTdLippHEpVt1vYWPOINjRO5SA4wFUd4CM3/n44pPMAUxmL6BDeDiKqJyrZ
3CsvrpszY6X3T0C/UgnsbgIHRDCqYe6nbHzByuEXziYmPVwrqeGBWG5htFWsWTxD
4gmOfrdwLPfUfWuj2oMo4lvKk4NZmH1WgIjy2H0sXwnXbDS7LB3Kn0V3fqIe31Qr
aG2jVv0j3zi76yHNAYdGUR+JVPdFczKN0WdMPj3qeIH/HrJge3A49wg7k6dhPFd+
yb6MQo5xZfP2WKyt2riVnklHkc1XQ1n9wJHyUnydUkUny1gSIrrGIxwMiHyGQG2R
iR2L92i5268H67t3YFTUF33csDwOh7NGUUS5fufm7OppA8Cq8Pu5BMmcji+TEoXR
k9Mkv2ByHqVgUcWALA7w+geI8LTJg1VQQ5rQiIymSbzHiTLqyua8Fe5jrcGeyFrS
VYAXBemEY6bZDlI6YZxnVHzN1mwRgpz+oXEi9I/5gOoRrrYbh9HnxPb0p0Ia5o6e
NZ/dsFsaHygtGOqVsHmS67hbjrJcecNmAZ1ZfQ/VlaTMhbLLB8Xp8IcpJrT5ehzX
4EQA4T+KYz9QL5jDG4gbeJuH9dPaQwKqGd8Onvo4eKw9NPDX4EDHMTh9BMu5P1dJ
qXXS6hlUkZrErcOUAoq6hiE8SF7GriSWp6/56++W965L+SxXYGiM+9krVBWwNb8d
vvfjd0u0mvPiAhcHqcCSBahO1PGDAtR0TMC6UZPfkW3hmI97X7+iMCijZMmEKmCf
8bcIyqX9MWM+FuT+Q6dr9rBvYGKpaalgVQ8gZA0E7RNXPlXSh/CbPDEEHy1NOSeZ
tcMIQi3Zgn7uR5FJC7YSpIN+BaMNm6KYf3fjPxQ91JbCeNukmyCiTDMJsGcEoJj2
sCmdbTGZf/Ir4gwA1U6qZuo/Ac0a8gbKDOtdlypJQRkWaihofqq/UDDH6NLmZyCa
38Bl/lYpfDhLvI+xODDPj4Uae2MEkgR2xYhlopmjUSB3CXeDrxDob8Pmy00Sj5yy
GQ2VlEwzu3RWLIstAVtGe1nn+ni3EwJdyjae4jeC0Er2xadd6AkpXOQjEpKbG6kv
dQc6M+BQoMFIjjOBj5ses3HEvfjpa6eMadK6Y1EIMm+zFt5v71RLA/J1rc4dihnx
zaoR3d8vXbCA5sMEtAIjDkqfPWUO7WNGbzAMf2uPp+ghYuA9IfM2NAL3E1glrcBa
nVQEyzbb9N4gIViZ6pD8bDg4II+DUMY7czoMLfhQ4557tlb/Aa15mEYH1YoPEwvD
sBglynMY8yUC0eQObo/hOn7kutX9gtF/r1HnxweeIPP312NZrruO69ce+xxZugSW
kbYEGhqEFp8sJDB4uwmKuNSXkgK+9j+SS9jaaWsRHfIqsufuE8fLDjXKSOC0FYNZ
ksMGD56CvZoBFBg6DPfHDHpw7IhzY2AaOu80u822KpywaIEo7QXx7ArwQF4rq+fI
kAKew1ZTIE4rBT/KNu5uOGkCTTCyopwpHc4J/PcjFTL89NDgQA2hR67BBjQxUhQU
k/rDJVIuLwNOB1fy0yVw0fqL1s1UE5WnIHbTB50LdKQeqysvduTcL3tNfUnfSNyK
oNd301M9KWjeHnqQgK8PTNrFaps+Bxqc5V1jBd/0korRR91+0N6MTLvNYppf6VW7
IfPQiNl8jLnYfu5qWqG+kj1r3Whtop44+Uuuq48dIQtwj7gHeNC8zLve+3pNtS+Z
Yb0m4H4T8iUmuKncOBhwTNr7STKSgrmZVBYyXx3Z2whu9+LgYlrU2x9tPRwVgMJa
bXJNNqwibm8LlyEg87RYxYEKeZOfRjVYAiqKUVDGWv1SeG7e5iyV06jKiqZvZkhW
JimLrvofr0ddA7q02vy/5h2g4Cm/1kxiLXvmwafMpRvI/Zu/AXDj+peGPLRL8UVc
NPcIDLPPo7V9nCd2721E/pVWit6NLSt5gd2oO9TMFIEitbYBojfKP1JNZBC1+qqK
SwhHmCe1BCR7Xd1n1VNsp98tsnDO/nZcIKFh/BEh/ICf9/HRIamxLoEhTXv83hLw
Zv6+TMpsAP1vhcdZ1PwA2vteL52b4Rzo2vvzzGM80YxMuH2yizPX17Rnusfs2AgL
HUAm2QkDr+bgmLSzVhRwnuo3Isi2Z50/lzQvoeIU4bGoGmnwdIB2CGMd7UejAcD7
RVwbOyr8e4z9vgqodjmxrTHaBH8DBFjL0n6QrtnYUDRPpe834DgWzyjf8vYvgbVC
7IokyEK7W5k8QbtrOe7BZLBr1GjKNGI1TDmiLmkyQYeCnlpkUHLGr6N37nAJ9atP
LoxNyVkfOrWfZwoCQ+uyMXOts6n69Bvrg4tiehfwH1D+kGVMfZBxcricO45tvAdz
FbjbJPDAhMQKgIOFVa0m1Di8JhKUnf1bBXB4/wJ8BaCOFjxKZAvaCsk93S89hhkK
V6O8+Dh8rxZkBrnnr0ByRGkxv7V59KC1wIN0TGLCiEt7nxw97nfT7GHo2JWbvnmc
DjmbfS0F+9NjpivnhN8wg5MekKaBYfRjF097OgeuLppr6qC8aK5G+9c1V1v/aZAK
CSuYru2U9rZ7Mh4JVWylLVEi+T5bUYvQnKIW1g11OGSWRtVFajDX2EmUqpygf0sZ
hIemcc0bqO8Ee3Bt+IK4+ZOmCnQaQ864XhQcJzwpyTa8xmqOlq07cRbwoF62BpUf
8buQO6HJZXC3WS2sRZR+azAaxw0mWe/JOJo1MCz3d0cAFNtOL6qNQXN5vBwt4WK2
ARk6JG9cq59ZjCFZGAN8CRsPpWFf7dUJ618kKyzNn4/h4nHp9tEuvoLsyiy/+CJI
bJIdylV815GN9UBTSXHV/xarBkbJ0PPe/sgWUOyXCvK5SpNP2mdxfA+yJpCfYUoD
HpccSbJfG55hmmEAWoMAzJvPIgGkiyDambu8XRzXHROVOqT32+sF1fThHZb1rubj
PCxEDGWO8aNF0jEd/xGZq74KTzYO8O6argVOcztdhcXMk4wKawkIEGOzcimqlhrn
kL/wFRs2yf8jNOm6tFX06knzkwH+cBCB8gsLl3JtDRpBcPelvlPJ/jIwJCZXl7WE
xNsLya3na3sKVo//qXBTRm5OWMJuLA8Td5NUWT4R5lAaAoJ4+fllfEX2eFD7LxOi
BXorKzUOKF/2lJueKo/EvzHwefadPt59eNgMF6jNW+19LeSQX2hMSb6QhFULJKgD
8jb+i7kEnccnMEwEYB+wu+m+XZ0BE12Cho2IsAeJm+3VHE36v+kMEwRv9zpclJKu
lQhJVAOm7Q39gqoeaXbnrhJ/TY0Sy/poChEpvZAR3fkWYC04e242auaX4J0c2VbL
XlaLKMkxsGJ2yn1W5N1nOZOOWJ/Z+iNfNgboRdWxdpoHD5Ssx4SwhoJ5SMqL0crU
1fZBn1F1eDUlXFnyLMj1WfUTi8Kd6nt3qAYatbz/G4K8IvyClzJoJooEUkjdfT2d
xTiRB4z6SzV+/bLtYbztRo0afXnrE5n3LMXa/vQpFluR8aRNVfLXB7cTcRe0K+T7
UpX0m/NVCQChEaAlW7rHZzJBdt6zH2qERetcBAyYp0159rtA05FPpNxg+IhFf+j0
qGo3LS8pfDTRsub1YeOie3a1/olov+NMu633MUA7CQOeLhzmeXojWY5vbedjarZ3
Kl6G6Q/G2mqu75cv8bMtjuLj6ltlFJ09oUFkiQiQZtYUrOVAA6uV/iEALO+X5h+x
Aom+28Tk2HRE3Yu8DSE+wz8m8Zn+/16SIqOKPb5Hi/YCo++P5t99sl17a69rFoxl
jjy+Wml353Yi9bNNLjC/z8THDZd+NhzOkxi841Qxgs7yy8hTJzpXj24NME2G5Atq
DNYHo2YGlQMi24OAlVMNbDJwgJ7RGQDVKu0numtZ6G4/byQiqWYDmWiwnN+waKKG
yulEtyVgS1976j2CsTMjKoI8PIn3HcYse1X+KZbaD2dKePEcrPe9UNvEJLJQ8+9F
sYzQXlcN/4ID0jNwG/HsyzA29nBKbgLKYIACYrRxJIQUTuhEGo3EFaEm23TCZnuZ
a4Zqp9p4wQa1gDXlbQHV+o/+fHmjP+yM/K4w2p7ULseXPGLZ6gp5RgBph+W4pmUc
cdiRdGkJ14ElkhINew1S/cdawN4ZtvfLpmU9gKKXwvyo4y63/ICK77AkX9WEgin3
5VRQjOzfN1dpx1A0tWZ2goKbcOvV4orXuSZQTwuJSRTKJJWcmttzfw8nDyPUJVau
FI9CVEpFdrySQ4dDDhQnN5AnfonEpazHNFE268Rp51v8bcmryRGi0mHF4E1EH9Hu
0vlktFFAVQARHo+6+i4a2uYrxFMj3kCcmeG7de1qeSG9bV5f3nAtkv1FfKM58qqq
AFZv+lZ2iO6nMv+sxZOUFaClE4DP9J/OFXWRTyV0eR94NT6tALpa78UnMDdfLcHX
jad0529XHOHKBQiYdTI5GxLgfdevtxWe5h6osV2bKPHKgCzpO5GrlvA/b32nQCG0
8OFvSXRVCE1xp8bJhXCYt1QxOrmJhMJhg21In/u/8NhKMgXZK21L1NgL6camG3UH
yolzP6A2XiModkLzXnsBPXmhCGx/0laY1wt8TKLbcnvaUV9V2JRwcmSrr1UteSjG
Q8bI1I0ddVR0/laDcNpCUJbnCycpy2ha8mi200mtx0QS7fbs6kqTETiBbEiWAv8i
Z6oqArZRGfBoWn0SHdts5dzgeHCzd0Zke8Brj8Br9oZMzsGDicugbUGqE5J6bITx
gOEfxWPWxsXLGYX1jnQbyARjH96FYLjHijnzrE0cMasuuEGGoPRGD9DH3o72KL/c
CcD3TcrpbeegvhbttPPJ/V0h1WyT0A8FSGAwmir+REmX+NOsdflwH1rIqzWCzNtf
I38vsG2hm0oSxW11FskyoEriOhltkswGfUdX0K8CojR1qf67wRCXqGUovYekhpFL
eOte6NCM/ZIbWcUm/on7NbxbT9i9vaGUX3sM5gW0zAIlWcIweoA0W1eu0HtlgLR0
KsA9KIVgSHY48Ie0K7cFWH+8q49FtoomnGCNi1OvCBg5LkwtN5po8L71fk2NTS4t
JIh8qNZfLoCDKqiWUrNK5fEGfwhpuRWQFL1/cL18UZwFTHmazpuOeZRi2eACfeD1
zXPEuZBDQCdum6RnuWWGtoDKodTnGVcd3goaxAOwHZYT1z7aaFMVCguFT06/BTZw
KNu0aBmj+ZsbVNaXZghVxLbaWPChXML1bzboGXacLsvFciyPkg06PmhEq/B05ke+
Ec5OUT5BF5gWbZ7mdpGhf8Zt7gwgwCMDDbULm1nUUcZyxLd/krmIO5w2tGoQWS+l
v+dALZgxxky+ObIS3GnIqyRYTKxAa2CP67U/xGnlQMApLazy4jhBwGrJQpHvzrwm
LG3u4Gka5m6L60b2lH7HT+WiiDBPYNIOZvIU0IHW6j5S89Pg13QPZd6HbUl/VwTy
aBub04K6HVpLuZsf7SUxhwXRiADyrKRKTLctRYkvX/A4dGsnen9ZMj/H7tBByU8+
jfFXWj/Lo0zMUXJrfv6N0fi9KFrraR6kVpn5FnWyHOWkzd7tJirmEnPhCGPIwUmY
qKlVpzsq/kN6QLzWFDyss8cuSrEp2gyrCJh/rCdIOP2stKgfrpgnP9I21ifZ5vo3
O+om24Ko0Nf3Rk9lWaa9rP2SRiKBB9fBuwifpeIOJhWfah2nKCUPmJBqhlPLkCyH
+ykun8HfN1Q8jsFbfbQANDcD1HxWvN3OLHknxg5HJOlK2Shv+wNzAnG1zbsL8w8E
YEGU1Pxe1s2g2bDMa5vKOxK7MwV+2IKmqXbmBrhtaX0NINOp8osaRT5PjW92T06J
kyQAfUuYt8tBfl5oG9uwG4hyos5EYLNsGMl0du6eTwYxS5HqEf5A8OFdNXc0Tms1
rf0yzBZ4tMahN7PIQO1t8URaK9PcKGeR54zs5X7b742EXrYpz2LxaVixeK6NT1CU
fTSCuIIxAwZKdSa2FgdCSQhqO96dWzD7q22QgOZqYgvBsiK3c6AF4PTom5rET2Ko
3S/ec+bOSYXrcDXYMqfWXITo00v/ihOfTbK1RbioDvHwpMKdAG24L2VZ6+Ke/pug
kQbj+1oPZwZkJnrtmL9eCo5iLiGe0pbGhVvSFW+liBu0HC9W1f+eI46c43SccLN+
Xw0T8Hoq/emxemdlAMAhyf9UL+B7tp3yh9brmNaUWeXf+GX2AD1f2L099AbYQMz8
q77tj4Bu3ZAPrQZmZ3h5Cz8NQXPIYMjOsRi/MmA0ReM15XV+VfgSRL/Rz50SxmSj
7KZEHNgdGlUpQDdZiV4a1dMHcuOHU1x6Kzk5L+dK0geexWvShnbu+WjTvPgyieJm
RRy+AnF13iv6qr3gAE9NowO3QA9X8XENK5VeCysMgZIzHJ4zQv8EELxGyauQbaZc
/r7NRQ7kT05Q64sBEHBck3lkvMlLaIGdCddbHPDgJRc2vjwPFaIDaKTpyMZKm8kd
0NHdMkz2hraX5NJqhkOchVJYk7scOjWuR7xvs1+M5xRJdO7eWZ6p5aAZ050kKXx0
E9xA9EjZ4Fa0GLJSEF7G0FDfhRNl/jevUqCq5OkN6kWu8Do1+4WMrdGz2NZY+A1M
zezDbI9YOQ2DB21m2K3sfq49Uuqt29SY288xLnLLchscu9w8P5lfuUQ1gyaAOcN7
sa8cFyxaQQT0b8FFCakQNaRJsrpLgtsiU3k4Q3trtaWEvj38jDOgGmda4WWA2SGn
5ZSnZofwsgEGyrquXRF05OYK9mUlgPJjKyo031PT0E+DeLRSUj+BfJ7AtS2nz1Nj
5kgpn9OpLCNLETMSs/Jo8KR5WeOKwbYpzkAsXQxfNIGdjcCxmT5tXFAY+Es8ppU9
nrzvSVV52V9ysIqPt2UVl2+Ap2MAwWpNjiulfD8Q63YbZdgA3yGIgF98ReDpkx26
V/UwHLKrX/Yox7gMiVPojx4NFquT+e0d/KHfcGt6KY2glwkqVOqQKqx6SkshDH+Q
6kgRxyhmbwbvsuThUhuYT9M8lcRFP4JVLYv2wVLPYbuGgMaS9LR2NSR2RyH6DwTM
d/93Lgr/wNp2277QU7zeu9yYJltXyrcHTh+AVjwGXIt+J2P02ZRwqktDB9QEJPrW
ajqHY8S7v5Ifq1DNzXmPcqkuQqL103vw0f5ASwIsFf481alwgd1OLP7s+58/sef9
KD85bXPYFtr9obJGt+8M2XDqOmYLm/et3gopf28pK46rijlSGINDwg1//wq7Ddv7
Jg2iUS/wGU/nUF8MfRVMneiHdR7l4zBpvGLY8ew8nddO1xc9QSuntCAJX0fA48QF
4iu1jOQhxiNovkbdmSyo0kemedxjgb3HZjBSyMyAkrtwQntVWM+QJHoSFmEelNRR
ON4zuCrSpz4YSLDDMeD8iAmWap9hbE8BX+dl/+owqCDWiTpYXGr5GtGUfCoRY5zb
CQco6Mo9dcDygnDlJvBd0XdekVnt1MpqmvEv+zAelUTI4mz8hImDzCAF85j1EBHJ
f9LUZJ91j1OiMWqv/5I6zba0wDib3qucYy5bKS3Ao790q5AmWZ2w+JTEbJLgkuez
c2Tho/mcmKttS89nJHblnbagnW9WhnVoqjFQBhOyxJjZq/QcxXNl+4K14wu2/5Oy
+0ARKQqj+Amvqjqk3a0a9Qig4LR5iHo34Ys6E6vhkqyyHeLSbPTAaFShlNC9VrfW
WDglORGjplTPk7nVv/wH8tLxljBWRW+5Bhwmln0ItbJndwAirGO7KtQIPHaeMzv8
ZJ9ans9i+jLFpw2b4mw4E/vzp1YVvnLqHE7kAtKodBcmzzj3dk4j8vwQ1IYLjb+b
3t3aAHCa9uaxt/MlQm+/bKiHL3X9SCaG54g7hNXtYlxVDQKzH+aqWABqA0VmETKq
9b3G4POyF1MzhMzDg/+HlOlzNTlmTfx/jbAlkucobkjCb9UyXvt1E9TY11XiVMic
yJE14nQHKWfjpuGxEwyM2L4HbLSUb48l3fsr3vgSjGXBfkNglRQLbFfAnky8alI5
U05IAwCDl27rDie9ICXaqsniCfb8ezdaLMoMNmhFYCwMo8A1qVJMDN++8TQQ/gXE
twkK1j7opgL8/ZqH8RohjuycPUVrLwqz7FweKIq9CD9M+wSgXkbkcuVdB0QDKnbF
Um4aboujhLXWHGGDGIN536L/dBRNJxcTC5dZVVi0nZr034E9q30qTrPXtlZammeQ
VHKTqWxS57OOuRnoLIh7Nl+0JaRhW/UBmX0ztLM4+rbfTjijfJE8kTDHw+ZvH3eN
wCNY99stEfyTPDlCW7L1eidLX71+uxyB7aXk14RvVo6UKIshYWxiQtck4KWxbzVK
QOxUE6gOiS6P4OgcsuZVDR7P5dffKCQmH8o2CIjrlPr3re1IrqIt/w0Smp4P2xSQ
iE/rqo86rLKYhIkS11wiJ4TUxJlmAmgmqyJ3bV9WQT4xgYXJDjX8u4aVDddtWJQN
uEOwHBf0uI+30H0netzqpPTIlYcl/GJ+kHrLjHGTb8CvR2myzjvAO2/qrd0dylG3
dIqfgTIGZRKCErkqRlAN92QLPncs1ZyDRiBNduJBkYoCyGnn6FBojnM5ikMN48dl
ol6MeDLn1Ss8cVShlV2pHw==
`protect end_protected