<<<<<<< HEAD:flexrio_deps/PkgChinch.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
qe1+t0GXQ5YjcbQQEHGgOYi0TZd/WF19sJ1AgVIdFvfBsp+qlYlkup4zsWoPpDIX
D+k8Kbn1b2edmiP8ax5syu38mBndf5dhhPksHIJ9gYwM+O0UPzw0eC8ICjh4Maiy
y7lu9Y4dxogZxU5wlZkrOFLg52Gd6KJ6OfokEJHXWnvccPLr8UWrQb6EwWdVGl5x
zLfht7xGAiL/gm7zqxAUbn5T7tkE0kvMbq9lYCxenBcOyvuNm9lSUGDDu/W5bVNQ
y04Qb8QqiRO3KxKohdR1Q47H+1Rxua9NZRQyCGATnDoMbTR+f85uQXOX/BaDS3cz
TWtfR5OTtpT1yte+DsN0/JQI/qYrEC5/BtjCd9ZXNezseQzHLtelZ4cgSrvrU570
VCuu9mYHBIWef9khVZ3AqNyNLeqxWy8BqlNyI2bpWR5+9WeBpCIGFeR+kSwFIGNv
01CSf+/oW/uNCQKJ5SmGxwE7AR1+mdmt9fePgCO2vr609xV8iRt4oHhlES4KsKNx
tP6+nBeRHTFc4ZJuSvoQ+VlHx8UO3iUvOPvpm8EGGxMcg6DcZMpguX2HFeX45FxC
1lWLpFNXNc4jGgarY5It+htlncAWjTqCkgeylLz+J0d5leuw1QwI3Bfj7sqHHiRO
6LnQjAiA7n1EBIQeq8zsk/ZLVZwszxihSzX8XP7tfVHGWOVTe1FIuHS0Wc0obWDb
nk/oESo3XqdZCPAfEkRUgukoZmE8N48sTNlTq7vifExT6qGqRyvmy86k1F64oNtE
ELl80nUgFcekxTwLMfg5hrMbbLoO5zQztKVWDB+05DS52yQJ1EFDqshyMhuFMO/y
EAOAfmjKjd8RMnwzYwERtyuewVAlPjp0bq4WiGgKwVloQTcabbcc7CgbITvR96Ni
BPt+Y7e3XUFThmzhFsKmWx/HS0uwbdSIttLlX4rGJZpQk5LQ1I16C25Y6gSz2nKD
I5fXIgH+/CihEKVRbkwqx/0y1ABWcTgZyJ/F6yx1nR4XEo6u8fVQ8U7qdCip2XE5
3a7+qQgCA87Rfw7GjT0NS+YiqnPbe8GMmsIkOGKE6x1As6c7pB5ydQkYcLE/NTva
2ww2n1uHqzWsSSZZ7ZeXFVQwn9yn6N79Le9UVcYt9Zx/zOT4TBeI5vpiJp38G0Rw
7+z5wGcABS9OZ7PY3YUpMUhEDI1QsJPT8fLOI8D2UgLwDQTK0kh5pPnf9OULvGTT
U3UkB5F4gXpfjtBdfhomqti5MqZRnS2UTSdgYRINexSRf+RVBzh9ydQLNkM6Vj/e
oKnVuIVgVDfi5gRe9eIeZYdZMhum0iAYRlBIsvMo+61XC7tsiqfbCvzksPSb88xC
+Bvm5lwR9wQOV1Y3ydvAy2pE+XfMA5QaXY7SpJH0ZJQ2ShGNheDQb1cS7+x3Q5S4
Vqe2oVa6/KoftLSTaAPQAuSxikiaaXF5eletUIjHOjNdFAcKLlyn8Z5Jqzxc9tBJ
pGye9HxcuKF/A6eRfXDoCuzmdXlhcJVSq6NMh+nc68SwxJXTM5gyr703qsq0TMSN
8wyLsdAjCVjdh+riIDeC5Sf75BKOqZ6vNVKPJJGej453vEaQnuG2YiUiMKz6UAP5
oO3WRITfTGgpvAWtVBLJvkNnp0+JDHiGtec9KBK0QfTGw5kN7pdvS/UjP+w5rXWO
gZMK2EjijPFUT6Gs4Cc5VhC+42ecK5zcTPoTdNv+g5w9dZrPF3SA7p4G2R5rVruc
ICR9Ulb+S60CVOi4T3yhqtz/RxUnwljPhpiARpJQRSGaGM15hCsZcKkXipxVRC6Y
JuFdNoJzhUhp9QlsS/qJrJaDbawLn2l0qZEGDwQQ0GYmlrFm269gDoPl2j+0L0K7
xLvqKLrp9lbg93Bvr29RlJxNq/uskAblvee+ovDVyLmADRMMvJE05/+S3PQSKiWk
Ov/S6oiImYOAsc0p2/q+a8F0X+uC3DbfBPiv9oCYG7iPTCbLnFzu4BUpJRqSxaSD
j/Cvl08s6wG6uCEkVPpxamVHrfASGWVDGiJZPWA8DS4tk8DsVBVyfIfRJ4xdpEeE
oodvPNYXAUdhGEbDuGrdsg+Z+f+VyKLguNn7rTaPDwzu/dkwPjS6sHUYqOgsomgz
osvAPr3nos334srDhlwmV7vCicpg65/Fjw+7M/1GUKMcXji5MjULZT37/CNtYSib
xyKutQwgPXom8Fjym5ECV13mduMQVy+t/O4UiQ3M7aM4S2cnBQWxtjP2A+tZ7afO
J0DUo5WgOp2iIzIqutXfVZHanOXetWhg2H8K2XkkOa1C78HMvGX2qnk/TZoEgqGW
0Jk2gD5M5FxEQ0ynxqqWQQQcaCEsZ+wH/3AwNJOUlDH0nJ5LI2oW/zrPqFQKr33T
mnbqd1tODbk452rzs04iJ9NOZ7jflvuV3TW2272/yymgt6jKKz4fiRATAdlkJiMd
DTtN+K/cFH2CFtt8kgbsW2tg9dqiEUXrPqDPysyXL9B6ay/lO0qYJWUI0BtWaeOC
3E5rPGr6ynzSi+sx7ru7fL7eKwek/7xx40fKoq5p/2IOJgkVZNMn2z0vk2I7xMd7
+WI98L+K8wU8BY4UsLbW1+oWMB6O6LDnLMS6M6Lm6kPH8k0hxpfOUZnAj3Z/y0Ku
kZmcj5kVklEdYI89cfzjUfRSIZ3c2v1xaCbH8ValWr9cqV0Oc70B6+nto00gLJZt
23faY1aRKoafIqEjKXP5mtksmoqHNcNVB8HSdBFxNRGbdaSvtThDCAEBY9HPu3cz
sifyUMJmH9EdwOGfNuVpVGxSHKUIODMibJ6mHEiKUpVcU4bhkDvIZ7lH3j5TMTFN
bPEX+h4ayNNGVuAxhUXYPcsCW/giyFWQIo1o7rTw46NBKyBdZF0BPVk1UiVOuXP0
X0M7BOz1eFTCAgeBXRevaZP9zGwuRQfciU76nrXBFVcAHjY8g5tZGtPEL3Xiybxn
QoxD8Zq+60nXXdGlsMnsaEtcDIMvId35vou0xW4l/fIPoytRyI1XYoXGEyiwxHxS
MuDw1WfSSxrMI/g3ssBsb8g3G+s8zhOdHFGpcMUstz8dCIMi0XNt56LDbcy/LFRb
fxBb9Mjbplrnafz3l1yCL+7R6hq209zZQ0P+cIc0eGbpHiVKqKAS4+M7g5A+8MUL
g8O5gfG3o7QCTRThEX8hOLEHosySDSP2Ms8Qh1xmmMRUvsSchw85Z9UUKFge6w2J
f6qiQJYs24KUYLdwbEvtaxj5pLLQ+0eUtNs9EsMM/aXGrxX2NvQjfJSKbztgoYvf
6fjnQUC82hTQsqwKoCkbL3WvAD3c/H0/J6K/KzuM6ADKEhSrXuKAGnE+qpRkV/rH
dz0O357NvnSB0FyssCkcio8PpTHRpKaVFSb7Mmu75Dv9wnibrxybY5tkpq9qF+o7
DQphQ6IdQIoEOe1rxVW3O09ST0TWuubQ9ez3engHl56EbUxx7cf9FvkSKL6AOIRA
HEDurgJCICOe2GdJ/EdizJvIHmOf0QJvwda5I7lRKkAuP98hVqLafv6/eVRQXIyK
E8iM07jz8MTDx/xmc8r2N+z6Hfzn3jO/IBcllTjfPdpujSjJ5HrMNiMU+t3VN5P1
K8jMu8x2W4ZnTQDBnLnz/nJehn3gm4IsQPQ4881W3G/komeQRF567TIzAJ6iwUsP
rmH1yevl+TrmTiqG5nHkMA9l3pIKUknxZDufByGICW4PBL+DEFmUdquuIRxLeVXL
MirPsLWt+xHHsdrEb/ZedBf7t5sFfnReudDRN/x6d1qvaL5D75Ydc2YpcYOkeOpE
bKTC6w2trrGH7RBqMLOry6r3Po3YSMJ73/t1btV5S1xsx06wzebygXkv55+qCQhS
4NLkKa/ZUkcT7paDdISoEx7AEG5rQoz/wyvw7XbVQ5M0jSQW8O0HK3bCyT6y6dMv
eSGR+iw0xd0ziS9HoZWQdvv/4I/+Zug8Yli5qQsg435pCJSBqcdJ3uSxHy0lD9dG
xnMA+gi7mI3POt/ATKbcg8nbNdQ+sA0SIFaZ1e3iimPK6y9YmuMDdEi4YB1hvMGT
WJPgrrXzoEAkXAW2vsRgWy58Xr0h740rGtZipKCnef2OzlmxTptiB/7I8H3TV7Sf
69zyFB33Y92BYC4Auy6b6q1nQzj3oDanw2ESnQOZy1gnQs8Y/5lJIL2d8zoOsrO/
tHL7br0IYdQORB5O9w9QwGgm1zkvqHb6/ixggsX7Og9wmNNUuAoAMijRYzpLgaP9
1m0VfallKYc1GymIj38aY6bDhu8nKGJ7W98WUrxsWMVKjj1KBTXA3WgZcDtPrb07
1vjUG16TcNZE2GBWytU2nktmJjfXtgQdEXQF4FjfFtD+4+oIk4xFuF0Usb+PcKa3
hOMr70r1V0J7HTGnphiG00i7W1GtIP6JAO6u34m6KrxxoedFzAw2LD8NRGMZmgBj
rhpX1S6fsf3Ooj0VyrbaZ4OOrtc8jDPdr1kI0aoL+trTR980PUOY1mmfBuNYecgG
OlHCcK+DMh1p2GPa7/WwA/MnQcFTttsSS9PB3cQOcUcr4PMIbX76o1o/y2lnDr6m
k6SUTZgapXPzTkZyyhF4dUDiAuVF+PEUjfNxRGamunHvbl5pswTlqnjF7FTG6ElD
mLTmjZTUJOT6aBUBXqDZg9YvzOpIz8UEZRrPcmw/vcjlPnj3m9VrkR/WNuv50giu
sMYBghH/XJTo15TVCmE2usF8QdoX7mfgeJayXVcb0+Ux7W2zHpGLXxKWIWwCXLp7
nfj8aLsHDOxCwfm0hAr30FcLFexdkEP99glsSFy3Zheh9PBJv4466Tr7GOYmg4i0
OJrWNXsU5Lk72O4IvWuBTbeHoIkwpXXdFoMo8E4c9IlSsM+buidbix5DLBn2ZGMs
1scwdGPpa5zuneJOPq40vxsfENceokCq05jjAKVdWnAG5zEVbzckPn9IKAanlVqW
lq/NwV4gh6hY/cYFczkZRBQi483cDaQlK1x/6qZ19UfZqW1VOQGLYiGnl3aZ3MIb
g+hn2rl+BWkKb4QfSHrsvKpbjaXtiZ5g1rWqLnZ7qICGmD5ImjQ75WytKoIaYQ3E
3X31L9X7AFLsgkfHSIrHvNyLs/9Hh0MW/yZ4DZ+5cp68TypdJYmHgbyrExvY6kU2
zi1FdGcTxnOc66N0bHgmplJusMLnzNOF6CJSEd5list0sM5AYPn/Jgn5Xohh5WNY
R3WGVsfva3qymrchfhcpmZR7+vX8Q9hvApAe/drMEQXa24dpfFZbnCJnmny9yv1p
TVQe9K7LIQJ9x2Uk4q5kfV7nK+4j5+pQ80XUr2zzIiWHvtJjc3ea162TU5/T1Q5S
A2N9qDEMJwjRM5OzKoXGGJdH1cGIAb/7I1yycKXn8Yf39Qq0+u2EdFbBTDmKEY/S
CXz4SUXtnC7V9DbBk/5zJtGqGh7p+ciDe7vjBErXLc80+5pbtsy+me8y0HDBlYor
3dX941YSLxFnW4Q1Jo7ol/yOeaSLykr40Uz6unUZB4pkH5J+kkpCqRVthCRdyj8x
KLcDGxgAEJJmFPApi1ECylfoMumRCELkbkJbRECV/k0kxILOd0G1TZbk/iQfLXM3
bYeJYUneQVW7HKzA1OVDi0dCkD/KrARCYu5HhRWosaEdcxKNgaptcwcvdRPpS+Jf
EUFAWIUtoeQViEpoXuJR+E/HyA2jb5/U7/Nl47Jqrq9MQtmlU7PZ9hKDTR8lj6hd
6OuF2y0KahH09TneNIcXhIFqPo9wBDXNVEijaCGNelYmhED4gLoVXemjwC7XEX+k
isjBBeiVfD+2UzOMgk7QQC92vkPBWJbe0M7kBAfdoaUHnQuOcKwNL9sJ+qeON16R
Qn/cDHgoCp2soS7YoH9UfOq2gbQB2tS1BMrIDbf+3WwpWRRR9v5kA201SYqNphkM
p4g8jXvFNVd+NeaDdlg12nZjS6TjboqdRQ6luFsSYmgBnvBM9XbVoWOSOtI/JBQF
xG3Wb27wsTVzN+Ju+o8pFOYqp3UBD8yA+S7n1Ur9Z6pZDtwWv7hfNyjuN/opAHKA
L4wAUCN5d25BCDq/W65BhUpvvzLYHHkpHEr1XrNGX9mrqgbWXP02+JJSzRn3ESAz
o8Cq7d8ibuQi/7D6oiiLJZVatFGA8K/5231bPoiXSEEGnKqGm96URj3tQNYxOg7x
Etkl47qOB79+WAXUBZBOWNaC1WZBfscVoe4vlDZl59aCHkA9QojkjMcaWeS6g0le
9O6xdDwVBftV9DqdLWtbPH41adGBADWm+UuhnOTT+XISPNf7XnlWi/MmfgSQDq0p
bphP+tLL0nVB0oB5X5sp2KX24wwRXXUlU24k5Zla1jKM/N9hFqPERZQhHc+6yBI7
jdpLqCTnm9+vnLgYIwEB+KHsMYFbBI++I6SyMJSYXZ4C16dH4yzQ6f1bU+rqIDjg
0cWWETud6Rl6qkujWPqfHN6Hn4dMkTSFGxC17c50VkFQXIyZ0FhYu31T4L1xAOn4
pZzP2myFjDGrV60QkogKAbE5TTDXBdGG9xRDYDSzUiN2dT8PfZPcHLth8LDV1bqQ
WPo69maliwRfMKOC00FIPDMi1AUoOBLDmsn+6Ir4mXoNlHhmoRfF4L6ijqW4bOKf
h14R656CAyWu5sbwOe0pV0uupDaq6i/Uqed6bE6d6u9TLZjwoy3ml6V1qtZoWB+l
zFIVQwu2jtjU2IOtXPP/1fawyJ3GZTHBSLS2zPM7oYLFkkMMEOtdcAjVlvo5ykUz
wQd+v+DvMslBN7NleUl41+h8ut24QDgAp5JO4ImXtdklKgc41VMxUBXTygBIf2jV
SwaOQ53Jo5kSuna784XtYj64BeOzP8UcClLcgZoSpAOXt1jpzkqx3qWzEN3lB7R0
doKjI6xC1WLafTkRPiCsteYPm8JK0/SszlHN3hHhko7hHZRz1/l/uS84iFbwvc/e
Mq3AQX+K6G/BEl8GiIXw6ANAt7mNGdy+rnXl5hVA+0+h2aqDxwtSixTyXlIM7/0N
QPlJWSkO4ZWYXVPU6wcDnLipNh8hUxWE0lVPze4dr9GmVLN0i/ru8HiWG2pz1ruu
SQyTPskmucuki3muAz4Qx831r1LJg85RJ/UNVVuZhxHm5nMRUIVnRIcnrGt3zLzC
m/7w5MJaeUCbyPnt28BW5Y2ROge6gqu72p5cNuKM+cxmXnw4/PSYdy7o6jGYU6PD
wtqO5lGs4u752XgMsbBRPFq3WI0L5lcw5VwD2Ov4IvApSMcL03r5HnrIPVHqGEgx
TcLZMKmnrh2EzLir4CfviGp6HqnCi2Z5xLLqDmtEtGOgtInCIQCNu1i7KCuGBG6a
YqTiKDICyco1jAneQEk/LmYNmpxg2XWnbGNHotVeehx0R+XH+OY7ayRZZbgCn6M0
b5AEN1/ZRWClm5O3LJSK5wNqfmvJSycnlDmswbiS/nebumNTNoQTqIHqR6WzrKvS
o2cQdEmXDHE9p/5IcNeYn4Voyu3UiAcqCYSe6QCdxnF0dOWJwcjUIRcIcKjARdNn
R0ydtT/yNXxBwkTazx5Zik33uFlqrv6jeaeOj7a+LXsSUnYX+ji6qK/Grg51d5Rv
Z3ouajMqdD8uK2odAhGP1fnEHrsz9F2dozKY+8ZtXZl9UIGQLPX53EY6or/J1NrS
fkFpdCnsc24LoERJMjCnb6/MGxNy13oUELljJj6ELCoCUxwgESWLL9n6017Ngjz7
AJ8bK8gZJJZEqJvquTzryxJtk5RHgD+y0OQD5rI/qFzEaPcXLGqeJ//y8im5exef
fvI7nrAT+//siaOjiEKhS3w9kz8lXqb74p07NQoABArrdNcAzx1M1L0T5Ndr+2mg
KS29HHC2alG/rAZ7dNqcb4DGFBDM2QzODGZNSsWuaIBiScQ1o4l9SeeMlB5Lhzbj
Oxc+ZQgjN2ZSXF/50XyfHQVmzCBkWS1n70oUmXvnWRlaGWKFPMOyx+J//U01tGCx
LYWMnVppD+ih9AquuijS7MH8SrBD7XTQFzGi0n4chimLlR/JipRNmAv3HWIhZnmR
R0os5fp2HnjSENwEZIVomm/ZNc17eVDli2lmHVlwJx81qf/cXPZrglX/eyB89DuH
P9gAwdaeeMwzSsOLMdtKfc9fjTYSPxZ9BlANZpwW6JbWi+9KmkzYluLlBJ8xDWs3
zKK15HZtaY/RKcw+ukQ+5Z3a5EapcVPWqz9kwAzWPXgyIeWvOKs5haw0gJblorSQ
K5MV5Ay5dk7pElh8L/9OSTFjXTr93jMZN+BfJA4wOGTr3IDA1U/HRnEEB030eBlS
PaZ66oj60zqqVTGidnMIVRiv5TD5eG96CfEd6DlrGohm3/YXFbvO/A6F7u/VrhGL
w/+PRwM+UP+ePQvHus87Cl4ok4oq5siRWs65yQjDlII/x3gTuQoUivmVU0SqpFY2
gxbdYyq1EOIQNDido7T+XQ1a8cjSh8GxobuBCYXaJ23TJiX3VV0PFV/j8/Mn45RF
0b/iTto5CD+Y/ROi111JvIxQH7H6/0+6HYEqVnRjzZF8X+QlQ/IAPHXkim3DRZ1+
Bt+f7r9v7iZPm3sy8J4/jqAt2r3rH4K4cQ0k9gH581+0iNpPNbJ9TuH8H6Z93Ppp
ycdR3A1u+73ZbnszRqTU06LMqzKWx9mdgJhF8f4Epl6afN9/RP9rKcJvnfuQ4RlX
Rf1YFiHAarVL8bN+k5AO6CP5K6fvdgC34xDwfu5xeF3a2ZVjDT/FevbQUFcy1Jd7
SX9j+ffrnuN0ER9KjrNSZroD1RYjlsyWAhXRSqB6AhktjWspAiHGtJkfT0NHvy3b
sO/t9FuRhevzY544nAFYJoH7RFKg/IoqZwMprwVrK1yCuoagq4CVLmqqqjVmiF8B
U5daHn9Yg/hdyduD/bRrSD08tZp3FR46KOb/A2R3JPa1LmLY9UcvZd7woc4iTdKj
gQgSwg4XB4M7BBDwtFhxVqVbZ/zLTWSL4sioVNojWKsfkaGPgGvqanOItCnCuI7n
xi8tmDRBK2mQQn9MrSLrUOxXc9ByJ36bufUVvRrunXZvfVg48geUTxD5uzH8WgD3
8X6nbc2hH5W2g7YoF3R7wmC6HWTQHDlFuSn40a5sr1uEX/oEK1h95tpHygQsOBrO
I/R+W8Qt94MGNM5k745AGPtnnYb3M7TpGXpjEgB0t44Tr1TZh6fb84Zs0QQ2OO2f
7kgOpvyiKwb2lN3StLkupqoTZqYgYMwPapsaUSAXlhopkUfb71g/8Pa2f/gbnYdf
5F4MAk2lIJ6B0xXy3mCjzBmrAJ28KBYkKihrOegre4y22m5nYKHm2OvGhU4WWZo7
vWOhniXDvkRUGw9/XkFLfOWvFT/XIZt3fwWiSLILtYioo5jlcw6H778bjAkm/8uv
VepdHnVFQYnAAQYmZ6VAtfmX50mXEnDDMYnWNqL8sIMEskAQ2JLnOUn98iPiBsqS
LOFyp8UG9dPyHNlNdwSw+5rGaXAQ4+As4aW6a4fHPMtayDpAiZPtUhIVpKBFs96K
vMitYXuhlOEvWvhLo9Hltv+CHtFEnr29+Di/8j+HwIOFF7JtEcYcBq1Vykf6jN8y
EVXGVqhor/WIOBCaFModpV0yL4RUfeOI78SEZWN4QnVkbV+Upp6A10gGtV4RdYZ5
p+5KKDwdRWd8BQj38pMm99JAYAFLnRXPtZ0hN1xafUO77/8lbcgFUg6NagxWoXlK
Gy18GH/S0eh5hwgEgoXIFpkc3S3tyYhXNqVO2+i69oSjOhBJa30K4uaIIQF1fimb
94MfYpKghw7/TCtZISCFs7ZC4Th9HsTrHwBP/ihm7+x7TBomsUFH264SnddTOziE
+IeCl1RjXIIEkdwn3X+I5Lyb5mtLEtw63RnzpPez8cHVLUGE2SwhfxHtZ4EYtlP3
Dc8tf8ikkl3OVF/+RSFi6h6H9N4InC8F5qCljTS3VRfpWaOfR6113Nab36gr5ru9
gUWhrzQKI1hd6K74KddyUdQth8vyb2wbvxGxFM35rSx5peyLsZhm7wPexSmQATtb
ifStAAoLBI7NsBXCWiv0ffvYIM2hFZQgeU5IffZhhG3nk/1B/7b6Yq4uyPb/cKk4
NsHyymL5xA+jlWa4IEQ0QTw7EujCPz3km2kHhhOBfwNp3qoZujdzWSEI8u2J+nOT
NzEjpUCed49X15JHxKQg+upJOu57xcqnUgcBlRcyorzaW7cky3Ld5mPhRzEx3Yc8
OT4aurxx+7cftdUD4goG8P0PujAWsd3CnOmbXT/eC4Y5Qo6+e59bc4A+w07OkNqN
F/xCDH+33yEM4OaivZQ5iV5gEk6TzfKnhOq68eT/FqJLHotQ81WOYqVcknRPSmHJ
bCp5qAJianNcm7AMUG9ubuQ0wgSfJKPSX2AS3e8c15jxCDKTUj8VjVbLDyhaxLp9
OHhgLQ1xYtKXyTlc4BDlvAKl2BFSrDAoJn6lw3Vyoy69DhimrGw6NEUvTcaG0Bc6
N1ycUpRXhkvPD1bESRbgnEIOpNGJx1ePa+0P48G/eRB5CMXQEndO9KfyBsgRF4ei
LFk/3UKQoIBJdVvtvHDlT7E8Axyl+ZZCx64+ZeKDDedPp492QlZwQfDYfA+MxmgF
pwm7I0mUuyQibCmExD4iFUdWst0QYz95MKUurjFX/EB8fkF0seAz4IFa1UL3Lnfr
YZ30k3vYPzxHIvO27YNMogqS8TbXjZv/b19WGWioBM+S1sAlSLWDQJL2zreB5pL+
Y8W7HxdJ/quQXwDK2504CRi8l31Ts4SAoqYfzk7Z/M/G2+XU3lw90PdcwNMzcBL6
z6MeZn7THeCSz5ZlUhHpykeJF2Kp8anbE/Jcb2jio8VU1iRBz5mqi6EF+wL+l4NA
xR3YQxD/CwuKTensstgiAFDKKLMWNvnFuRT2jKJIwZhPQCeiPQQ17BIjVdG0E0X4
maZGecnttErCIAZrqMBmoBZWa8bZHoT2lYopWzNMRy0b7l2hP4LMgTC0CAHUU29b
eG2JRGEy+6qiZdkV+abqwV4+eD7NLqIWRvf5qfyaRr6unIxz7dM9wqwfgyThfhOD
LnrwQCS+dhFeR2bLMSoL6fiDGJLXdpqw6a6GFnErHasyxD9ulffsfOODH0Fau75+
4+exZ/DkkqjweZgqkSLKvaB81ZOeg9AQZFDoznxmpH6Bqw4MJPt43Qryrh96FFM1
mRI30P1XEEjQFy7PUe4P40Gh5CKGrWJJDhu2Oe1IQz8ze53180lTbnpg205MTdGi
j1FWQMHBGoVRRQENFbAJtRS6PiZj7tOzOPGDRVXBFnac8aDi+85SRPIbD5Wm/3p4
vRWzX3e31B5l0FD8DHbf5gD5VCbpopckRJK+pAVEg6Ru8vwqJU6FmwMoupIgCQFQ
fEQKznmo/3v1LirFQA3DxnJfvDScztl0SbwHmx8Jrhv1ieDEYjc79WazTTWcd5qp
wQiV7HrU5yROQI34FD1KK+K+UDOG0jKaAu214aEisbqsoCD/utN9dc7T225evikp
wZsFDmVTSZ3Ntfn/k5AfzpYg7R7pbw+dWV25h38bVKF5uUtecutLHlqZeQZg6zyl
l/rYogodH8tKLHjClIhVaODa8WRRX5cEC/jqOQ/RunGFfGjXQwmbMPlf+pZL4XaA
AKR2LZM01AySpuCUnKbb/CXQ9ghP1zNGLZJ7WrXqHR+blRynI1MRk1Aeu8K18v2Z
/D+quNJHOPt0SpiwvflFJoXf9LfEHpe6n69DxYtbewdmkDHy3dmmf/wVHa4eOzkb
OUKu+vfHJi7oaWV3OWAqEWKIa/ZEX3mmqSK6mamg94WdjIhPNxRZrfT069L8AjX8
Ms2grYuN5wy3GGlWCtVSJzUzLjqCmuJgcfhig2e4ZzJcjIysS1aipZak9UBtRJQN
qHMugFWKL5NtRJ7C4mxgpqG2Z9fC8qPZ73xNV4WmML8csXfeCxQwaQeqzXSWErE0
ARaxbj4vumRnXNi+qgkLm9ElqAZxx7/n7NeUIimJW4Ycd6An76GZGP/w0tuD+3zT
le3XGCIrm/BCCcjudBx46BSuPOLA5nUer3X7WAzwSqX5OXviJr068i9aINGpF/NJ
XwBLF4FUkOXaM9I4SXCjxzVajpI9K8fWnug8rDVQpVzuMER6AYnyXhkMbbB9A1Bl
4AJtGjli+f2hB3AejdDA7Ri9NMjS7pxls4mVfCLfNRni34dJAWWuUsso7TEusj1m
qbrMmh7ccsMvoor4zEZCzf5Z1LhDAuH8Nj1KZz1n9NVQqYjaC5I+OvGfqhqBlew/
B+U5acvNHhK67eoLM543MSZcaPTbtDVRq9etRbdu2+WuOPy/dR9RV0RW5hLrgJmS
7V4Z1BlZFgUOah/gbIDfcu1VGguZG/bEMxZ3J+FCCVB1u6wv7dGz0G4KOkqRdetV
tcJVA/CXGPXcOOZw2VcwH2iPhdVsP6YuDoxsrrA2MGNYFg7zhoDXKAb3z9JuMCAN
mft8KbJvUZBFX5Ut7jf6hEGeKsSevkKtl+NNG+sgcYJMCR/3HlZgpHGlzIok6zfL
C6nk6f/w0t7Zi0q5ZAeY0eDK68WHOcxMO4FZov2JUE1HGk31r/VLqrTa46hhxdIk
3mZbgEubE1jWdm/6WKSkhhObLVmyAgz2qAzSX7X0YHyfP3XpkRYz37qvh0Zhh1Fd
GOILgz17q24NPpQFz2nhINf2bP3KdkC+wYEXAs+WOSR+0ipykW8UbFmAIZrikUa1
WHi/fBrwCGn7i1vCJ+bjuAUL+6DrFfa39mMavgEcIwtPGFO1hu0Th8ech+no+WhC
siXq9bnWpabre0TChGrdgZphusuCnvqY5HIL0AKJoamK0wAmeHkSt107ktaBaPlJ
fzeyBvsjTVwSPrgAoNRNxG0JUk1yGPXRs1YrIBudnlz7yyjNvxImCHq+vpqv18Of
sLcPYB8SfEJnX5rsvuk+8+MLcCOTJ6hSSFyNpSe0ldj08FNQyid+uA9O0AW5GjFo
+u72mw8t/SMFx8BBuj86+zwI9g8eyML3qiIN78W2uI49zfvm/S7Heut4ZgZHSTOg
K0e5+1BXphG46+O67K3X0jN2SNHqC1OXd1SBpWq92P9ptmRZlCKE1zFj4E0hYMSF
7jHN9pC9n/Mc2sRbSNTP6s+ahDBTy7H5zlGq4s1/Xasq37fxZ+cLd0NvNNAMafYQ
VSw9gpyGZib7VULwv9is9/z72FaiBz7Lkkvf/sg9Ku/0gDDfpUmx+Rd8uBS0rZ77
vPAVJ8APQxPppX3e14yndVy2kRvEaDKKIfyfbAiS7pyF9bmtgJdE5tClcjUPKx5d
n8wNIPjVvCu9l9RsM9FHJDb7MDr7qvJhomcqBZRygU0fXiysuzoVLAbeXVFZ5e0I
NS1fOrkUQU8uJbTqMgTSQHZNzg9CQIwbUgR1zyTWNLkRkOAhh/6OeGf736FCELua
dhwkrtUhqUHlp5T8UEyjseF0JJxcoyVsr1mF2BvubtRufNVu6XI4eFyvf349NvtN
YRq93YEe/7ZLJYI7zIZcAoUq8+p7pTFHiHYkqTFsKW6BqOREKpiQCZZrcwYB6Hv+
WmQCoRfbJ7nKya5k4W1UtUBSExkAFkEFZOfRtwLUV+Rtbk9Qu1fNlFgA1VdLoOkQ
g3Ao2Ekf4rLOvsT7lGs6QbPBPcp5iOul3jM9GtZGMmOdT1rZtPL5xkzj6X0uzEmI
o1DE6aYBdnbU20HnZnpCIkqsDvMA/NhuQsRhdjROj4OijsjN5locaLwf2WinJb8c
NJh2ffzTMfD0p2+RbE0O01TeF7V0ekzHWc+gRIo4pV3TOzFcPKCm7FpT9bwXH/KC
3iGUZQNexbJ/fDDKzjiMyBkfnu/09mnmXWhckwKolgqrvJJWkptm95EcEtUjWwKJ
oMMvi5V+fuBHksMh0abCk4LzUpW2wmGtch2aRPDaLUCuHKNx8UksXCie9ibLgg+R
06DloliBUO0pMwu/YcOuiK/dc/XTU4MztEySns68dybN+O9Q0Wwk7BTB5mkEPMUS
CZbPKwKxzOXDzKhTprIXDya6qmX516zXTw525h849o21S/85PWl7OWMN3io+BAFQ
1F4xENOY57q1QAyR/u++/MuDSjLOS+UTahxigkjEmWMyxBvusJc+j+lM0rbDeTpa
LQpUlRvhI+yQ9nLjkHCTik1PtrmA2Y33cJt1dF8/u4+4Bz35+ot9X+VPEocCR1qa
x1z1meihDnXwXMu6PKyszDvwm8OpFacjhmdI7DIWJE22KPicTFDUpJ+CNOODJUCT
FStAo3AtgXlv8bF7gCY2l0fapg+NYI6o1uD8Z+niqSuiEmd/Slnf2ikstOgQFzs4
9IGKztWbZ/EvcDoSirXCLpgnBPNI3/0p6JNTUMXb9PWBjvtpokYMG5umIDp5sOA1
THS90gDVtoB0vH7N5GJRQeDDTN/cQAfcjteSOV5bP6XdMkUhIOkXVvR7C9IZ2LCc
fXmMsoZ+uRWWbhACOkctOrwxiHQymo1H+11kD6O3oy03hhPH45c+rhj+dKMEt3jH
trL5KK4URmxirIHIWceYhklm6YE8o+JtKj2BJ3xZYS3kxMozhLuG0gi5ZC77OoFK
jpDUziISVdfVlwd6pV/U5rtfZBamt1Q2UF20UtWujNab1zEDTml7NThBBhSurO+j
WFY2Ll+5j2SdqNRQZVRTWkevd1qwsA32boHKsrDathV6MurWPal6ISQsMTBnwPh5
kHD36L4G9Xj5QTeQrCw0jBSa+XLVlg6GjvfqCdv/YBw5jWaKLdjaOi0pHCIS5RD6
VFvBXd/EC8MkzHhW2/Df0FtV5GTWDFOXChyxRrdqRaNUNk6IS92yEDedOUzLMRcA
1mHg16fFg+cqV23QgRSo8VGmqj6KCE/KODiZNraeZFUxVjTzc5+Z8jDTqJ74Nlvl
ho81JYPus1wp9RI5fnKuXTD/Ncu1nnuw2AdSSy2Ls9SP7w/SLpwfM6caLWPfpf1f
LbZ8UE2zcikKcS4t5VEyvy9f0aD4xMSdBxIGTjRwGehrDtlWlJ1Fs1lVDxxp+bCv
V4leUqtOFecB3DWv2rjxu0KkXR0QyDomTzX1C8hac54iHMiFcn4iYM/I+qfpgbqw
tzC4BE2BJNFvFVe8dQliYgTiuOzXzyTvtTKDvZM5CjvBEgZueM7dpdPRKWWVinva
Lt4jNkJdxYYDfolFbGQvrNTBI9BG0/DI1JaCikGi3eOuVXPsFMye9L96O+O9EpGO
JLVY/zx2n1e5lYcWM6Gf4P+0nC/qtACUqbgvQl5WN3FN/9d6FgC0gUxk8P6EQIhS
8/6qW6lAKDoWATl4Q/vss/yAPVQmTF1sXI4hVu+0uH/EieOkNf293R3yb1qP6w97
ErqBHbWeBXYSbsK5Z5X6gNi678fRucicVQPixNHTI6xLU789i5Z7RLXC/F+zgwBl
VCN7H87CFpeA8kBoDCz+QYAFVX8U8ictUqw5PWP4zJsKWJgc82LjH0J0EuLA7g/3
R96VRQKgXatTYC9FShp9fDMk7gcXDO3NiXVhhnqlxIC6lSjT+HP07i+xFal2W182
id1luP1nyrX9z3HTEPmYc0uFU1mN36fQ72FEmOla6Hwkj2ntL70RnYeEYfBdvpaV
HYT+KsPuk4iJEEEw+aZObwfUHTxh+F/WhQDWASesCE9Ra72hRA6m+Sr7y2FlO5it
KoTf5W10oqzGh151aBtibovr6GnDJ63OTYAqkH1C6CIeADdFqT5PbvJThVgK4u+S
cDXmi9Hjnzrs25DxJzd+HCjidBmu24LdLik8fZXqjS2VTR67m6sg5WZKttPzvNol
+W/gJz0CNBRt6hoIXKADAW/J7gOwDaH9gByR1/xuiejZXgcQIbefPgzHMvbClK/s
cTiIOpsFhxMFiANtaU8oeW+xMZwAdJptdnSjeZeo8You4O1iR7AHaVcJ06yFMhB1
hUjvgT1fKFNy59Jhr81/U7CF0h8z5CQ77zX7NU+OZz6yasts0PxPjEZSVDaBGMsL
c9Ak1R3OQH3ftln+hRcSNOoDkB15QTpjiPuMCEIMH6ziellxDA+INx3AaGSBd0dz
61g5kKzdPYTfHSGZlfQvJXhv9xMfGD/afnujCMcBcrh8+pHHnrKcm163qEPwrCLc
ThRNKtPEAtWHl/PHWY3erpCFaEty098OL5U2kTtU9PzgSjvgY8Hk9me9XuFgWxiN
usXXHARIpsiQfQx7Wl/fcd7oPsnrWQhp6JAlr1feqLW/2531cEQTCLCUM0qh+oOR
xinDihkrPtHuMnPA83HlvEy3A9SM8KCV3HzBxUnjG2bhSCSQBRP1DPt30a8hZHy7
qMjxS5SeqvHleEe0eQ1txecSU/wpSvSljD8ce0A0Q0CAHQ5/u5V8q0gU19V8RDEf
5aiL4Z6sAg/O0fT/BGTUG/Xd1kvwpOnHCSzTVbgrHOkd19hSEIpuOluh9CuKvXAo
hsQkiS9TYMAzsSwonm+mlUCB7DB3t/KPCEsq3MdmLYTx8MEiR4Hrh/QEnFOnxZsU
odA1CUY7zKJis9iRywACHi66sOX+sroDVRlaKbgRXby+2Z41MLzFQ+xLdOanmSvj
vH93kxtZJQ01DK3RkYNVUduxQY6e9l2nO9eYoeGoSCuNI8yw129wIhN4WG6f0LRZ
PEzKxZPiq+Clvw9aYojKhcJtqCUQUWeSDt3xquXUD+oAbtb8ok8T7+X6BddZV3Yk
rPZ8rT++sudjjScWkJ8aRcFpT+3zE0ZBETCXDVvpk4jtY3eU7AQ3OrF5p1BpilG1
yxKkp1IIwW8ck20WQv7XMEkZdrpdtFRcE2xA95nQbokX6ceIM2FsYpRn180jHeIX
/XrOF4eGcCjiNCapQxNL8dcViV1s6U+5p8kIJkavc9A64INeHtBUVuBogxdw7Wrn
GcgMS9s6P+8aDJ55HtuOFm4U+Q2t2Hba9UhG/bS7f4p4f9IWTQYLeKIuryGE2pT7
AR4mvo6eygjEaxszH668s350PYyd5FwHmg4EoAQrYCA3BOChHXhzCshITsDM+3bx
PTGM6++2pCkYO/ABGwnoxpgHoZfU9NwEcTupLfm9oswhCeZU9C9Ak+2dgztrP156
i0tbhHnK9t+l/Gfonxi8oLTTsE66Fl9+vFIlorDll8FIIH8jwm9O9GSKxcLH8Ewl
a/aQHhouxCiLDarzvQvgzN6CGK/8jzu4IaCw0tchrLa8kAiUN+1lxH6qciNQ6ucD
P2m6BAOMRKfpNiqDBxo+YsuNvI+SWLleRW74l4B/OWvJ7AyTaCGcC4z/lFsCoELg
RrYK3o4eYxk4K+0t2jAJy+z6zNhu5oc0mdBqB/AXzYSuMckzn/JPgsbbvXokzVlv
Oh6nKLNkcuV395Hpbwmnb+NoHfZPu4ndwL+OCOuYG5ftADkG4+FG3DnkKGF++3FH
2EoOvkd+PPzcEgpo2wgiP98VppbAgwzPZakW6dxkCButZyGqRBNBxEkDvxwGEUUL
XPX9kQCd3YtLQzIK1JoUQujAyqLenj5unthysPYLs8FH1jBoIiEv8mwnAAflJDtz
fWyvoZPI4RvuxG54fx+tGwiAKDxMMg/2oFsWVyx3XQvySClzh5VmSPKC5eN8+3b0
L6R9nYOopbwzUPyTkG8w7jcCgRzhsQpaEEAm/ubU4nMniRr/a+anQdC+vHtDZLHf
Wsi3NlgIXY+iUG6dCdk5XDXKiqG2x65BJSUCeyUtO6KazJsuat5dH+PyhGOueFGR
fwdjjGZgQAMQDIEeOuxB89+1t/R218QT70G9LhbZ1BYtgrsVJqqnIkfrW+QBNJaz
hhlnuP6QouFAVnmkCHwbcYi1iEmfLPI9XJy5tNxQHbAsy6ZHIgSOttM6LPI6aiy4
XComRyiX51KGkrpIZhnvMMQv1icxAT4KQ+qr50mjgiOJ8BChpyGhllUMeaSfit3T
NdBH/4c2NxAVV+mnVxEJjQSl83maQbRuLg8YTeDOjshNjIOdITV9HzInbiURFN64
np/UfGY0hE/teeWxBghFl1meui8F6eVr3P7mp9Ry98sX0DG7b3TKLkc1vZLcdjmr
fv1JbR+XKfcMhf1QzbcIgoTDmw7ZV05i5ceMrkiJPmKCxoNpFVlaIoYBaNxlqS6Y
JEgscu7H9p++u45k+gneKFMjY+AlZoU5gDpvYtwYeBck/3jUIKsX/sRm12a3doXI
E1ayRIl6w4cRpgLPYfLkithqwOFW9tMUGwcihKnNG1LYpj8O6F3QubVx4DJt1XkN
dUuhKR+659X0elXhdrChu39ybw2a7Pyy04zh7t2iHmFd9mIpfygdzs68tIX0wS3M
YsaXmm8Imlnx4qsoyVKCAWnlePu8XynIX3EYCNoW5GsC95kLXXHAP4qmXFbAOSrQ
xpj8QXSK8GcVS5CCwJs+SuF4hKlxZg0bY7wgMzuYvVy3lqqviUmVjvJkf0mfM+Wu
RFxJin7bDtUZ42XeLGZpvht+b/VPP0oUeQsrNGLir4JSZ8X/4LV2KEDOIEAUCoL5
2KsJzKBcR1TGBBS+OkYMy8l+qc8RlFrtZc5d9XthaMKfLZfay+qm8OoZJCB5aDvN
vQsJ1r3+RYQtBgI5TjEBl1Fpzq8wlTIBaCy+lG9I+gPLjaQRdfhES1IYUwZ4V1Tk
ew0fIRRAtrc9G2KhwM1H9OjtPQXAChchxiKCh9VD7yV17dxypX9gLzFr/204Wxkn
9wdeJ5YskmFCQo/poB5RRzn3rE5JnmTGfbWO+K2YDLA3tgrvDMWn5WbZ3OayZNCQ
OaGRLbzPnAMRGPm0Pp/IcsfpoEx0Ivo8/Obcf3weRmPHaliVRW5iyqtgz+dUczMD
dOMW8pOr17sCI5O3270zVLX/2gdwl8lrC7IQG3AuvMdzGAfhAA9Blzi8Se/5AtPL
vL0LNAOa1QhIA6M/GF+qpWSEJAyWHn3wwl14wx8kncA81+PYzZL/WN8/+/hN2gRb
y0s1u7jK4R7upNYg2ECAKpivM9z3mJdw2Bs1DT0NZzud5LWnwDu/RR+niBHMCCO6
oWqE5geERuRqk//Awa+/JkxX7XtyR+1u8oNEmG0B+8c1kD0WJLQxieCZKeirLLMe
Sa18F1N2T0tAGcQJFg8zTXJOHGbijvh8u/VgGidnOe6RveeM24c81wRrAmGA9tl3
34NUou9WS4ZHv1h5N7xZAT9/Hei8Md0kHE/7q38GoHd0SbAOv8T0bcclW+Y2FAR1
wMdBoJXy28IWNlpVVre8QWBxoleUgZdzheHfu/9gd7VSxY8DFSWJaOI3+RtsYCMN
Rvo7cRhL+2wz2f6HMfWJZ06uNa0dL2YonIIqDjt1OeCc9bXRPUB7FqCJTfEwwgVj
6WCiOkQ8oTYsdAr/Fd6dpKmUHljHjdv9qTGj8axuobB7SHT6T9PQqhwAsivGMclh
DdcUK/un59imuGrCw+U4IiaEo3E+krLuSVAmW+wFg/EePMEwZC9yhjmeOdM5GodW
y2c9T7z6ahPy0uZ7ySTkg3t12mtmSfW3JoFktmYNiTKX68VtCPLeG+JQ2ihnMc6K
UbJHTPj/MsXqlKOi0smIbPkgpqiCotaTz/sChkRvaB8pJpr2UqCGKvrPF6eyylxI
c9Rcqzb4UJWp6yiNj/oFkj8jMQBaX5LrAmfGY42tJC4tqhj9PB7of3D3/nqYe8ji
am0G+Z6BaqUphOOoci5ZmETMjiUlK3TS7rW+Rd2mxK8rf953xXH4YZWZTYSncFvr
asELBadthnhgtOp/ZVIfVbh92e+OyoPOEw1NLV9DT3qHkVNNrgXSzyOCiwYOQoTY
rCetD7tiSyVh13bIvRmHJH/6BUf8ip6zrTKphXS008j0L74VzFZRLHu++XiOxpEW
MXjphrleOvG53oS5q+yCf5qKO2lJx9kL9dr2Z+3bUI3BGFUqCA1S4qjYj1627Zme
6ITT/2jJ5zCEHrUSqIsIPO44iOQ/KqPFM8ghhjZEEslmkKr/f+vg2GQUrJje+5lR
VPA28OGgqdhhrM8q1FX1NFHsv+ftzdU1cnfFHzy8nrlhphw3BJfVEo2bMo6maVav
JHfF9Bzojz0IvPKcmx+D+5ZbLsMWS5cVLeNREtAdi5LFjGxeScHYqAh4lovozIh+
QvKMJOjiHTXMfTbgG5729oTioivIzdD/Ti3+WXFAA2o7LjXdd0jrvGBrbu/ZrTzk
fhKfAedXdC4KzIJrUaDEAZDeVD9AbR+FduxgCkdQUb9+MZtH2fSCVTZyZrw21pIa
GspDS8Ptj/7DgKiGCSX6IsjbjeoI6ASfmJvgQ2WF8q7B9DG+cF/8yqI3qmrPofrf
MaEVDvGCDCs9xMUBXW2/OhASn6W8QfYgf6U5eNTmbEWOB7qSNeSaO6rBHVwZS/9K
pvdMJfiZewymfGx4TFb6nNXG1EsiP/6aJQPm/001Jiba+6pevZ6ZXe0W7cjBuPNm
M1rek8wMNcusxSJTWyKD/8BR9HWj/3iA7WRhdMFC2S/FVgmIXZedwhAVzyPzqd2U
j3jpH3uOpCeIPTFX7cRYiCzbAMJTeKb64Xv0SsxcUcdXbMH15dT6QDEQHskVdv28
U1Qa4SRnAPM3VQe10R9wZH6+MxaP4iIJ7IxIVfLD4uhGZt6M9Az975dqJRzZ45qJ
yeKmCXjacPhXJvIiEo1tJNo/Aob59zJoLs34p69zOYbxGRkq4SECqkz7Q9houV3F
Vr1zLAljBruNf+XykyjvuAjRJ/c2MFYb97MXURHqn3FcrPP1dysCeX8NTld2oYmj
+eVL3SLFuL6lNWAlDNh6KhW2C887qoru1hrx44PVfZJj9qyN2SWUSVx2MT/N5WY5
GCHRlGJl2TSYVz4fWWbGcPecOMtmyRJ6Iye6/FvzPfKJf1CeLgiyPaN1o5ir32bc
GVawvm8NYJCfNeABrJEG1WwME3y6yG2s2OykuSGq8kWLY7GMGiEB4XQFytqnftnj
2eTWJ6S+hgMaYHSQFd+UW8SgXy+PGnOk0nKvdSm1S/3Lyc0jfqDaEbuOd348HGnD
8NMU2nWpIqOKlNflmIIRQUblXi2bspTNwRAiLjf97IyZd9uv2eXgaD0UuGZsKbBM
ZFLRpsqCHtyCCX8IdzQWBPj37hdi+yzzfoBawla1aDOHK4C1rkOgMpGVWoroD3Mr
xeotlD66JTVwnz5tmCfJhn9erD8PD6wysw1dTwC2UR7M0YGr1U/hYvGEExnynOUG
SgTfd5nyPVXCobSEiOjxp0t2c5YnWhCN/fetc6bPSauUTJ8q2GKCmja5E5ey9VKR
emRIdIwmk1TexSfY92IkxjfDlpyMuoQIsrK6pU5bTJFF1OEIMNzHa9W/fXqx9Ul8
j6e0b4AuFpBkZcdkaCAXJuYhSV9CS7R2pcwHQTwzlgpf898/m3NuEXOMYIM9tlsW
uriLZ3wZGLHZvikQohfzmm2FC0cdhdk0HezsjO1X/AAWVlVtrECMriDuvNmn6x3F
Pp2w6oh+UGZHvcZ7X6Nr4eHAqTxI2Iz2NDIhGmmgsgUFePBb6dt7oSOKVF92B38R
+bp4jHIUKxx2F8G942c1GLwNUYin2cnYm3sUWclBeq6O0PEKnlDLtR0q2k0JxtHd
6bcbg2mcE5gSdc/hvWml9mt9oKcHAFNx4/dTJe5G+hM65qbAwKi2hqj2uSw+ko1v
uuS1AAzjmTBaRRC7e5kz1lU1JAYBK7nqobkrQroYNzPnXQynn4GwVXDcK+yD36ry
XkSLrDU69GrGCMfI7L6b/HQns1AZFpyDgQZv3FA69EyEL224BZ7cDGN6GfO4VwZB
v0syPw4/eSmAjlU6oYeWAOcPALgNCGPlwN6cK0BYpnRLZj27abSAFG3/PPVjuqG6
DDJl4m2Y+CbudZbwEPEPTuYBnRo24uzw4a1dNqjtXIfc7aYx7t8bhdVzC+fMR5gy
V1F99OF6Rg7eKc9thnUIU7lXAUUpkBUAMxn+wZuntU5RXXQv/lsiW8L1DcdlwMwT
Bstf+MBb39FQ4Ncs4QMCtgr8sc2O3yO1XZCV4aiFLF2WlkIXPV5diNUQFwNV2ZrY
iNWKzNnvfW0K1LQZBJFV5SCUE43uHf50Af+OVVE8zts5cAKi4AnL9TgqFAiX9R8b
za7aSF37//5LGUWWQxLC3HK0qN+N9PbtZZLz13KixphpbVnKpkKEQfe3nyNdebpl
kv9eA7QwHQxk9/Wm0dlqbG35XlZA+PHpIGA9pAzGpxv1vCjP59iV5B/iCFO2Ev41
5V5dRYKECWW9i+erl5rYxBpBTK8yIpuOLeGHPena6LalFcA2SEhQo+OqdW7HnMct
X4PqROm0OHdIbufzb8V1tN5CM5iNRjJDu+dBYYklDYpMPc8o5DB62sEmhe02gqLh
LqckDIlq/FvVo2BSIu+HMmN3mXTYNwvPYjKF+7etoqdZ65DG31l1/WlArGri1lA9
CLgoTokzZ23so0li5YyndM0FokP5fDWLgcl6vWQUJIoKh3lh1VUc+zY5Sk2BuGRB
4jwB3UxuxuTBS/bfD6bIio/1SPRBFGYrqlDRtMqWG9z1+VDSw8S0B7iYljhLWoti
gXPI8n/+HKmq2J4rS8SWfe51V9CCnCwEkRVSsJpCtcBvVMDPo2c/VOEqA39PKj+T
Uz+vWxwERoA57L8uHM/Nk39DsI3cY2IVdpIIA8Z0c/rUbfDB6hGN5SW9CET8OTaM
Hs43+bLtD36GMqBczcvEsm3/RLFbV5sxbWFpdnpE6wZ4on0lnMEyUs8AE/PDgAvJ
Be2e91+2OXH1DoLe/pzw0UsOYkLlaXJGnBFVySfnRViOscXz4Grw9VfO+Wspkjm+
P7H3dxCjHRly6MLu1tzws01rpbo8xvgREO8qXFpza+t9S+rg9BJHSKWaTjX3pf+b
nmJKYBIkTTFXBFTGo+0M64zQqIVu0AVIs/X8e3JrVyS8wGNej371SftePR4WqIs+
/l0fReQEr1koI8OGZ44EsmfPcYQXdoLRePu7ljZ+m39JBCqt5bBHhnBpu3fVYuQR
ZvGl3Ue5Qea8REpL/2g7Qdxxqs0wn2LumjjVUfps9CIE8NsWMpulZDbdCJWvgJUR
MsXCk0PBKPnHBUleajU1YQciOvEc28DxWlzuAhHuGfB7JH0mms8P4r2cC68PYMjJ
+VYfsg0Dd8w+CU00sDTa+/4O546diZkW+MScN/M96YWNGs5dEnlFtBooPR5tVxf7
2ANT1T3ZTX29Hpf2WnsXh63Z5h5LCEtFJomfl3APXnlzPOfBaNj4Lp+EssC+EcWa
IYfkvFhOP1GJvIgV7YucRLX1MBMiEMYS8PO13MWF61Bp/Hwz2LuMA0X6l7wzfzZW
CpG998W/Dc14xkuBA2bx5XgUm94gODc7XZLYYNDFOWimahUKZWxRYVfDZ2RyAi1d
JWWvO6XW4gACcfDaFsPQd0gebmfrBBYwGuDsW78VZpcuFdoprkh99LPhaLvg+uHi
U3Cz3cnubnTEFaPOHZMRfBOpQ9bHUrms58cpDAT+vJfVL3rAjdP+GbwaKIEMoejl
6xn941iTe+DUFeG769aXQ4GS5cXMLxWMqxkqdqI309+w0g/R11kIrer5rkcHAxK7
3LrMR+5FzpTVyXPJIozyxvL9qE7UNOJUFGqLVxb7pO90qouWbmdipFHLw05mwpZ5
YgqRf9S/SMONmDVbvbilx3lAXVSIprGvr6PPWotap1cbPz0Lx5YjDqCAkpW+lLNy
9pAkfEwXgzT8pcQGzNsNcNPvULUXyjTA94igJ6oI/c2OjnLKe24/Tm8DitQ2dHAQ
8+q673tXnEDlZ0trLVKYYRSIROo5FUn99Us0IJu549+6LJ9oGn1szJDDeBz0Xt1u
NzTnKtFSRZaUGMsImgC/9GnfobWGEKFheLK9lCR1vewVp7/OHfKX+2mlzVyiPV8l
XpRr4ygUf1S1mKTUA0Qv7+VQa7ueCvE3JoTH0cXthbgzdecT4VXA4YXRP6s4cGFM
jwjY+Y6rAsqda7mgl1JSJtMOsALzAWBgNkO5kdVaoTaPnf/9umW0NM8mh+qFGToy
i3w0eyeiWTgiYsX1nuR2u2uVGFfvJuopktFcr4H+IRDs4GqFHDIfd1HK2IR/pIwi
tk5RT0BHHyww9k4hTqE4UH1tczxqCjNAs2S5Kf7hFjXfmMPBiz7B9HZuxWe+tx2M
vIsxMEXo52aGxnbuVmWMuHZD3E41shW1vuvo+gw4+qnK1RQoAzZTWJCip+DL+NrM
dNy2hxqwXqYvRo3HGLEmKJ/xN2sZ33kzKO0v629JepbGS62QQsmADND/6thIWa3d
kDWdxYAgKd7qe1XwkYKHCPL0+nbe1VY63wtqrny9kbdhy5xoNrVznZoJaHd8Q+76
lhjcXM9MJbegFS9cPG26k5+E3KdAA3aiuTfw2Y38uF/3qWE/txloDM2xopltamso
Rau30fNs2RGsQTW8ZLt75CvIDiIjHaDLV+ZULzhe2thhEsCDXScD6FPEaJnpoUBC
LZmGA3mxmi0OMjKOPUXCXUnun/qqeMug58HTsBkIPkKwsuVy5/cmv4ZlV81bfj3p
a0ZBwO8/XiDZKz3ZtUCyQa3SSw0X7oWkutU5ybkAbDAabPjGEqjmPEgJES9ZmSbL
j88iZbqcr5i+C2rNf4VPJ/Ia+WRF2miQLablWfLuvux9m99IQmleoSAjzRqqdSGr
SWWgt17OwL6IbARzojwFqTunpxVr7oosh7z1t+WCnhCgmpm0XFfH/LjXvwaRvosK
c8lj7gaEMsJtaNEH1rqoP/4Ku5VJLbfOOhCZC/TAlwDqf+dpr9Ne0Q77cSIfke+L
r1riJ9OFwl1D6HgV9c72YaxRqIkYllKszWpI+3XP3Ihb6gWc2QIJuwisw2kJrrPI
I8eaoC9THTeSw3xr06foEVZvXWi/YAFc3iKSTRBua28fTTlPSD0Cox6XMLESjrp0
iZHJSkGuuquBfVXAbr7OUXcEcgFpaQgtwHZvcf1i3/trR4F/HNfSqx8LpkjJwWji
5fZQdGpP4KX9Z9OJvysaTQvQsBD/lJZQ//EQQKnUQ/jMnxsmfeLNKmwoxtnXkz2j
e+ckmILX1Qsww87HzlzAAJgSLkCYqX4bu8ntRLO/Nrj9DOl5AkecKRBU1rX+XUrU
JL0OqqbsV/FguurEfjBqE3XAOnSlWefLWRJildo8GGyDAbAkr21eL5Qo+rZx1GWg
Wb6Bz9R9JJHeURiAHRU9GhYqLDp2zkhP604W68Vb0xKHJADiPLANZI9/74r8UHD6
PX1HRfXjY+XzF0VT2jsPg3+7xWpij/4LqgfAtNZ1iRc8R3U6/HjXp3DTlvxQQOSX
qakbpG5eMYA46KdeRBIrDCO2WiHj2Oq445gDOA51AJ8kP8gZl7fI3KzQwxhFB8HQ
cDjkxo49xEYj54uFM07JN5XOD7CvkLdlGUZL2IrDW9O6KmQBNwJom118eT/QGCfy
Yh/pcGLZWWnRyXJHu08hnBTUkvXU2RbXLglE9hukROHruOAqtN15aLg2NCLvMlte
l0guVqwwbBckoQZ3rD0lZls+EKiQpD6QQYK/iLVu39Cv2miVs+j/4XPq9MDKa8Ht
j0jJ5JO0sewQmuidtcON8wV0aAhTsTqN/J7nu4pd9T896Fm2pwQPo1ETjQLb5wwf
3AOXhvzv2U02rHF/I/gz79MP8GSxCKQUccDIiykf1t/rga8H13i8RQ2mWEjzVM0S
W+6xkAeLkoLyFx3+9R/vSemNMHnSQK0Q2MJwtXi3+F0w4g0hSc4KyMzgz5hcgsdj
6ypcG54a/NlHvon7HlMXilth3WrlXs7MWwjqhE/ofQgpuKSNUQIdQbJOfU2i8eRF
KwE8yhYXXUNkf1CxSaRbM20QqGhX6wDuj4u4NqjczC+lfFbZCr7c5vHmaikoMfTl
7tjK02zhGSmpumN70xgWMa7Tl9R0ac5JnkNW4krL9ZRJ3iAV6fnMsauoYxuFIlLm
ovS2EdL58iJ4bhsaCVfuOgqTowA4/9aw/HaN2zvHh52Sisn0frcYPyVqkZaZ5Ppi
cUF+6qPde8ntf+3d061SBDI+K2MZDwJ3jUWgHUKMsJwsv3YKWvucQyAoCSKk1sJZ
+S4XjYur3ke1av6+WHmtEJ4cu2SSZL2YOI9i7m6Aif8YRtT+2k8lUpx3e9me+Etp
hHMCIM6r0Dy4Ssn1WdOa7JcqnP+opMPDhWEq5S9I40sbRcDWVFJZT0YNpK5AFFxY
trGw2V08YWS173TUEl3hvl+0EzDYwEL0EVu90RqlY+pVvx0SDEX7ZoV2n+v12Lbd
MLrhHu1X9F0TPQjwzcip5AcQGBceXrzJp5vHb5Vuud2IjeFRQc2o4FHKnJfFyhAg
B/n/logtCf7PnbawRv6yjlCzfsvSTljmzs/J2G9K7pPnCiUHO+Nhzo8bauRRgYXQ
vb584aN7kG7s5n5dIA6rNRW5KJZax4rKUyfHIM3hUsC4QhxbYOXCf8HWhFmdUr0q
PRT3y/YUcRbK88lskqFRj/riN5lbdp9KoOhSGUkcyzeW7JNQrvKRi+x72pomRtyZ
aOLeMcYpl63HPLDi7KACnmOUgwsUslutKA9OPNlvhctOp17+10bT7qX70uP//X39
5E0oNdlywooH09o82nv2X4apbwaX4zZjWRlZiQj9SfmKoRg76ZtszoOGldX3HHHq
wFCmNGtuqE5GS01S8FMMLm8vKWOm0KbpVhAxNYBfxFR1eN0JR477NZMPe/0Y+W01
gAGqvp4xxgjCR8zeXRYAgqWm8MMt5dDK/A3YVqW90IzcKe+Mz4D3eSeTaJtL/k5P
C5S9O2zdqz6Tft2NqzJcbtWDL+8YHF0K1KvHYzAqOR2OErEqx4Mqx15ZBMIHP+DV
X2yYXR9IxjnPL2RBADCnEgU5SfI9QcvN/osc9wUyhofngj0JW4+wRc4VxuoV5ipo
8eFngyUD7xVN0ugPDbXmUDpwGbE6HdHQc7Q3fyseA+AOUDUruA3f6MAxgCZjEvb5
SThfVonhC8pTnjB82ELRBFmsNey7NJSxYfk//Ie93fwb9+RnU2uStgMQpK4RPTRu
/d+BQzKEr1DvvLwYpEIB2m1odcVBy3RjZ92hgmROblaXO85EQrJDJSS6Ouiwf5iP
F3UllLy6AIoefWbO8cLV+xz15s8hvRy2Ul5r8Kuu7zzYw3FOAmmFMDY7qjGbRFk+
Xn4ZJqP2vrJjo+niTiXCAJGu7I31WpRkaBJvjjpuuKd3b/XcJ8xH+Xn27AO4Pzp5
DCsdCoIWgzP4Nw4V62CCowbZESRs0Rn9mv5hMFJWUWfR3qu3BcK7Qsj5gRO2w36U
M4/36Dg8ClQ4TJ+f0XxHNbTZDRIH0Kpa9dyQhM1QzPmH3SB0dtYS2u4+AvzY6F8Q
eZQOzweyojnHGsh092Iam6VZhwpH0TI/j58qqR8oZYjJtPGZadsT3o+FH5++s0ZX
kgY9BGznO0x/OBoTMhUy12OGa4Sq1hU9L16PXvFYqy9KlqmYfXl0CxcQt5gaQLSG
vfmzUFL034pPpEgoL6upOO2BTVOaxUgynjvdvu/ivlWs6eFLcfQdmpzz7NUT3zXa
9hqmZwGzzrPRl3h0YB/jplHjMQ3wEeupWXr1vzdT0JthJENPgtzLfILYR1KJYGs/
xFWnijZ4ALvDn7qQ30wcbtONwLwIuU582N+rwQUsitP6cE2FyAaEuW5UurLw4weC
ILZTrWPEnaUsrXawFXGK3Ad0oYBbeENY3hdF5M7KZKRx7uUsZe2FoF7gg5zGBpbD
sKVpfj8jlaPxSP/wb5lSRLg70LJmKiOzp+fn2wclvThjjKH3UAeLp8iJ8SLvVka/
StDs104TQ4dRurb7L9LOrfZ1wUqQB8hDPKOK1AdmldPJOn9cXF1srSdvGBr2/7gZ
z6Tqjhw/YpTuTX0AgKgthMTQ/0RyaJqFnNs8U/x3KNkuTS6YKBDfB/PFDpKGKSGf
2zVlNbjcAUbY509CLhaVTm7nF3ebgQVIJUYA8mGRD6n8qMdSSbu2wucP3Iesux/3
xUOp72AePq9e5lLA9SJCxyuy2bSEoI9Lol/zeEFHijpKGNKTLtYKAaCUE39OVpi7
66g4ByjMxrNRIVQjTvctO8KWwJpWCEJ5+NHgMWDFAcXjaTCgztv+ESmUpMxvyjV0
dEqDPbCL6ST12rUBx9ekqr3HdoZ5oHJehiGR58EM0r79bHaUOTNS71pFmyOyOGJ4
d7oYP2lDmhi8fHhiVge3lLVI/GYoI4bhyccE0ILjx1z+EpYj7CgIh8kWU0a+bARI
0dBkE1Toz3bTazAuNPkSxlYxWECEb5swQ65UGmfn7gj7ltIR57QACE2PouNKZgaA
3egDMqsvhJ5Uxalvcwf9QscAePyfzm2pM3rWLvFrm7qwlI/ydSmnLAiakjMaLVcq
m57Ocw1pAXQmhM6mMUDC6BEZ9GzBRzTr04m8Ec743kfOcDu8YT1DxrhT2NM0nUIZ
HaSe0T88Ts/Vq4JIVNJ1PDPvUf3cHc4Ntlev/g0Wo0WUw6y6f7xTDaOLqcKEip6J
7nMKnBo1BVpEFBWtUd5+EdP/GEeYDiuo5ki7ejeSXuo7cP+zCYDvMwHeUFQNLeyV
2zTz7ccS+ugHw85JojpqtVuNamCCL6iorGrX9PMWGfWdRULjV4BgWVWPbSbv4RlL
f3Jsu+SvpNJSmtOAS4rikw8pLz38qpg82/+N0juIdp2TsGrmqKHO88s3+Cw4iZB7
1SDqPqRXFQmFGicbo1ttpJCpjfI2Qmle00YK/mWJCNS5WSVsZ24/LciMYjyrESmb
bZcQVr62zo1r29tfG+EANG1oO9YLU9XFZKzNLZmiQ+wxwFuDMGHwbt7x++uWEDwt
gaK4DB+RTTskbR4V1mgWdwioMbxiFtA6eKJ3BC68YzXHdZiomwX2HK+kcveRK9ka
fkb6GKGPvr+3tWLQ/hueWJiZd03roS/Fyf9KkqLj8lLE1c7M6LinGRXFR5PEv6Vh
Oq0vxh/Mjq05LU7X8oMI5kxd5bQBeqGU8Bqt3bHaZO7+SmBL7N0nmairLZwWu+yj
yyaBRQYArlUz4BzP6sOBue8OH9mFloHgHdPLaoX/WYjdmNdM11T5h+G5Q4h+QiTW
J1US29A2WfIXESEWBc8EwwUjmViVJvD4npHfZWIAVNXYOTcPA3aq4y+0IT/eI1uY
sgvZI+8QTI8M57ciQUikqPV+Je8w4UgOlQwn6eRR/dP/qTTSl5bdc/tK9U6OqcBW
0Tj4mPufiUsUvQlgSrLR955Wo28WsEjjCe34713xlJJTPgurEbN2CXnOvZXcrfq0
x+O6Yjs05KaKDKMx02g6HcxQn5uZqh9RDLSrufu1m6vfKHj3lOKWvS0o9D0MT3/f
0Z+bfjnZ3WUJuTK4ki29bLkbrxUApFVrkwImCkZ51FBIoRMllx8O5OKDCF096/cH
dtqM0z7dHUcx+kuucDsYeFytWRyMJfq/4E8RrYCItDqYk08kNBXHiMGGZg1ZsGJq
xnXZzAMPFqeXmAY3fJ/wJILeZ4YrbuuveoZKXbUknd3xxJ4HuvySlrpWl1pq2NJO
Xi/U78qTqd9LHJVfhgWvp0hLpys2J1SPIeBKL47s60Q5KsuqosxPLpdosB2jTgBG
bYJUpFKwjybYRCzn+C/zlGmhEmk56xi0Eg25XsJPO5vENRApOkUVw2YgAkWFiYK3
VqbHms1IDqpyD0g6r+MEYlWaQDXtSLekYGtU+WMXK0nwtk30dDx6SgcLJQ1maGUJ
YW9vyshbz0fZtrQD+fbKCgsB5mgjjpSGeHbHM/jUM5TKNiK2tOVEM0Kv896iI4ix
OPSyXTTUgmIRR8EMWVgnQnkYjPs2U+rPEkmsOBuzhqRSKzQmB5F/os8E1GRYhmuY
Mx5BRBjRm2q2eN8tyFpf2w17L84kGXBL8CkEFjvyidhpb7CEdh+2rTBet/YwrHtO
YOzBmw5PkFriCgGvdEq/tr9v8cTiUlEn454zNMzwLoBt7CgjUNainh2ITdQ+AXTs
kVa1Ip34qf/g2fqt/KMyu1s2TFI/QKIqJWrNIMV1VhrgrPfyeBm0b3tgVS+WkN9C
CnWmJz9LNhNh32Od6mFtQPSCWnTZvfYBaUemNX6daQ6K5LtD4wjQBqDfeeFS7Ymu
e/BmcskctPY/IiusKC4TgtuFM41HZFM8N8kw5cz7mzWydqnvmkdH/ex/5ULifJKM
dphhtUnqWB1rEAZ3EO7n6ax5EtDE5Ek95Dg5Ij46O/F+FCpyQeIusQ//0Myba5Fd
V3lPI2lHuP6G0QQcODYdyBnZYF7m2kzbOVUMVyGgmlEw0B3dWE7Svaenx6VPy8p5
5gd9mO0iKhCGVuq6tUPa1YBXutKpQd7VVIdY0fXAhmboa10z06IdhSX4rGW1Dt+K
4TIIxZbJ9i+Akj1q+QJhqYbvDwB4lKsVLsIY/fSB1A6EjTe6DFdXgP8l7r/Tn1H8
yRaVsyokSsqLUx+r96vuUWeuajW86PHCvioGde2WDHAsY3WwGEZXiqjjIQveE3BS
gZk/9BETVu/kL+WAN/3kf39ouHDrIngiSPB3bFKBlxCNyVVeq/9+8XJ6pFkqbfHd
6m1pnfzVW0S9s+qoV72eAvCEYi+tAs7TI7KjczrW0ND84KldNL3JEtK245x68KRQ
r5dZcl1bMNEaEYZbaQXImAHtvqqDX3/7sC1S4+MrUyx6uyvQIiUqKwXhthy2CGhW
gOceUKDM14Fio8FcU1tNWmaRn+r/Qr0X0qrZJU7hBET4t/6cj8xdZR3KYT23fD+K
2I1Mz2INIG/byffY97fSKj7gsNieUKgFAeGOO/TTOIieu7OODDxr98rAyZhnDTr9
Ff5BZG6XmXqxpkDFCUgdQEZwdLev8gPxhfzY4cePB9KXYjvXOU3MEpGowrW5/pRB
OLiv8JjdNdUt10Cb6mhFaUSJUMehYVg6uo9USNA8oVEWLNSGojJsY9Y8gSXkcrFD
wguyQLksbZS0yG5xFCBnNtMsyWujjuwmUvQH5MXdeqTsIItlgdwBPb0Muju4+QtN
B4eKMxuoei1/DunZ+RDlai4fX5eMYrtyDM9UWgw2qUqWqLqlvxZRzlrmw1C2698c
HST/Szu952T6k5+sfUCf4dyvVfDwf27HUGAyiGwJSDU/8OzbjjLiBku56MXd+aCn
SwHoetD8cIgUysEt0XMmqv2xkn8o9Lxkweylvp8FiTW2KMbJNdR/Xflh0o9adElr
DGl0YvVfDo1tZdJfu4DNcf7IEHNePDUqWO86/SX3ajVF+xj2SJgEICuTNXtMpBGm
WFCRGdHdfzeCUaB06F0U5Dbu3lCmib6KQEvzrs/WV63Agh1jVDGU13PP/454PDON
pDdGwMTi5LRsfzniyZDciTzD0lSsDqeA+11bpZEUjrOVpjBUc4DrLpHYtNOKrOsS
Z8+zZ6RpDpkMnnS26IPhHUd1n8iJvL4CplaewSkVy+Yfh2lhXpLnmTtRMNSTpDmj
LTTVXI87ip5VaVsa65ZwX9pKWDRge4mzUt/lc03CpQcHbBPKEBkJom3+7Fx8QNH+
7B8Nn+VKLykVQ4VqL2/axp2PqrZIRVPxIcF8dPmO50cIW32tas2TZvWcrw09kSmT
r9hotB8W0ntTkywFRIHxmND3AvVWVYM71twE4bWUNAFpukkvZmHN78mK6mQbnrbU
tX4QJGSr1OLpnoouT2EHntvEV4a2SclBsrQJj7Jne2/JvKHT9htnw9VERlPfc68h
98dZUYXiNjKq8/Kc/QpSvBVnG9cxg7R7slq0EesG7Rud1LDIviS2PGZDT1GZ5zWi
3z5/00D43ejjcduKSBbBTFmZAcRlUxxQyTOgdKo+Tc601OVqD3Q5rrohm2C+Qfz7
sB+oY4ZFU1MFt4usNW+Tgz0bdSw3fafkTdkNc6JDQDdL7B/P3gvC69XUDRnlpRdV
PlUDY2xwDMZyo2r3Yxckc7CqiMr6DUUpRKbvSVPfM+DD2KQbwqowmB+qlbwpyp5v
5yw6ZonxzU6anDcQ0yhVIp3MG8xzPppCNTxLlQFnKIFFOXTfz8h+5MY4QkZft3Hf
9rVqXZgBlXkL5u5fZU0zK3fgarJwzwldFEpXNqj+dr1JNt7qlD0TEa9z6Cc5B57d
CIgGvZCM9HinKptKn+gF4zsyC3n9xNHZ1k6u7EtVHZTgXAoNjI19f8WY6FpF16x2
GII1Cdu5dderaCIwL18gDVd/vlJVeLJ1SMh+P+c4oBW1hTqCSx1dBHzGnUeM8rNm
n2d1UxbvJR9h40L9M542u7g4ODXlhtmG5KAphVi0aPiGEdPqOuh3Aej70nB9vEOt
mJFls6HRmbfXd7MUWeNGlUH6K6/aeucK6Of8uCw5SVNNCbCQUBye/CGrtt8yOtkF
hpaIV+7cPfzz4E40SV0D59dlLds+m+Uyg2ubuNUe3LSHyCDB/XrCU21Z+DpkJvf9
1MU7koibH9K5OyzhHoAiJT7/qq4vYHN+eW11PJMlA0fFsgYFyp1rfIYsnJbiw4kY
mFgYQkr18KJ2YqilTTc3m5OvZM8nhjgXAeCrxairdxNUaPKISja98CTB0bUbGsO3
AGOWHtV4P5dUt5IpTPnNS69UfmPC3riJHDFCCpv1kyF1ZU5X66rEyZpf1E0TC54y
QSzj+uzJ/niNctwcUjb8ywHFlNHOIDOGGHmIuzW01+sT6IiHQXo0JXck7UGyEPJQ
70ZR1LE9edQ8yHx46qlTAVuhsKFkSkhI6tMVDGZT9SiMdmyzl3oG00cviA1Hkm28
O3cFHPzT/JnLB4unmoQMWfaiIFwZrYG6PTtyfZjGHquRnMd8RJP+Tbch2OnPNftb
6eEMeqW+4Nkx7PmsY1MLv7MhnFIQpEbts8ok67nHNyi05PWaVcYDyZJl++fgXx4B
PPqBUkRfcWRvUDEmZE6TCHyIeTCb1VEEqF3Dq9M4HWvuxaKbMkkZIuUvIjMxW32N
8dAK5iuIZEbTYVuSX+kHiBNlxXrEZ4F1npuUxv/CCyfGtJF+fU+mwOknMjJ0lYuH
fKuqnB2kKyn9+/PzXvjcGRckhnH37lj+CcaKMFBeFNIQwixzd6veEN/IdSMaTpyY
F+683xJW35dbmjoT7qnnWpilMicAEkrxhS4WfuxuHJV+uAun6yTO3+bdpfWZx+VA
KqRHDrx6CJG3vLhlP/x86Qw9D1YzVax+E44X0lgbsYEY49V5mBFoS4gjiS0RtiXx
SgOJ6DIcqJoMrop2mh7fa9Kt8TXvI70weK9WkoMc5W1jB8M3YAShO14T+b9ByAQ7
Ps5Erg3LJ9W+Qn07XqtgUYPpp6d3fPHZpyIrvIZrYOAMroQ6tka85zL6XTjG97Lz
Hromjx8Bi6gvoQaKTRAStIqju7L6mKYjrKoirAZS6DZoC/AnXrtuFQhBb3VqN1iR
XrAOfay5VMsfgiM8bFvMoBXItDeq+snO93nV5ykQu+VZJVb25Fzzaxb4zI+7FZEW
UWXdDM9lJK0yh646DvtjR0h/ythlzARPipgL4phJ4XBVvEoElluIMTyLpXXheRuK
hSx4V+fFmhVYQecxtovlxyDoFjqdUEvRai2xURjdsWfFBuwvt7M5mqk3ODmB46V4
pBL72y3dEx8im/NyHW3iB7GyayFkd5viCTFVo27beIlf/kHw68B6oTc44kLWiqBU
qV+FGO1vkeAOYA2Yydise88GddRKLvfvmyg6k0If1iaqrkPwSBI4GWdt4lPjqfdw
zK+HYS68vDhRatRN40cE2PjfWM82HpUIzb9UjU1UWgOBUxWyxNQ8mXlLtsbvoAo8
d7gA2rxHhPtylQywNwPI60G4cMffn7zbahtqvczxm6DBgyFqNsoNyTghv3VzG+o1
+azRMpWPdvEITXZY/tfPRlwGkxx71eoPjGiSNW+Z3BZ6/qvts9oCs4nd0UER++sN
q3uJ0tjJhyFFF2Q871XPslfZLx7BL7vmJNH2VAbJAqmvRNYmj+FxGwm0O3Wz8qPx
K7H/f944JA+g6lo2qj4UVd4MzGQpoha8SSrf6P0GwyLRz11PwWZWVhO12p1u6SvK
/zaxH7Eu/8w+z84Rqg0h+taWsmTllGzCgL3Mo7f+DSZqH58beODXfpspkLZVeeO1
nmCVCW0VfbY24fzRstUcbeZbNcDWHPRLOAWCvPhvTndh2l/6lMpLEf8bIIJQYTUI
W3W5frvdojHd0kbS57rFbnpOh+Lk7j4voP/EJQ7lzO6fwK6cCR6tTp23nsfkCW08
TAc8zMhfJBcDXDtTkBP+RjnsXXKQXglw7ZJu0NVWSH1LWrY2ayi3NF273H2s1apW
mhpvtOVO1oEjuK6R/AUqaXEr6Gucad0Qp8S1zyfnHGjeS5t7lDsl5dfRmYcanjBY
MnXijHDwQYU8l9PWljewHiH9NTxedeDP5jsGQeZDaljEFy+XlZlh2TGmSq6VERbD
9QLPR87msnM95DYRJ5in53kRMN08HVXUt87CJy+QPr/2+SYbhPVXkUUD3wRMPwMw
mLhWmyMkCVZxxR2VmX0CYsnZA8DbKIa33kpMDg+VNsTN5sk2VtmkWf8YCpdKQ4wO
Gk3W52DgF5EvYqspHmjWplL3HL5No0oo0oXMjC2UDIF+nJ4xyqa9IFEvJFXk4zO0
xDKOJClay87OsH0JEIfK71ef2z87N3Tz3SXbrgl3yDCPYctDC+pIaPjeUQpQ5iPP
r15/t5PM7yZ7xILJrQiE/P98LbbC2VDI5awGkvQFoWwaEjwQNtAaBqE1ad0eu9DN
/+S6k6fKRiOTBLmYko9jMb1G148wBrLqGyMcquw7c0IUg16AyDjLSi7XXKub0Zcq
ONT3nIUda7pG3jUlT1+XqUpRlt1HQfoOz4BwdTGLUwZCBaNFFZijQmaz/clD1PlA
JGJaBKTmf5DMR5tzNmU0js7wdg9zXHjKCYRzTWR4offCgaV6bFVpyT86du4dkHcZ
n9ObaT5ac7m9y+5wJNSs49Sr7kNZMA7ngS9EdnyKPHfqByxg0iwZI1BeFg+3kKJL
JB7AgjvBf3XKgXx1jfmJen+JMfzvymTKIb3SsBq4wo2LNDaz/3A1efR2PC2LoS14
fdJv37qPIsq5RL4mJd+ijcIXSZLBTqgSyA0q4Or0/zTlSbXnX34bKO8f2Cbqdg3l
FJenzL24LF8IQeY80/cdDsxer67j+yysk+BKIxUytTKWjjw9z3dAOYcJCjY4Qucv
Dm16QSJ/gJZWVFZ+slOY0UZJYd1jNXDzhRbqFQ5zujM7k2ICa0KniDFOgs+GOrlq
sxDo2iBDfPCI9oS2Y4JmWD0knVxhMJZ0mJLmr+8buVZx1zQTS1NyD62q9mYnwpPL
by3yKQ5L3S8apea9zNwW0YXjfhYe6Zp5Jbu/qRpnz8S0rMKvD3nC7DObkZVXns98
uwNKszndiiGh4OHvjPxJz3xf+8mxLJc2itsViTDjU+crfdeV9NcoQb6F6jrtDhXd
xk1Vjtm2uLISFGIYilf+xoJbXbNcsi4+K8ilsbGgnqXWpyej2XHORkqkgT2jlleO
DKsdYZewPO4rZ43bUiXdE7oG8rE68csRyrCoGPg9uEmCXMbHNwVKCIPz6xR6nx3U
nRzu1Op1dRW68mkQUnNint+9ca4koMZroGliRgZMvjvlzf2fMvv6vey2ys3wf8H/
XThso0t2VujNGFhvNk/cR3IRXV5TUuTSvFweoOSy9zcGusAmMHToD3jnjSEL23rE
43j9ppw2BSk0TrK3TeBVsbHmkbzv2lX2PGD4EU8VTGNGBi+NmiBTU6T2YeDOFt6d
7veysMJu6xLS7QFCJnKkYColMPQ1rpKkLFaxX8qP6mDb7HmX9m+GLTzBnynHkOVN
WhhlY7f3SP7cW/hSNMb/ZBX9gFBoK9vq3xiqMaAG4gUge04f4WBywat6LhxDJZ3E
wJumRi/hrJxoqmyImB9VQ9Tv2T+b2OkPiUq7cgOq1+7JPlzBbvX25RBhG1oRp7sg
08RamrKJnOm1e5+2anjeI0fwSkoXebQqjboit5yaRhzwirHFauisNBEIB0lK0zU4
K9aNkBlKZxSbMvIs4DfBgxcb2LSfJmKG9l7yfCq3awJ87LytUKRjlfXnn94peV1d
09fw+aRrvJLOLT5F6YjhIMAOpYl1GhWyJzRHBe9Iahl9kzPnJbPAdXEO54kIRzQY
IIX5DyWVbFKABwHUm2TbvvnGimGBidEgO/xFAXY2JTrYgycwTgy+YW7wR7VDdPks
sYjKOZZOPF+oyIYMBZPMBN6CpEd6pn8CyKsfow6IEK7+fDbZNgDrXh4MCBvq1cx2
RbW8VTT869NQblytYnC6CC556OQ+lqdtu7P+dnSlsQQEt1v+Hvz/wHH8MrR+k0h6
3EMWEMirPGN/s8iJ4PzcawHadstpLHbgoOIN9mhs2avfBbfaZCU7j+IOE5i1dKkP
bCaHh0niiMNCqAnUCDl8zDEkSiSlO3XLfWBZnJnpfvBoxAjzAj7QK/ZRCOfJLp7k
S8RfY2exNe7KrGAqoOjbnJhQQge2vtI1BOGpTyha3Q/vBhEbxdFOtY5sWXRP7Xzt
gymNW4hXxoYPfBO/8++VmJ6CcKiX/XDfx3DeXuhyIL29SzFkEQMZnQHeOWCh6Tow
Lu/SesVDuW3gVk23aXVLq4htC/cjhz/MGWmO3RXTzuL7JGYX3vO79MTcAdRft/js
xnGhq7DQuH3qPERWylFl4iVwLqbPKj7vwWAr9vdwJdjouY8HUn/+vX/YZbbOeZrZ
F0BSqrS1SeE49+kxcNDNXEhgE4HzWcJ0odhlZPPHNUuHN3VFGvc0J8nx34WWVswe
0+IlKcp2XfYfop9Ohu74Gk0Sy2IgameEnlMGuT1/+IRpQpf56VC8HD3qaR03AG01
AJZCopOzDIqFe5/Tvgw4bBUsnBPO6pQ85yZtDotyEwCmpCIZrkek55HtUAL1oV7D
6pATnDT22by1fAZPAdKu2V4nMLrmc9g6iAZzTwuuTHJAXIcUKCqnf2z/Of6TbexO
tt2krGUGDczkeQZRC9goBLMmYiUtCQWdeuxzm1JxP8VTpXpcPYvrxE9+n+wxWHYl
/MxpIG0D327dxnurQOQuQWwXWcvZmnv5rSXZ1zldG8lsYfmQWsIdw0YUvbHrRu6C
QQhsm+2OSKYJyBbysHNBAN55tF5nttmazlufRb2Ei/XmzSlHXbAQNh05JTYTIg3y
I8i/AlmQsh6/2cwcUMskswxkuGrYlZzLXZz00pgvGfcFas2ulXAgN86ZEvuY6FsC
l7zuzOymRMrPtPoFDeyJD5ixUGl2cYw62vf6Ggoi0vbxbeLbFDPLHlu2jhCLng0a
2RsACYMVq5bQirgSudWC72+5A9Nst1HYgo1q+DMeS0hzq1PI4Sn/HrknXTXMugHs
KCy5Xg9SMb1pQZulfHjw2bngToSRNvjWqUkCmFtFHgF3QLMw8yW/e7QexxVsMr1f
Ta1mM5LLiDmVTelQOfpy7haskfNqB5R+XUWWduGgGJqS/Fr+LLRleXLoKgwZ5RdA
lPhW1BufmBYtWRvxTzfp7/yh0f83tUeKZPRxeCa/ICT+mJ5t7axVa3xvknfVw4Uf
W9i43Dhpw7Cv2GEqcUAXpj1mS2SRnr7fAFoJ5QEF4jjNRSo3cRIcPEq6SczlF5Fy
YFf1vmLcL0radOnwwejppRshYvq1UenjrVECZo92vUC2X3xlzTLqcbC1F1JiOdUt
LbF3cLWg6ngf0g3lKxNK7hu1IeaZm0eZ9dytJdPFzvLfoO9WD8MJW+NQUiSPYGvS
NaD1axqecsC/EbvF726RbYu48FGNYPiUZpdw5IfpXqj+09Z1pKy5f3F3G90pr13s
uaegjX74ePqISBVLZxwvqKNtXdT9qeGFRgL650TvpTaZ8WZPJyQyqdhp5ON4S7VH
L3hbxyYgQJoVKOJ5U9K76QWSRWks2P6YIUGNmelpYn8UoXJMiU4oSWJyX/wWSXCQ
WH0vKpoKbfoid09gDHpiYZ44FBBF5EOaXwjPz+8PO7iiPsr6qQ6RRQesdXnilklI
OMTqR+KQyz8LSmky2oNk/fhI0CL7GxmdSoL4/i361r/Xim4+2zCIVOul5hsOWXhE
3uiwmQQKcK7xIxsVA55vZZSG3A89dGhQcdDFcQb+Xxrua7UrCDLdudI4RCW6d8TB
/5AnXo73P6Wkg0E9Sa+RxpExyPEa/t8LddmlXETBMVLNNT4dwF+A1CVsM+vEwk1N
eUcJoLtBvACfQnhrRx1DJ+cOJ3S8lYurtYAjbCFm72UDb3Vbs3vIt9+asDC9AVIb
XOvB+AHl2WAy9NNtcF1qvwIJaeNmmpolA7+l4Lc2bTk+y48EViu9QbFRJwQT2q7Q
AEsea3vhBnsCcW9yUHV4oj9Ur/cLg29qlw7EHIzqQhD4txTG9OJVoBxgWJj9S0Y/
8D+Ddjm1DOO40hExH3su5qm6cGwiCsrtqvQSJXOSki4iA5AWGhW7hxHYiRSmQLfP
d8RDYs02jO0Rv/a11t9nvWKDRg/db0479ywceuPcfwqu1o5oqWr784lOvK/xa/Eo
3aCqFya6ZdbJ418sPngx42KPZGi/VI+XWbRssRq2uLb2GVdDEiEoEVNoqTO3N77/
9Mt4uj4rnfG4VIrL1xEiVPkttQuKSOhCZYd83chisPc71H9CWKFEI31ZPaaGxF0x
DuDc5rmTBy+U4phHNkQnWpfXKlQlRMybZQ4ffpwj7PQOUjjpwZ4MCmbnFx3xpnQS
2MzGg6sduPF9c3WJbT9nPKq0v9Z55rsIJ0Kz/qaPVH3jfcJ0yAzZ+/oWJVLN980n
MBG0cQR6SKJBi4EJAfntGd9ccnQjjGnnwd1b78F48gssNwbtyJbysmwnffL7xuKP
egNg6Rt6ekwAc7vlf0MtnnsqRXPRh/Pe/dIBHJ4mLhC6YBkZ+JvQMi1WXRPUO1OW
Kfn+Xk3JkA2/5gc9F13ulOKOEUhSxu5H6qbwlb31XOSjIh7R3F+oYTMx4iMvcgkH
6DzJtfsZ32TboJqrV+++QYo/HKRTfuFbhBDv0bOQTVvCko8EysXIoFt9fMH/i6nT
tPOcKDh06e8wtrgF+X9Z4E/JglGhJZmmQxPy7cRrbKxuC76AyoxPTQIlX30Vh6p1
vylkJxQIxa5QyqmadZxcMnUTbmUiIxniXA8V7gXI2RKpBrsYKnM1xEE+DKYhDjT+
vlFyBCzPbl0WVAWS4zx4uosgyzjpunJqb+yKaS8LQJVkpREENhnKXvx9WjzzYQfM
V6wdw0rUmroug09boDmJcOEYcxpMepNBEtXHRoRPvSZGUrYMIxNM4A9blerARuHm
IcQAiEUE+YoNz/GLlS/TJ392I4jfiJ/vhUVWHWmZRuhpsjGymI7NZ1409SXELrNN
wcCQ+fWR6zoT4I+K/shccF63y+cXonWLZx3A4Zu0U+Cwji2N4yy4sxfey4hXZVH3
8DXqBXWA+S6fsdP6w44hMqGIwfmSRU0K9XmlzS5yBP+BnRafxtyav7hl/0wWFLQh
bbcUcyECm/KuHf+imjg6X+1Gpm9wRRpI0wBGF4jBVi5DprsdhobOFGcmSr6ihmvS
i0Row1qhIGeLb50lI9Vndow9/rrH6dYWdKHjptBCSY39sttkvsia7lUtM1+rLtNH
7Dq8Qt69Mnl+l63EXWEg4f1V3c/+1gErWXWzwawQEaBeIpeXlX1EAQFfExPtocnA
XLEuWQVp/mUywFjuihVGNcPDN+rS9CB44zIOUTrT8/kuqV8Q2sRHrNOcY7TmR4OW
ktQunqgE8Z9ff7ylZ10blj0qOcmAW5Rx81+DgmvmvjPI8RHsnqESrayzEt8yP+Q/
Pto58fnmDGgsircobM4RaEXAsvXP3tRTa9qa+rm91VPgCjrYh0Ok54MyUsctauoQ
cYJldZLORWONuzwPvvil8uXDR4S9QPySWVQqfRiHqC3gskhBYHysyHktg12r2OpN
vBfhFUhh5ipgVIPyz1ZwP7PDxH/1mATbPQMLEdEuL2bN3s99jnKxtKnl3jxNTw5T
msFTZlSSMY3USNpwigGsGCrrU67lIBcuO7xSOtvP5nRslrIlCSfo9ncgH+8cRkcM
ra0k37aJJINH/lwfK7G9TwmqxYMrpd2SG7jW/0UzHeqZIZK2dhPcYv24YRPFFpOL
p2+uqVvc/xKrT2iZVLJl4/MaFHVsp+Fi59hJC2SxGlAJRrxIxmVmhYMgkkZud6eu
i1tW5VjKgRh9IZAOgxNGcn9oFgd5g48TjoNwUmEqD/OoPIpowFb1rq26F2oBKPlM
RCQK2bzV0QI38wO8WYPlsDzKaaCBatX8HBhNGsUuA+z+R3B+8HAQgtG9ZvWCu+Ip
s9xyh81olUgs95vjQ4ISLqPDOAr6WNdrjbxZ0D3RkFngtUS31tJmShbOf99hP4uf
St7EHnW6XX4uVOtKJw2WCP4PtyMZN+hffLA6mTZArMrwfrPj012Zt+vU2Fm/BBpr
yLD1yCEXDg7aYX2iHPjp7WrUWTkYUCBQf67GWWnpVEabliNix20hf+T0LEQTNrgi
nb93n+5mjg4RaKXyJpZ6Bxm45D6noglPstwTX2XMNbiCnd+hNcXJbXW+Iw6TsO3I
LB6iGdBfU99dJfdSvY0kcTflqxMUavvWCfQdKFfB2y+G9YlYAC/zv/puX1UazOAO
J/LYaTqeSTwfA1uZawv4Uwp5Ws35tUR3mrU8CSDGWZW3n2cjz6rtVQoPVmfDVThw
cwMBLclkFpnjYZ07saMsjfV0KiJDAzWJ00C8seMlAPyTHBl9ctwbIeq6NJMVaBEm
g1YBp6a+IGzoCyNS/ZmLHeXjYQ7blMMGit1VgQsMVCG88Z1/UUMDzYHVKn+JIzd4
MWM5JKS01KxkHHkGE9JzOzk0tsEAZzZ/QbzjSbIIza1EjRxA+900YssvpPKKEwTj
R22BrTdsEyOTzyoHM1kS+YJgd1k/B/gYuvY9OyeGfRBfyOhwnwnAhYkQPH+WUQKR
VweKVt9kWSQ4DBGahaNa4BUcd3NJ5ftZYYhTnMqfqoHJCBpJCCo4NNXYuOKhDPXa
QdTF70mX2zJNyyUKiiIxW5OiOKKNoTD1BujVRQq/PCbqE4TnJGmzCii3zy4UzzWo
waL4egqLJ3eFWRuOIqQfQ9eSzo+d8EbBhMDbrVktndLvmvrFqmtjwDt1mhZkCnTz
7XQpTiHdQmdALC3dFEaOj3ZQ6jhGQEhHJNjgv5kFFopVWsBIHdMcdXd6Ducheals
ghZdINXTmjGGI7SgPBBbiUSCztQ4NcnaSJR8oQDrjkZIYtm7rjdPN9aJKoNmptq0
zsVFygVO/nRQZx+14KyJPQ5GpFE8gBeTefevuipzf06cv6WRtd8QaC/wr4Gq+mZ8
eDqdHb8UTEoIlIP7xnzmS8J5Rp9bY5IYfoPwmt+Tn731O82nzwYh97bJ2MxG6K8j
7Qp+sFVFNemuZxtadgVO/Kv/jsFTJ3MLYMo4BPBf965AYybaHWXhRFuR7r2ZO483
gfp07oyHX8t1k0E7jxn5mVIQD8L8MpVgJrZ9GPF2wjegXTHp/Li5vHlgHfgfDz3G
A/MzmaXKPkfKLqhtqUFQBP7DLj62ACx7QJa3GJJ36r9PLMCg+73oTXEjIV4/lmIU
AOiDosKyNpZHb0GGyF+phwqD81/bojjmcjY5MuwHm64vn1XSom7FgO9G1DG2bJMI
+5XOwPwJPVW5UbGHRI+SInP4OOVBRNXdm8c1Wxdv6tduuqmHPLtD3wIJDq31d4gh
83MK7gsH0Vn5v0awsZFiuyVdkCDd8cJChuNxgXbukxOsaku2ZWvzmaQ/zJQTfI6v
2jGo/TuOMLsY1v2ck4tcLNbVxXaoes0EbvK2cZdYeNoELlUh5IAe2QeDtzLRDd1g
PiCaj0XOXD4MN1MzdZwoGgTVwcygbMoy77xwQhtvzvz/yI8I8/uCVy54t+bdGBcO
5iWuG6Ox1kTaPDlm43ZLXtuLFjc86gOBHJvcM8BkP150b7ZN9G/4wFwwYDnF5rEi
NE7Oou3WhmMLc0zBct4v6GuzC0fM3VTzhJDgrre5TEPJrRNL7ChqdtN4Ined50W8
G6rxTlEwgCY0de5bb5dQOiB52DbTZnuXGlAsDGwQrqZEsuA3uIX6TpZm9EOrgtbm
9fwSeLf+kqyrAwJ3jemx4jutpC1b6hLaOJrPZbhrP7HgOc8jOMiZpmLEpBvMjkPS
+eVXBq5u3eQKDbTxJSSWribvLx0suQrrD6ATyNv91CHqIyNcP+O0vJLlKB2kGiPv
Vb+VNp/s7eaOd/P/+HRUxu/hyki+WOf20lRNiGqpFe/H3UYcXAe2GBiMmhph8ijj
l1Tq/7gzWj0D4nfN04EBL+Ff/37bCrrcNZTIeNUQkPdaAWBET4Va7epJjFs4a7RM
Sy2WwM9o0OpOSzkqK8hfz3TROYfKpuRX8mu+0SnEa1I8cG7GQhsRhT+sLErJY7O0
cdGgDa9HmxBEZD2NQjPsKC7ZY7IhaUuh3/+5YBEYkGvDwfmTRQxV+QxT7wr6LIdw
J0y/oCSDBDwe431jZvJTbca+K5GFiQkY6umtfhRuBAuA9UMBtwoa63/++gJrJVW6
87tY1AKkhxf1+3hRqn5bJrkWQCPp8s7mjOtT6Oc8o9qh+1ufWKagsc8gyWXTTt5S
R4Ly8/ZjffWLzt+lFdHN6NCdLUZ8pcyAViYryH9GGTJWvLup3XfZ3YYl4HoFrHL+
KF4SGB0hWa+Low2hgkgRTvIXcLlf9f4IkVnOwNoUIKapgZ7vhK01Zk8daVo7VM0/
/ToerMh+SLYS6tL/00Co1nae1TnH9hUed4tUO5budN0+1iukF8b34BRbIpvY4sbW
IEJnmv6bOoIMcXaF7o/lx2CWpOVh/HmIs7oB13uy/POm3PzHKQ1mr7litwQ7Y0ww
0nn+oP1m6+fK2nmkrCM5F/F4KQRGuB7Vws4XZ+1qommmE2Z2lG4r+nNi7YW+UmR7
kq2JUZvnqaFdCwj00kCrSViID14/SlDt+vatkqjspLUCmcRKIy15tRNzmXEDz5N3
P4RHLWJ3Vv9aMd4/6EpolToofsSxsNiELr1YmWjwRzUENPcEIPo1uC/Suqm/FHym
JkdwHHzr0yZY2BMyMykSkhYvfsSsDYDXHZd/MbapeJo6HJh3/obXiSEigyftaFkZ
hW8+ebgQYByYvoMv0rRdb5C6cG8ES5sj0zzZCfY1+TFbJRVfE0Il+D9kUKiV6/lI
WV8r/C7WRqW5P1ZacpSlPkXGw0trKrYa+/+IXRvHaejrx6LPsGD2tP7eHnR0kMOv
ZcYZA8NFbcuLpkGSGrj2HyBL/fBcUJ1B9IUKyPq8VsrdB2QWc/Tj4XXzsT9+H1aD
UL0lotKiB8/WOVIzEO1YHE8QEmsj2Fla+MHjP7aST+ZYuImYXdrruv7X4G3V/UOO
kBEQT6lI+Gb7FZDxsc4Bl/2BqmM4CnSv0JGnlJmdJBE8P4HnU//XzwNg1Mn0a8YM
p7DAxRD6a9N+hPzy8zE4bEixA91Q7iYALA50WWek4GVH4MGPY+U12fXeZ++pfSw0
tdUDDG4xZSdlRFHY9j+TQ31kc4h+MdtOlGQAuXITfl43XbPAKiCTIedK23ON5+Ar
nx7jvxELoWKfZOLwCxNgGRyX3FpK0hnkGQMubnpXRl09+b/h7+SXvDrrG1CQHC24
PsKsF7RUkFvuc47yk/vjNi5yCcPt7bdvrBOS9qxvMLnGgmrCv29F1FblqyUksTOo
m+WmRzzHUoev6zg726mU1S3Z5B2kL2H8hMw6HDQOKzAPn3ecwBNbf0uqBDRO7hlP
xb9/lgLLHQqZcj+60ze4Ro74TAsnMQUQFIFmpLoEtTjJzVUJxFnHyqEQkWNOPhK3
N7lqjzUFEsLkOcGHVGn5GASTuvVuar9GXUNv1BG4rEPUy8D0tLthTlBv6D9FIwqf
KoSfq3rZk+Yrhz9L9Xy6dhfbRBwnL719Q9C6VVeNvNC+oHtCbqRaHAWKznQ8wkT/
kUEMGfh+sxcQafsUQw/lst+8cgcKscfoSX/PF7Z7jfX0l44LOePt8qXsd28Vw5i6
uMFe8N3XxHVajPAxm5UXWRL8tTH1YAdWTux4HExGhm5UY9Lnpq2EW/fLxSKW4H3x
4R0GKvWDSLID0URJBNw8lj307FAA3/qZQxarCQsUcWb8opBThbold1pCrIcXdNer
WhWAvUOseccHRd0506SXmZbe2e9wWQY/+duLJdCz/mIZ0O2nIsRUC1I/BYhFiLNB
E+y+6oeMeESIVTi5iaYx9ekbLQKyqGhGDpz49OqpZeRlFz9qXVx2dDlYnbMJd21L
LPKFDV2SgdWv6ZgDbLhaMDrsJxWkkhs+ohGJkmniNpNjDy0JlxIbZL3sJNjTPTJs
UVVkh8toVFKzt2LiLdVBdAXrALIFen2VoCPBJHpO0Gze0Nruv1Nt053uXf8t+Va1
0ZyTdRC5cA2rxiaOsU9HWkjnlWSGqxIGxBSCxeVAEXutZA8LX1fHfooO9Kjar62c
C7LC2ab7hg3bTQhVo196dS+OEUGblHqUoy8bMt3rI4PYVv9D/82rK4WaSrprwaYv
rNwSNynVsePnQ5XQhZ6aCcDEtKCoZnpcZfqFjQP7AyCBupuV8BrlMA+Tx4ducg21
Gc9zxzk6TV1xQrTfBJWEeUUC9uoVNVdWJX3MjN+paYB7DzZ8LIs9oPEXGl2Y39/O
wIvSzTugq5tjzxKX9YMuJiLcKgYaxkluAcwTzyDVfGj25824X8I9tDgOmfuDJckD
fUYOyDs7p11BsDfDnSlMxeRHJ0pHUiXHwyxBk6BN5CoOVUtE3jCvFc4vdN6uLfPb
8uPNMNczG1+1WJ6RpMUrXHN62wW1ElIEN6zvszYGf00QkUhJa8JNEBuYtg7akRTR
KIkTujB+lY68u8qjks0ZMXGEoTGcksbUmXcNft+LeBUudYkvUSK+YdPmTM8HUUBO
X0yEg5z95xCXzoWBpfGDWTDQMJn22ZbQRsghqUWc8cSWqv1vZsp3ftJv3CsdZu8c
P4BQ+amfbrsu4FqNjMK7W+5qKZoKYHK7M1mgwIXsgvOTfF4czbPoso9YXIZiJZho
HHVH+k5oVnnLgItEiqPw1b48DSpvdnyjxfckN++LUxiKEjzM+bzC0HkRlZPMBT1+
itNkBr9XO1Sa9mWuVABvOrKsQ/xR5pu9G1WJ2aiPpyWq0jfdBfizDDK3cgXuKb1p
QNGNLzKCCS81uBfapst7EO/O4IwQ2dbQceYun5aLtP69gtpVKxQZGlW/bHJ3GO+E
p6pkCgIQgMPKj3ao0a9PAelhyfekrB+86dNN4ImuMD3VTqgvpgQYx+EJBfCJskcJ
Yyqchcy18N/yYBSjTytWtnuHwzDmIdCyQamauFy94B0DBjdhcsQlUm+nSMamDHkw
oB3U43HODyoe4iFuvKCaOx4WtwkLgYssZEappy4raB7gUG7KxgVZl5C1BCcuEl21
N+IcfFXaobC2IRJwssgj6HoVVn8FdC5COeunDfsqgqxD40F7h155k1gwVhFvr5dL
CEXNtfQKEZODau5uPjLFkDVOeNiZq5mZDaBmxrPJQleFaVAyDk1GCR725ITgm+BH
ooCzYfdgCWQpUJulKzMRAc6M1K4cUHWGv9W6jYGgjhcqqcQaRGIZsVDoMj1ZQ397
HicU1/vyBfruo0JqwTNZY9ZOD6I8CkJ32JPI4A9lcdPXpZ3afFDQ79UpgcDimxa3
caxi/vliNbY3fxiiEhd7BXchBQhLgXtcFavdv8co0cFe+240sydNNBecj09o/bW6
2jux0UoTf7ghCMx1Mqd6OdIFQtWNHHtqWftDJVgBpRc05aKJmUjTzDUmH3BhHJWk
sdzveW9MokcVgB8ZV9P841gzI/lsa7lj6LIqvNGqgbRWa5XMeaizMEogho9GyQwB
fIcCO0BPCQfvQC+R0o8zcs0rFyxgbEryj6aV8sRrw7anc0jixZVs0bKltvuFhc0C
MLhOtu/wigW48+tkV1dRMbrOM5bm5EePc+91tjtYKE7Kq5y+HcD6O9PnJiKM0pEH
0s7HEnFoUfFrwJ4Lp8R/rGdyh3V36vWfohecnbhT/tEdMF+oQ9FfZvVfRg5M1YhR
69t8ABz1cnj4VFW0AHc+zwQyCvtlfcV7VGvg+190MgopSNs3+vkyWala4XB1dh02
wb0S1YOTTKhAdw7fveJBXcqgWK0qq+IoKGAuFltggf17Kg0NBJLmwv4TTmcXEENS
JvgFjn6EmyVTVXey4p3C6c4Dnpg2UiyCxZRc9RzoGVtWpwFvoc4ZZYgSE8FIjobS
nAEFoGTdsr82WGgMkAjKepdNUB2Hf8dbyvSf5EXqnH3WMbuCOXo0543hPVbOLDKC
tBzvdUBAw+epv3/6eo1VSRqs0TPBYAKKF2DvcD8jNEqbL8xU6X6if7uhw2VSKC0F
8eiztQS2rjN3VZDafHGYPMPmzRgrfdbZwi+q4ZBZeJ1Vvw9qTyLIkw9Ypu6uBXkH
TWzfJU4avp4xbU2aA+YehfPomFNf+9wqK6bEUPeGjX8CYE4C/UInknv6B5oIyswo
9qYR6vOA3qTdA0Z9XOB6pd5lIzKX+Xbt16Fx55OfYtwzAuwpVpuX2Fo1f3iuORkW
7+3STqCClaZ/BVljzoifYyyNrHAnvvFfT7shuepLnaA9eX/X7PaCGNuWkRLJaka6
ySsnoCf8NbGdENIw0GVuKUUFj1F1ufYO5Pda1Ktp2CTaYmExxxazL9OnLaMKNJBB
vbB+u2buoBgr8llNj8QH+nbU/KE9tbcLDJGys7r1be4zEsx64ITNZGQ6PBPnyfLu
fPGQd6RvtHxyuzlr0YFMsA4CqSbNlnNJldAb/VptK7gNkih+D4h/4N8B2FBTQVg/
8Pa+u6e/N2Fvtme9Mowg4h7vVUUJJX+JUSsV+LkXaYN4lQJ3OmyJdwXfY8KNvmEK
+iwhHn1jgAbYXBmy9SqOeqfz7yRITlrFSS7PYrd7gEvOEHNEX3+U5+kovrb8oSaY
jn4x7G0gVbr9sfrJMPyU2JFlLBJha2HD72Z9VsFHHUVpgLsJH4Zu1jVlTObUkD7J
viCjC+IpRgP9BOkqad0Vf2VxHHLFlaCF9tJk8VD4qvenCiNUQriI0Co1NpwskSXL
pjvCQ9J1UWaZ2CIJdW6jC1M5rg9pgtGvU+eGnvtty1XTPhK9ONGkmiQtnNqb10ZD
7/NHFspuyTvZZUHFBdd+jefO/1raIS/wPx56YlxQOq1EVg60JIE3MMZyofCkkoIl
d78nF0FsXjeJy09X5QYBueAT0Bj6jLzdCDClXZsYeqWuHrlRIrtfzMgEcXRSPswk
8AKkkby68c5JvbDabwacM4sdi2fa1EhcQSG7YiIJWuiZl6EEEkUv1C95eG9U8Dwq
z+0Db5QMLPyTkUFASk98aSXwtqIHqgVVesEy1uTxkxQ94NXyXHnOy+xSsTSC1LNX
Nd4+Hlx/F8HBMU+2cV3xWXOhu0HCmfJ+i7f+h4FY8qFxadqyLR3BvQe+n9/bNUVV
wD4DGban+1ZQWN30KWQtz6xiimUQhkLlX3w/QfJH+Yo8VlVkukp71EDWksSTWIjl
SSfUjL08IrY2zLDzRJxLqqixvKHDQcNo6V3/8xUZdXX6lVFYBRTSjlUAnjm+2hLu
q4Ne/pAg5b/BiAg97XCa9r1uElY6OOiTHVDOGokpZiqfsoDbrLbz7GDLLBM/wLF4
BFVFgNwBxpqzz/3aOfCxH2SCqSkbrpBEfvLIHHHkFpivDUzs8W5wqvfHCyMb427E
SreJFgz3LF3pY2rfQPA3CkIpjA/05HKEELPFL07DxPbQW8g6SjBljljKR2Lh6FLQ
KmnX+iK3UsJqw52DMDQQCHniEE8x3cy+yjXjbEFaidmFXWVZ25O31DF7CMFmfLJZ
s8kYmLjmF/IP4zzUcZbu2FM9+11vzzuCgG+GUsswX3D9i5tVsK25f8xAnwSjM+yO
SoXAJGQ4eZmfnhzjQjDGdrNxsjLN0JD0M973OI1GuCF2INStnr1vEy1sAoaigJN9
MZ+WOADQVMKdGCe5oVDVAlXEJdk4vJirG90Fke74qxjcoghrgRDKuslX7EFH+HZQ
hr8wjnMXMv3/mu6NODdE6gPxCKscpAzbLzp9pEIoJyihzwIFS/KP2NMnBgUYNeI5
/d6Jw8WkI3LgCQyriBSCOyT0t4801aPdgrbzxPs3t4/4EYK2Stbz0WdDb97sstSj
IaKWH3dcFpApiF+T2BsqX0X2zfXl+ZtWwFcPOXYBp4MTf8+paKlY+Ltyi/l0gQcH
s67RC3TILJwxx9fe108Jvm1z0v8Vg1LeJsdb8iO4Wr6iWh5699nD97n68iQyVgR0
hr4NN7mawVcQPKLaBaweSc36y3X/elkXysLYnB34Uab7BjuP3b9GSmqdtAhJKltv
rJsDrbT7SQqFWuw3NbnWCgrxfyC3S/Eo49Z38HqtsXqiWFdj4T+YhFoCE1H/HAIT
aXwa/mFj8bLMPuT58u2qVlItBPPWztnGxAKQq9WKo5OHEe1bs4/7ofwyki42ieoG
X0WzT30XBrZ9nOLyD1McZ9URvbpdD5tIzwBMieOxBuPEJ9SqlU7YHo4qE2v2BlZ3
bhdSu7O2zR8OXiJJH0FGSnlUaNR3tJtzdKQ2TA/GFciLKfbDxEm4hTDMh22237Yk
Qwouo2Or6Ws5llqxyTgmVJdcZX8eopr0XkwCNzXk8vodfzzpNT/27V/zzXbhWtTW
zKc5VaCKmP70KYs+pIkTZoCbbCacUiKnPVUY4YSTYzJtx4xv7OMeK5p918yjUlVT
wC+IVjLsiRU5Qe2veZKzJXNNuAAQqlzmtudIfeqB9u0KZF8J9UNI1gYnvNC1NGPJ
ZBm1QhgNCH7SaL0GdL6UH7S3/C/r5HshrF5dprcSp9rwXNSFckOB+G4hX78I7HEC
RV6u+AjEueQx8d490nAQp6NJukWgsHYBw1icUBRH9Uw=
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
7d1aayJWrMXzpB8QUg69LEGhkdg8kTVcSgErrhWC9h5ktvf28mB+Fzkz7OFSzaZs
80IyvnCzp+zC2zh8fwuHo4COAY6oRjnq/LP6i3+HDMDH54Poimqpv1cbnyOG/d8p
h7FEnApMTB0Na6uLXNCyFr+/j0RVPLBRnvBaJgy/IIdLIqplmbefsjGGV6h18FkB
8LcV/KXBQ6YigTcr+36rpFlgYqD3a5TOUXWPkd5uzGE3Vp2ho1T4C9FFaS0Gc9hU
v/z9pTs0tGrsLBTSpvyLQUtOKmYtT2PYoq5mL13dhf5c9O8Sbd6GtDp3MnSpFu1/
iPlP+DSDf4wZTrkhclS3eJBzDXz/FtSlL9ti2ZNdSOvQ/5OIMJoJ9wg21DWvRB7w
2glXJ3Qv5itZJgdpYCTYa+WwI5558A2aCMrmWqhMkPR+vNU+WvZAH/J+Z0Qm5/oZ
1xI3Dzme+JIOEnpdnDhpKL77zgixAO2m+8C+6YasAB9Z2OW1pUP8dfreah8I7XLz
bSQqyXrDR8H6Qvj9XpGJm4CzTcALDqK8f+5IMc+Pwe8WbmT2YCLPcOdd+w9z99TL
vKgv+6IYBwDnFUGWKkS9t9e81ESbHHIBJCwy+Bhi7OSZK03KrV4KmqXRTX/Oglrt
7MHih1HY/pAitWT2zBBNjaRDx8EfBrBT36IAe5sV22D00rtBUIR2HSu2FDa4e/DI
50Kg9bR0ZsHFx2qG57cA7qpYNF7zpr+46JOle6Hes/Sj0bRZFw3Lbs1/b4idkhJl
7PwwplxpMQMH8+RAMknJr6ZIIIZ8BJGa7BIN48NJbPS+E4owMmLXYAVW5ecUf+Zn
k8xUzXulfvboFX/T3d9UVA3/ahpabTbH4+91Zj0wjqIDSaJwfXvUc/1O1adsWfcl
NSFSjEA8WOSHjapxYwVcAYiTeV/fiY/5twNcGvLZ2UUPodGaATyHNr4tuH4YFA68
9SrTFTp2wffDTKVd3z5zS65IRdXY/U2U/9wqMih9PWLuZgFK0fIELEnjThhJAY9M
tge6ZWPFLqHmvQt3aOdclNbp2EvsuZ2teoduVMAY7GdVtxq4HxzRgkfsVlbZ8ffD
xMuMJtXwXxPkRwzAETL34hkl/cNcINhhFQJLbiASE+RtRAaxupsLAGz46uUk0ZXE
iFCRbanBiT37cHMeyJGIqkyGjT1jOvsDao84LK8bfjdNiUUz4C/r5K/b0lqHQ6I3
WKrZzLl6aRcTDLTNS33yx+DnBWC+roZ3n+Bu9GPD8ZI8tfAE86dpZTorlelstNpb
KVxeZ4fdace/rx6LLVmNz9r+J60MwJAiFdiQzbn3nwE+kPN02J+xjQLQ1JIysRUR
dFWrrZDAWhDCVKLe03/wpwXTGitKpwKlSE0BV12113uvwDNJz/ueTvJHq6gkzgZG
DEvRc2xOvmvcDi458mkIHcDoCN4JoXJVXUyPsVe2c9rWSnvDv/VACyKnIcfQ66fl
+4khvbRKSO0LleMP9ECFT9PDET+TqIfCQXi89ijYa1GNvpFPGAGxPAhJ7ZIJeQqx
twzF6G9gQsYhVb7If/O8MHpMvOWTe9fyFnhmgHvFzbHocHiOm0hkzt5i3PsokWt4
4SNeV/k+axGTmmnDm75OqOvPv2e2zGIpaPVnXMxeFQLjCmvWjoT1o0jGZtNJitXC
IpgH211ML9GbEFt6JMecQW1TmR+yjWq9Hkq20v4NB47Q7Rs3XUtGyYIlwWl7NKWI
X8d+y23eE9LvIu0fUtsWa9Tts7hAOrgOxWME5hKRw6PbK5fmVRC65tUMVXWdEoSt
GU6ndhOXbfd3rM3c2yYCM97gvHxA/OVfIhRVc2sbA/rxow0A+8wO7Xb+k7g+dl6M
ZW1GAouIFAMzQnzMaH61u0HDrT3o+S73bTOytzfnRRfgaT6mjlnkd/e1TMnSnDpG
1slbRdA66mSuN467uLNSXbRpdy3PHk7A2/XcQqAIeekHjJgPjblZBZy0r+r3K+0U
pJ9mTL0bsf7IC0XFHhWzSnmr23ZFa28MR9ww3M66io2vuqr2X1459FzlzpchUeVP
CJLDyvIFnYJcLjV/bZXM6Ps0MppHGiB7pcvmPomfPhwAdLb/XgYbrs+YpWM/KhfJ
pQrNjsdsi0liraU48WMhp895Y17lOtrbDGuWQTjbqNhE2YErwYpyywmy3lt4TQtO
dn+9qtrDgvDhFBTo+TWbb4pbTtFHNlQhsy8GY02/032hvW+xsx17mJ8xPqnjIbC7
o+EyroqDD50vKSx9VLrn77YatOfPiSnamJJoYYwzv5ZALnKrzPan1iJUmNqTeG21
/yNA/fTN0/8Ecq2M4vYXNl8c57JXOq4/I9R8jwF2DIQH/RNiRRlj67yReggJkeKD
7vnju2UaHWM/kAzAJzn1SFgSw32gBJF6GT90JU/owtWdRbKyolexx4H4IHTlXnnk
b0gl9/d4qtLwoFZYt3tPHBe+W4Y2D2z6i6UTyr7n7xgxfsjk5SZaMYG734Xpik2n
Z00WGBFc7ArTTWG/Lg05xngBLRF/aFWv//BrAusZ8SdVnffWS6MqaNNp0CiU5iEo
vnwaFtCPIORmWfv+1dbx4z4cEdxC4dQ86Gre+25XtpeS9SNQAlEFRPucUF2ns0Eu
K6GUQKWEyTjpejSgezGlsSWHToD4FVGKcUGGolHiFR9+GGuehEBvySmnxt+Bj8Mr
FsIzRX4PtLSRMlRdTLxbyOhjc5UapZF3Cy//0jNWNufdhLXZI64p17F9R5UDqGMw
tvsObbU+nKq0i0sT2btyW0EKdAMSMGmw1dkuSM04H09p04FjZ42VwB7H+Eu+2nGt
v2HEVXZobpxFRbC6RA/Bx/jyzz7bsBCA/c7wZ9QNbwMq0B1q4qxo6WKACkxTmr8x
q1XADKUM9KIzaXMgD26FEtC3vBNCjxmJBjhmZTvEUwo46rOhcJSCmpLXeyMs4tVx
o4Q2T9AtrDZyEDGFqBSw4p8EhUjIUDVTB9c+8TpBjrZwne6iq2nVQaqqdfbHnSzn
uFBTZWb7P5xJXMqB/EoWhRps2c74gjx0T6QrVHygtjJRmQidc/7w1/1AL5VH6nph
VyYYgM/NRxu2ynLOTTdoN7y/RKmR2eV+jQyQDhEjdo7wZa7eCMVoHoi/k6ftLS3D
cqZsDvg6lfZujHEWCr5i+ThoTYWMsy1SvZBRRPfHxOCwNLc926Kt+8UDfDQoY26M
iPiACsfqaNHI94Nb0jiFwUU9xZj3Y0armBFZuMHWlsFstcxddRVQq1njP2VC8L/r
O3hVyx3eCjk+HCMVSg4p/an6d2TZ+ViSL6ustkBKxvMFyVsCWSX4qWYaWda4dAbD
0ByH16mtsiUbTRmRU0vnciHPIDyODQHXRKugk1uk6T008clD5EOy+IOT9TEPaqTV
GqwcmBRE8/eTN927ktl6UpyKCq4EnYf8jr1bKrVWmzbSh0N3CinUcUgzlIUr7IqG
sLEtxeHr30FhV0YLuxPqlgr+jE9CJXhU8nODqGrs3ClBG1LVv5fbjI4k+gNxMBcc
5Jul2oDbWxsO4NZ4vSw4E0RKgoFRtSi1DC615ASUPZ8CISAfjy5eZBc+75uGREVV
sln5T3ig/EH6PdC91jDDsVVWLlSRTGEKyS1DInbNfzyB2c5IwZFdEMdtqPWrwa0m
VwNJdtCIjDMdVSZPKdn3dDFJGSnp316bLWsW4p6Xq9kWpI3dNTRXM4+vV5UqXBpQ
mph0qzx33wp50ISaXRb0KzP5pduV4Tfsu9RW4GN8/gs5z/EJMwlR3TAC9FHWDEQN
1LrI1LnDDhuILZwP2qwVHVkpeoCj+GdpwsRLJn7tdqnYeJeq2/9nZHRfPmZ303O1
AC4PbRqgAyo4BpYh/OhPXH+L0/Yz/qfnqMNz5kirWqUdtQ7nndiC6pRHjvKY2vm7
H+yuou9C6hx9FKE7DqY+BNeXzL/yiy7c2hPADfRZI+Gknpknhhya2T3T9RceeJlg
JY5JPFRqU6XhQVEUmYIyVsr7AqJv1LAKtdgcPb/Xz6ObAP53tdgO9aTk3mJt9sn8
8cqXm2Xmi1xObRVG+9tTfOmk1gPgkdMHVZXdRYX1pA03AXjEFZqUwLw0v1i2mzBW
edCq4N2B5ESwNmYvRxzNbNVjceC7Hf2T85UYRebN0e36bHC4+ZCEwF3zvmtz+yeO
xFoFMQ01usxzd29L7VYcr/3OAZ8GdPjdWfm3k6Zw4oh9mDbcN6t+39CtQ28hulPW
5z3Q68e31BNAuKMrJX7izOOQxV0RaO7+8m+AcsqGO0kd0/lyNH7C9Og2rX7PPI6D
x+H6OKPsB1TulHhZ2sHe0cDZMCKW3+VNPnMJ0T9IuA7XnUk+XDSJDIrUokouN4Gj
BOLGTngcUiJyaQ/DQc95aE3Zr5a+f1zw5JX9azXsTsu9nPM+lC7BiWgII9IQS7qm
JPan4t/iGT2QAH+u7PFcfaRrr2AMHfKOee5dKJg/4kpmgj4FPuAWaKi+kCxO8Q6A
/j0/yEluYJKDRCN3hYXRADit2iSfYF66TB44NhDo7dLlI58OoFf3Vi+/bVrD2LET
XUW4sT78qY9hA9I7Q4kxkNpyKZxzA5JzmY7KDZBk1DRiatVkY3+MhQdr/esG5zql
6QBz6GbzsNsCpTzZmGnOxeXLTNS8aW/4ZKUCj8UlsXE0qvHZvN+Kj96veJSMg/Rw
EbJT10b6bfNrtL4Sn7kxCJozvxwek8POwPBPAGvTtR6AqlmhYCL7or27AYdKJrAH
Tv8I4JLuxYCfcIfG9IoWeoCNlWnbMTznNfH8G2BpUk5UYCoyXbwR4whXf0yN9vVE
buAtUns+QsMQBrfZrB8P5Ed6kBFDRNMCssFQmTaB8GNZmJzZIDVYgfNnwtMIViAC
hgSGQ9GfLAU97LHSLJTnPiSH3sXd0768nahL9dXmSbGWJOu1XA8nj8nyrWFQce4W
MbKJ86hXqWXpeh5fvX/d/ZQlk2+9UPkDpQIRGeEZs0QXXAUaHwAv15v5/4l9OkmV
gyFEKsBSoFVn6miVO2bcQiNVI1ANfoULj7VqZJki3zL68p/mhz+yerBZbV4VOL2R
OigeNdbMlsZop7I67WFD+3u7+VcZTrgnn4CzZ4vJKe2Tn99A06T5GflJRgDrhUYt
Kfkzfgqo9D4zLMlaT1Gs5VMRbM9ku0zMGko1/gJ08JEFgB5Taq3BXWsGIE/XGQNe
qKQmELsdUeEfePT3t4QxEad01VAVSL9KwKuCbxgm/GtHjG/AqA/P8JZPhrtMyh94
xbs8mV/mHke1J97JYR7anygsl/J1XgyBmfQy5WgSMXoKTksQzgs1HbL/S2NPiwki
PyEDPkzT8p9yy5B82X/cyTjbLXteF+fu3T5r5RVAPOpuGC+Mavksz/Famyx9gnMH
s+9Cjf1BNrXofuob4Nv8qWWYa0cgxkUhB8DD5+KUhG8hSazxqdYzlRYyi+V7N7GI
6Zb7YsIg/OYRLxnOa2pvVoml2gvJBl/jnjd2maQn0BqAEU0yNk7xw1MFKY/mK3OC
F1XRJt1WiKSUxZYyj4QpnLsOodUUylhcu6dXrXQ5arbhU+zNUzkEkFbPWH8+09Tm
gckNgs12VcdfdkW8nAvWnBlKXDDoCtnmmIEY6HAoPO22xcA4OV1WNk2EDBmEESTL
i1C+T6AksrYwl+g8eBSnDkqjSz0OTiO84XhINUjPtkFQu+xUw7exKfgbwvvHPE3T
8b1HdchPzBCCCuh6ItCLk3bDNNLNMlMpDDlIt0Uvxg35Fe1gqyzA7zezx7pmXlqE
07k2Op7cEFGbUFKzyqlEMuSNvezLUI5ORkVszOXx4w07lsoJj5z8PDihDh73Ii92
mGAbKFFyXglLAr90THA3PALMT//z6vVaAkJKCrV1YrErp+P3Hp79GcUPuRS4Fq+H
RRMv3bzK7HNHIfZsioV4OcBCGHwW6oqqktpBs+DUhI9M7cem6gwB8xelcmm1oFTb
fkXnvkqavmMs/IycFnbbCRdqeHKjCQDoC1YMFOr58pMTfa0QLOKTJP0zHI1uFHXH
ge9/IS4IFscYy8VX30Vom60Wzr4V9L5q1wvir1yB/jT8PIQCB3HQ9sIHhlzKMusP
oQZlItIejNff+kVKoHFXGkZFmCL9wgMKQpERS7MchUrwkSg8aersJvUnzaRHzfrC
GvKCdhXCL7mEVI/t47LQi0ajv5LlHCvMkkjnZjQR3QvrTHFSEZXfnZZmPsmV9BFn
wyP2QMriydVtTtGq+QUxcKtSjsWcbS35qf/hRKALBd3XFVKzhpZcYmB/LyOvyUP1
pmFJ/U0BoxY7bLMD5nwkyAlPyqsYofo0aHuQLRbj1HPebyjeGZMgfwl4MwnjyF6k
p1BGNUjmHXUotIFw9j3mEYZveNd1PSE3Wg53Yo7+ipG3KzG+9sKLSsxD3Of02iPn
qbo6/w1Q8pI4zlctaKqnL7P36M2Ze7iIyTP0+7L/jMAXPprKao8PwDjtBMucIoOd
b9BqdnbrJ3S9/Y7yPoRPamCG4PyMD0R8S6KWGxSuVKr+VIZCsVZ4g5yf3NouHyVg
etOEazW11iprw7JfTPr8gn7kJjXp34TC7WLjbiLWiNrrLkE0b1SM3zKcCjIeBFNx
kAbycMf71PErH3y2sISGb8Jba8GD2G2ru7VKBnWoOpKDBRQWt1RkT/9OmfGiJD0/
FNFMSgb7w1KWNOnZi5PnAaB2S9WGU+z55/YMinLGDarIifg6sWxiq4AEkrUfn/pA
6ER6YJIXjzuU1XIaDh3KWEQPOpjd3kRHbcM68X5RdiTDFH1rJzZLbe8MXKd4GHZd
5viPRpTOL96blXtdef08vuqhd7yY5PVVkjIE5CkSFwy4vUIJZ8y2wkiRcQt2G/Lv
PNRXVpO58N3IzmLtxQSyamNVJx1b/bO2wxaefagwgwi72SCkqkZ4c5IuEwAR0F7o
2Y74UlOkrpRSXez9fezDDsaCpZTQpaf1H+pUJTFaNrNaW/QWZYc6bpcdXuIiFl4N
blZLM41AC+o9ZlRvDXcZjMh4UIwTmKkEDSF3bULTobqEQfVtniMwMKbp0g8k1vdW
LaAbsqRwr8nxqMtuqAShT3FSwqtN4+cG6SSazXrocSOWe5UpgT+OLVikNdU0fkpk
XOZwk7xxnnppvtsw9gCRBH5FOp78xnyc+bpwaoh1lMmfY1vvRHTJeorseP2ycaYY
00oZtTr/LWf1FN4V63ZFFWRuyK0elCqRPGi7h21kX3uelRauCxasaz/RKaYZImca
n4QwFAwUf8EWGkK4/HCteMNyBfh05/z6I+dUUdWeKSQ9CXNf1dxosqjTdN3/EZt+
Yc1rE1kQYl6XSyf3caSzYf0Ua8DAkjzBmcGNTXyqWpNxyCh1ty1A22ASU6jhs8fy
bP59p/9IBD6WtN115hcgOBKWUjqHrG7P3+QuCht+08YatZPH1y3/04QgRbp8xQMH
w/cIY5ZzDMNJJNu9ByA9WFeSiA0YZNDEclUfgMfqb0IP4/+EdcJaUgA2N/vyt9k+
9xNEaHLfupUbLMyzH8fefbF1J1MZsYxOscjkX7wPcv+68B81EAfJ2hRYZfwbFvf4
LtqmXgMlUPwQ5IoGCU5cGoWxpfiycRZ4F937gVLOo4eW4Sn+07L3LFOCBpF13kC7
JhKrt5annlgTMjz16DrTW3jUb3SwOf5bxUZ5+6AZh9TTtDitur+pX9SYBVEI8apD
LnHsrajYB9kiyTz4L0/0OMU61cjU/iGd78WAn/n3TmYWOSPUmamHoLrIdW+zMSZQ
ixgYSqqk1UINH3uB4mXRLkXI5OaLrwYJts10OmioTW6P9kPjHf6CfRImn0jFvLzL
+ktbFfe9Tt1cRLrTzkKLgGPq87FtiJIs3DmOprFsjH7HurPjq1brL+CSJV70qsHB
EbRCrJrL8ON+lB6nFCY4pqZC4eeXjFMtvzGJgcnN7injmd1IaN7iSaU+Qt/JU7eh
6ogvHRT8FIuuyus37LBYwupMG2rOIe1UH5stGzaKhr7Ud1XFNEE8sX3DJ//DpDsw
sj+6Y4yyJUSClmmW28fWRU7YCMoSDoeLz5BokiK6juN/pR+qYd87Ps/H+loVZIDX
uVSAilgmb8Qc1QdiWI8B3M1r7DoiZsjonRLD8TKxfTi3VYYu3zmSVaCzFJC099DC
vIiGEqz4QDxW0Jqx28s6DT+LqkSeqznnXtoEZDAI4Zjw1FCT5j6VlZoxmFkS0S2L
Zud92/3b1vIUjhvqcp6xtbsuXCNyOYuwEvJYMAZ5X09PNdnemmDLZ7LQ0VQim5nD
Ngpl4PJjxlGgTG5+3FS7r5xjQhBGqqe2dFLFzY1gwK/2SMAU8/CfSPTlbo0Pt0SN
X9Lf3eFOWa3xkoour/PLQKzYjUc9kNnZWGova/3YHKMgSu9oO3hlodelFShSTDHn
Zh1buM5pu1tju/qIlrpt10KoUqZHonmNSx8lURlnRaoy/3yD8tA8zmNIN37HwW0j
d1bc7RGEH2bqkUouMUhXZvFOWRXkpfPeEbbX4sdBssWqmteDnkf1fO3n/5u+qOSm
kqZMDyNtxBVPNxcaLzmarNnx45R2AoGJ1P2YkvTYNXb93UB1/1eCcOHE0SwnF5Ds
iNemwr7RvkaLAgtdw2jZAXYGMmTdtYkHeW68P2D/3G4/UQAR6SNorM9es5v0QDdY
sPj7EIu8YZcdE3bhyi2Zb0h3uFx39fR+UAvZbVxj95NUnRsh49++p3eXogUYkdma
M2idLbCR8juVm9C/HARPDmJXriRizRKhFMRev9nyeALL49OBkm9Np55YmCkUNKHq
FPMB3XGXIrOwbp7j4bRs2Dpv16SXtV+Ft09pWmd5lox8OK1jtNJ/cXtGxqvXCkv4
8fEwaU8WWnDV2Xc9s38I04pMcFK27fwu+i8oqdnieA7Ftcva/EebE1pohomFbhCu
8d07FdA74Tt4+R0qzIz/+04hwN+wqlhgAqWJYbT3u2cl+ko5p2XUoWq7YsBhz/8S
syltBMox3NnGHWozY7DeW8Uf3nvCxHtYqh4izVVr5jzRdGJx5kF2rjA5q8RuhVfd
6PnW133uSzEei9jre+Gzt9L+Ozz5xYPTI59RUOkpe/111pX1neL8BjD1N+kol5gR
aTYKeHwtUrF4u8kDk1JHL6umDBGELToi4tQ6xq1r32PK+zia03r2/u4xixIOhcTW
YojNKt+xlrr3bH7PpT96eZ6dmXyc7VAwUqufHjV1X9U1hKqw5FqPs7prbTrYUZDx
urtVIkxbq4m2OafQxraju7XV0NEN2qDT1zaJ4Elypwbc9FIRKP0ybsqfEpSPV3Li
rr/XFp75+f6zsjVBNtVxYUr+/rCkKjSeyup7fvBkh7PMte4j19qHW9uoozCZEBm1
FBm39nHrbreZ536voudB+AO+u7sGVIeO63GwOzr0Awv6z0dIMHubX6iu4Og1rzKS
U9rzE2NjQz9uh2PsjtvsPSMul6ecf2557PbIWcIPurQxnHJcyWuZB8xL7sy9UiEI
mLPaARqKyvBonZwB7v9/Ryq0EJU/TojzxRxPW9K5I3/r1Lisck6T01GbqgYzK/Xc
3R8TKF/Ttbu9dnsV42+T8DIlbcXRtEX3gBOt3JtQ7js9UH4q3GJBsqhp3Y2Qi2y+
1TTtwBQxUtRVoPsDNOaOQhRsMktA6tzxtrcIBmD4KMh19kmEO9twSNN6ziV1nUvN
K9iYxxc7KYbj8frhxLQsxcsyCn+qfyu+6w7tS5KYMZHdn47U0yhbFKS9vMao5RSo
NZDKnH5DZmWY7aDQrvQY5auMmNZNCoLWplo1vRWKvZNvUdD1SF6tmvTwNMP4IE96
6CjvjHB2opzw0M83a0m1PgwvdgSDw9MHXoJK5drHadhMzT2N2e3weItv8yWupVTi
oAUVogtP2F2sjD2wn447XN+sU542iF6Nq+W+NYgPv4I/nBQsWI60BFYdgGNqz22G
30y17SCCEwsE9mZ0QfVjZx2BudUpFHebQUnRQWZxMdNt1nI9xYWQd7hhXHKQbrd9
ubXeQnMGrWpq98EW9pVLayP3bJmJWAsbBSNgQsnGeufkyCH9StMYKaotkb8Gzmrh
AYB+eAIRydd64GI4rJ+ONKx0K7qmo6csgWo3CjnsokrSy1Zk9ykGeVNjlFtxLDAl
RcS+aRP8Uo3iXp6pVLdFviSd0JSdcQUOgPMXYxQ/ms+vMcO1ZDnmJoEftGBdegWi
q12KKnbA4VZ1ndjunFBEYA+QMz0YmIEJ5EHL7lyMBHQB+mwNYDIqsnMtMADVbYx+
zd2toLCTHWWy5Q/zs8YK4ala573nA1yvB2OXttmqzbqlby0XDX1JUMsQuNOEsPx6
kGyR0I33JIABb1xkgZPjvanzM16r9P8/PYfwfV6iVifrKKWGkNkEIUNouHTStM8E
a+E4FcQWid69XIEVMz5mm+Es3+OSJwBAKca5seI8P52MUZeHRRnH2RJZhbuxwsi0
KWsLHB1AWwOUOLFLPKM8caIdgBOuoUmPh8PLSM1UpWJnx31xkWcHAEv/QUDChSR4
QFhaLynvjVfKzAncOZzsr4WsByE0GWFdfqSsc+Hs6DA5PemmUpScTMtwPa9PQflF
2Ofg/7Ot0iTHwJikgzpDVBtSqZOKONc2QVnCiOrab3/cq6pKwHH59vTdKH7aDytK
OaEyfur9A8n9WZZ0pm/wAbS2ePXLgL28Dcu6JeXQVBebmfdlUfY2XN5rX5F+2GTa
PsvGZEuE+FPxT29KaZaIIGPhBBefwGKwb492UZBNu3+8xT/bckKTu40osHOhTy4z
Wu9Z8z45UYeApF5gE9jak9NWXAeyCebrLWHnQHKKl9hUwfAgXSVOizVA3UNih9iY
mFFbx7Da0Y2n2ufpkgpdpS4xduglVUQvfUryRqi/gZu8n5DC+7MDD7kPxSM1nKY5
9ju0Ef6JwQMCzBku2zbhbB0hRwRpHEfTJ7sPNsWIp7Pmjt410smx/oiOJ3c+UhFp
7bzu5dRagtVwy7b/BlVZSJvk8AV6ILt2M+DocfK52g7rOC8O3aJVMeq8eF5e0IaC
2tIXCv5vsaYEzrQT7b+KkX8IlSBEyuiH/x+Wh4dn82hxa/SIu0MBwxlaNfF8D69P
oi1IYATmU5E5pcRlhCezTXIWFxS6XrCJsyRj0paQXtWAQPI6ttWw9VBkTm06lzfn
1kuvDSqqQpw8pnFwRcQR+aWDP6o4+Sp7Mpycm5spVoWW0Ad1Rks+06G2463P+eNm
becTWsNEpT8ZBCexoCBBuKlhJn35ijDjs5E42fit+mhBPRXqBmo1t7O1qHsG3MiB
M6pmSp2+52+8toN1ijK5U6fKeodwHnTIdR+mbwGQJQiceEcNwOPCPoqYykyHAEyZ
nMTPccDBuMME8+NdLHKULC5P8tBBiNQXPKt8GJPogh3dqOa67IE90/fKB/QeiuCa
CW+Caf2yB4IZfKFG3YQw6wqYLNyG3Wyl7yZ8tNNh070fEwKmTUA9+VYTTt7iWxZa
TbS9R2uNJuVljqC7z0VF3+o3K1Ywc4Mg2QK5cA68lSazKGLLN24rdm9Q4PAJJNqm
iLTC6EAAPmZ/dfB2jjXTNMn0H+v+4O4LqH1/8I3WaJOqNjaDY8B1gnlmYQxJaC/I
bEQjIyeKfuITd3zUy2IiSz3B0IPMMNukTlf/VpZWF2WxN+tGbA2SyTkzymM6oLSM
S3TQduWBg2Srd9Am8yK3mnmpJcJvhsYuYJT/KJVME/Z52S4ddBd24lvuENGG/ZHI
hCbUmhDGI+aZqgTtnRrUgpndMQA68a+Aq23MHgP0HI4dKam/u9jZY+1tDSFJxCEV
nZs7XbNQ+tI3kWafPBsn/lT7E3VR1xnNVm3YPXNqnpVgw1O0wAjZ2yfRkxn+iS7S
fEX3Hu6U7czLTcX1n88EDdfHYyK9gd2Xto2iBlnbJpNrW9C0728rgPJx3eZ3hhD/
WacZCHgYlCylygdXuPM09I9f80WFxoRsWjCFsTexgHyTaZw+LadmMr2ob8VlgUnP
K2wMrBih486XyNLhxk71VH5UyCYzPd6pTKM7n18ngvHY1VZtOY82eIJXgt8pLaK9
4ATTlhGGE+eHajRBD9CMEidR/jvrIQqNqcnl1BLUg5Ei1tUKWD/mTZoZi79tRMVM
Uq0VoKFo/yoVKF9GCy/ZykkYNv2anEJ9Y3HOj2MXB/fKs4tffBm9vTsprjLzuW3r
IgJZvhkltPYduqk4YArednb0EFaVLRgDdSjgJEHh7BixUOyVwkhMtrUObDMOKWVO
pu2eEOLESg3ng/Bmer+nDLch+epo4i7MnqYqbHiFNVR9fcBGtsR/FgFu0hcgV2oE
q6js29BdENb+JC+z5p/yS93PSZSQVhVqMjhMlQztuH6jVaNtDCDQ3QfqqFmm89d4
lEq5ushyMP9ukm8tT2+wseeSkFvRt47Seg9iFsov0On04d2P7c5yO24a4e6qhtE1
0Z2Ap9JMfsvkvyJQ89gh/n/CbgQco6D7E0oD0HZIMdVp/EUHxfiAfsYVXvsIpy9m
HLEZjLg63hXbDNYnJm8Y4iNFPASmMpvnyTbxL5MHaVZX4wdLZs/s6lIpb+QjiEES
HpuPqcpu3HntZoPOaFWALCNqgZdSJR0ndEerJLQIhcQ7W9d+O0yansxyHztl1fIC
vFeV6geRXvWWFgCUQm7JCnLFI5p48JF0F2YcSafHHGgmhhGEsEVvubd2LecDMwll
dlo32fY3UJ/rgg5Sx63B8Y2sS3ar2V4ndp95M4xMkbgVqM/OhktQui3nJGYDcTAA
uCwjnyvTV2ZIOXV/Zje50UyGO2LdIZzIPelVNLRlkGlca6eaJeQ2sjM13g15jeFc
QmibEFAKpp5GzaR3X3liG/LNwG1jOZ88EketKauFbNhCcdNG8mEsic5kPtILOoTE
UHREiauIm3FdeIx9azPRHUBZmz8fyRuiNKKMM5lYoHTqQcHJtn/XgPC5x9V1tHFJ
3Gbsrx/RlyXl8wiPJTV4uyFWjNRQGpLwxWOK8fI0wgUJi9Rnea17UxteuYX0F9Es
TpdSdKbTlKj/+CYiCTQMlg1b6UHyL7Z0i6b2UTJUttvwDx4HxFGojbIkoJZW86sE
eU3KEc84O4uw5rNgfmbfF1s2+1o0JlZwK93OUa9Q2CNp+uxGcx6wBNVihlq5DvQF
6CRX1WFCP+Lzr8UY15WnCgh4pVz6bft2/LuaTWmS2e8TQ8xXVx1jNK74zROSdCpp
ZnFjie0Jjao7liuM5NFM1HpEb9qD8K2KCy34eCAD3w2cfgrTQAFlN8E45NyXnVKk
6o/l2R5fELJBANvgPHBOJqPVmK7z93CAjAlNpPdkQ4qqwXe+OpucmB9qUDQzaPH0
KmNKBBrv+bLxTNJbCC9HX+YWDmfNrhcDqDnNdslpRxN8Lc74EV0iivzg8LJWflcV
nuUphR5zUTZBuENvn16U/rIRLoTWxphCE3clx8ARySZZnNUW98FhByONk/qZcV6s
P6S4hAl3SRsac3kAeH7pLGHUtyTBG23/ak/zsibQFb7Tsg/B46CJ5Qy+BA9afvQ4
NYdtEgvz8jRWqZM9KUF3IPZAwWedUWkmZghksqbr2Dkfxcma1M9acyYFblq3WgRc
yyS75GT/ChWMAt8+2sWg2Jwyw5ke2AzyyRUk5+6DHv8ERQY+72H/lj5dJbtImiGJ
1fSXXk1D8luEwhOvmE2FFq2clgHvT81gsYQTTtDoyWtTk50PBXTAS7OQgjHwbhXc
BAD0zLNGn8C3KaU59uB91NNCpXBAD2/1wMxSaC0XZelM/kFu3Gkfj4udSCMXDIlw
b9HcSJ+4jeyxMaNTEqdLdhafOoR1G8eVSngzVs70I7lF7yPkPLTLcZCavGzkKMkY
kydH9szIKPyhbOsTP3vCLX9eEV0cEZjx9i8hODkduNTFp3YKQlIMUXPO/EedzDUs
M5yDAC3BsVYt6z0FCA7a+aX1UzRYQJtan3pQk9fFvAyPqs11dT0UUFzsyBncmX0q
9ucp9OCrfkPXbz46Y5Bv0W0Lbdc0pHpkIJ3jUMFVWE4UAV4N9YAHKo5NGts4E3PE
aaZIaWMd5bFEMv10C/Bf6NyLkDUqqY5Kskkul7rRzbyfKPyMaQ8N9vBrLXt19A2I
K5IWbgzDwVmrr34WmvtowAP1ciQpijjlzkQQwWWFAykEWFiq3DKH0xZw3gMdOSX0
BaY9ojmnPlqlAs2j+nQ6xbvEJu3Ru0DZ9uzw3u2/gzskD4JxuL6kFNgCLgbFMWtg
QSjMMq4ccNLIJKuS8AiGu6/03PImmbspinrnfj6pK65SVT3rXJFYog9FyEBWc6Wq
YipTONrX22nXiJlduHC+9bNd0kVYL0D7+uq2tUmy35RSmckE+fbmGJoaDrooCyem
My1JFKvRi2tPxOyxFCv41ezK1xB57hq4RKM7UQ7E2hhzNJZhB/yuj5/RumBMUTNO
t+yDQV6mLiEWnnzPd6kb8yjHhiP0e2MNx8V/T+J86IxIxtpalvFuMXWLraquA7Yp
Hp5OmRL525CXYXGDNGLVxJVHZwizq3kwbVeAx5+wubidQPYGzrylsXI+zF7s+DBx
nAr9r8Znulf20x89ZVaa+jRNV2bkMs5M35zGPF/3f/jFaKrZnX6NX/7lUX7j8gE6
6+DZdGUC7MCd7276B4xxlloxZlEgPlp79tNrEcQqFp098uuUa1NsXwqITQlFrS3+
zb53cOKI357wXq0GUu8RJW2WYaMecVd3FN5otyDuGy/AMexc7IVRXhQZecz9OA6g
DA5toTb/+LvMUSJz6OuuLZYiGBHdg9vekrkIQnwWsFcAFxrnzVbqPcKkWCoBNddA
Se/EI8thJvKdI86g1DlXE23g8p6J13UiaBm0/yGaTieoG1DRgxasunveI+7RtGe1
WA+QYkLgIWshbSui9f6VP7TyoOXk0Wsxel922U+pVOmLaqnJZnO6+OH6D+MnXEAY
vnkv8Tr/EzHJfB7yUM+n4C7CdnckYEAU1+fMmh2C098LYNwWQfedw+JNIiOPaFj4
HqnLPLG/OtP1d18dnQEF5MWlxKbRM+DDHIt99O2r+NUquMT4ZfUQ5UdujDBbeK/C
CFVEy3X6HU4/MUfsEo1ImnDPPtWYmUundL0BXJpLK5ueMHZBp00+9l6Pc+2qIqXx
IVHxMWVELDEN6rKx4eMEzkBKfzjQzjRd8R9YgUeE4VWJDZHyJIUiE3souho7vRZc
f7KuhoSWtUwzZGBkiZgkPWH981+I1/NgVaNpq2SPxCAiSLWSA3iCZVaex8iIN9Gr
3CZBSiCNjfBBAMEUPbP/PqXx6XOUuV9B8kdWdW9mzuchtpRJUCYLjf+/GnC8+kay
sgGueIy9x8TmnLA7v23TBbTr5XiquFAEzClN9PYeGRcwLihVQpbfPNt8I+tYFYbb
Y+ciZbPqLUDdM689tREj+eckaMA8cli24a4DVPLVHAsV1gefy8j+nbxN8TxsPNcl
6aQW+sWRnwWPCDlw+YsS0MBH3vQ6HXOZ+4EA1krtfCZdiyuaAYYio9do6G4hDFvv
nQUjSxblSPgVjvh+0TUQiHn+PVPlQjyuz4mXdz9vQxO5SkIL9PX+ZMABJnwY9KnW
QGWM5mx6iqBLLC6P3SP3kH9ioelKx5aQFr22DbR2E76uNxIHxTbKw8iwN/z0ti+p
BO1nr5Q9RynJW2uw5CCafGuoW7F9q67YSM8nVtyj9ShaEjURId7VFS8oxv2+RI0p
SNQ+CGj9iKzKO+Q87hFP2slRxMf/YxDT9kLzQoIiu7cJeYMbSWEssRbgA2e0sunw
BRNJpCv2nWx42P3a/RVCLsPJQ07gqL62Lzq3WtUTM7zxuH91yBBDR3m9neIxFK75
vI5Dznwnaaq9aKFzBNF7ip5Mvm72rpM1cmTP2SDsrRqHTTfbAt+N2MRtHqCSs83v
Po4JDzK6LJSvTgG7B+28N+tU8fr1jCJ2+x/hzC2su2D67TYlZYJLpozZuJRcfi2i
4K6akMfapdNbUnjrIcnca2JRZ+uchn7PXNuB3sE0Js7ohG1fMVIevE2ijeV8Oejy
Wit7a+SwwshIS5s6nMT1c74nw15piI2cjEA539h70tROtPamzzaUlfDBxe3wcSqX
Y0/5XmCjSaxyugtKx+I5RBXjsyv6eOqtLtWlY1AloHZuGzAHtd4GmugQvxPCO/bv
BLBDH74YT7SqUzgBZMZqAfOvMg3e16z57Ax4htLJJVisib7rroOyDn5gVso4Szog
HZVySZ/ShzMfvZUSFxNAtOkqoM3KfAKZ9MB3UG3PMbo6KDPF2MHa9F//2PW38VFr
CvsT42Df65D0KkDoP27nmrKfyliD1MUwulJFRJiaC9B58lge93FBiqvW9682nhBH
jjPAdwEH8XyhhbzN6F1HQS9cMEqCYR2dVLwer+CsBBgRvC/KgtDc0LQwCB6L72hT
f/wvOSgircFj6ebjwNN2daHFQbGjME35LEHQJwJ4MIb3bLMmkKMXNpSzjqExUZcw
66gZzQtzv4x7PBFafg/1ge4vaTQNGh2iNcJEPaYucKgR+KfB0p/snnnBfnUbjxCx
s5Kw88oo26Pyk+3cQlJkSIbqHaw7OKASfrQ3PDKICVg5vjQ1959uFdKzCYvder2O
uv1vBVaVV9Hdd8Dz2OpBSKgtLOXFEKO6AItSX8WdldC6b5ip22bh3JOjAbd2JotK
R9LYI6B22EHsOaoN8Dvif8AuBPARKPSKthcz9KmmLkRLs6BZ9bB0OjE2dGpzKt/o
h6bN8vppXoOwU61v5rdMPkD7PZ6altBvnuZ1YrIbb1v4pA6845NZGaTePJVdoVG9
NZm0EU9xRjycVZTebgcUkAAE8/Z0p1OfDlrSYol4Fl6I5XVJe0eD/h/wukiNA3ko
wbY7APKpwX25LYO+0CPH/++WgvmBQaPEINuN8gccGrr9UkvQ3SCB9tk5p6Wwgb4V
qQxzmuKe+P6q/ZV2xXH1SApLNA973FuXqOmpScTubapJe7zZ6RzyP8pTsHBu2+gI
4PiUe19dmCooy0XdJoLOXXZsXCX4UkH0dA54T7dC4w434twwoMSDdbb43vggSkQe
CmQEUcsZRvrDBYNPv8VFyQCkKJPM6iLpb7CpQZXPziuVy7L4j2Hnif8BfPGDqrxs
gc+/Hu0d6hadn0gA0v2R6xnz/PD1rnLoqUysHT3x78OW8Pwav5qH2K1AzsjExnWl
PCBv+ha1gdBTG005MOMin1HIAZy8V6v3LumsfTKIWV0yqk/yBOVdeYl21GwKNYIL
AjAIvUSIy3BDSuTd/ZC7QkXU/jXk8LaRuFOH3Y1eOCvlspnWZ6aedgyH8xqwkDz6
Y0VNEADUqvvNyoKFCGIGDpKH6a/7F/nwnENliExiR0/bSqUqPq8qagwlH4Z6tPBv
bPFL/+2auOhuhI9dyK5Xgi1kAc2pZZ6EtRSxKAiKwKS7DS2TnEHHsA0sJPeJYCaH
jL2O19pTuUbIozjv4pPo0RYEkvkIfTIwse57/K2e/6GnNZ6nt5rldVLHaPFru3Pr
oCZz9Zq8pSI//UH2d1KT5nhgRVcqTY5FGZHHfMcitLB7sAvmGe4A71UAKiH58oI5
AqEIEdU7O3hyaIKreeQEJCPzY8CVSQ2L16yJjsdE5giMFjweMhY+I7ueLjgXD35h
f6oIc3FbA+PIQDSoOyQCbyT46wV/QRJrHQ4txneLY0xj3V0adApbUlstAoDcsYxI
wYGZdRMYNibeupcTUtFGbck0c/nO8tiUmFX9RCcEUQjyY6JBmPTY1JkB2VshSNwc
g+UAF167wwRpLnTahfa43dyM8QqxgfF2iawnjHNx2u3jV9ykJxtD7H2vY57dru51
+RPT6NU4u72lSZMoQJ5Vo8jR5UxXRU0bcOwwbo2fWQL6rJBfduToNkECnKUuico6
JvgRQT9yyRHI5HjsB2eHQPnug2jk1U6Mbp15nLt4R9Zk+oTdqD3mC/XlTgxyXjrk
faQpTf7gZ9bxQpPpGJhKTEZZ/NB2ktsp1brkARLFkZldvCfU0lqtruRMJj5tDjin
nt3GRnL6td/qNRuit9WUVK4mM/KmIVEbo2h3hnqaPzLrTvZGLtmxwq7jUvnlVE7k
/Fgn2niC8kVA/0rkDNzPqjQRbvSR8JaOHtA3Qp1AsIyic6pjKL3ZfZqpT7vITxSE
3RfzKReIjE2TRb/2M7t3IVZVBcS8yp1p8UP4V0ZFy5HGkv0aUqDiaV+2Gxe82LpS
qMtJ2b//akdHt+4pqIMmlPYFkN8AhEuIsVBLLz8A5kVFuJl+6E8LcxVrZX0ZxQ5I
Gr4A+jJ9Yy8OPaumwYGsVA0cnJnFBSTzuO0+d8nW92w7VYmE7xHiSGPbcdx6LiEa
MaIJVmf6NBi2eTWz0MgvXUPfY2+qGSbKdaJsdx/6mGkGswqWGXQZmN0oWTO1hvJh
Z3Vot3QeAotIIVRhG2cZySd0B2SUeAGDBPjLFtuYywn+Kpa1lsmhemSANet0OpVf
ucfqmha/m13gMBgV6crXVNVUEw1nSLs2b2hJXyDvNTBkrU84nRWu0uWAYTQO4nPS
F3+tZqkRtl0R4NG8ADknGw5A7mDVknpbpZitcd+ZirDpn0cseUCcJ57gpKvo+I+l
ghce6MqTs4oLqG6lPe3z5ZTxzoVVMdb9G7zedZ6qXU6MUEnDsulPOTyZrO8O9+X5
UYHIJ5ya3doLAQMSKsEYoU1jF5YMe2coIEJKxJRNiFfAZsgenpUsTyTK3Z2YnXP8
h8Aeu5qnFXwdlWDd8IkQvrb9oYBnZNQao3a3CmNGBqL8GlULVvA79spoKqvVbdX8
vK4yz8WmO65DFQ9+s14PTeFZB2DWVdZJ5C4QYUectiZ+Q3qDaotNxV0YyF5+qMUd
ELuiHzQmTMfKKPorXIA79NSA5dIltVcJpi0y/op8zkULm4b+C1zTZs7KvxWvBS6P
tJm8IUQDgJayRyd2+6zspZRzK9cqtdBp5UHP6N7fCSAHDh9tZMAV+A5grPWOExAE
uue/vBsE1jU/rFNrz33eTTojKz2mUpFOKEUWt9NFcPwvCW917ZhkpceP4QFfiBQp
UB7Y9dVOxTENOHE1hf4yFfa+sJ9vp9aJnNi1XaAjh+uQrVtMCTxtwm1GiSGZLF6j
JTNxix5Z55UGkeIdcgnqT+XJKV4HC8jOrXnxIa6RvpZ9LvIXUnLtyToUK6Ze572J
1mC7xl7HIfcXyRVf5J6RJv6i7oo4R01lPtUO+RAk1D7hlO/Tg98Gy8SNGa/HpNJR
POIhg+7uy+WdtOinS1AEQzyvG50X6pGpdrpENz1d3eWnl/E6k+Rm0QQhGvXHLCos
Fj9Y+ybEloSL2eBlRAwGIQlT/Q+EOn+fvQb2u4bVY1UdTwRjse3qaA8E/llsKkF/
PlP2nRwFTSWBSeJb4XcdewyTUyynKBw/4yI0yXN4iBO/M4pv7V3sLFZrqrFqFpX4
/TbtB/tyJtjRRclF8A9mu4TA9VQlP30A9AiFD2SubX0LbbyOI7Rzlj8YPADvs7ZC
LlKxHl9ZMyJyiIhH2RTD3wKKhMb3D5PVWm+97ZaV5g+PxPAKNGNOfQFox466MOKe
P2TQ8aujHThHT0iaPmDhSYNJIuzt46Fw9kx8xL3g05RYXkt/HYN8n6eYjs4gzPXu
g0dgMdQ5q969igkiwnLgUdVeMmkyx67x4yi0duhgHgRh+l5JXQlbkaSxlfu4K3FT
iWTw0ukiJwSd8DBIEEs1DM7TFA2XDXuhk3AQZDdeNzynYR3O9RP+93cPoF8vKg98
pwR0UfpKR1WYepeTysQQXHfQFAfTMl58zCXfaLPhykKvTjQ/TK7Vo/fL8x794EjE
ewBD0FG7GzL/OB3aACEUVVjyriJQQGBv2D88JpkpAJnjM7mjR0YMFqviVJO8lE1D
wetw9stKsVOKmanYweDwWBJCLQJDCSloLbOq+LXkWHgDwn+XERUXX5Nn+9HMe9do
+ltVdmD+EiB/gkqvyAsU2E1uGcx6JxOhOMCbIkHIZDGm+HaBEmn65WJ1x5XQ+e4Z
8YGlRtww15NbLJZz+wCkF67KqLeLLsfEwbcC+Zp+idAKEWfEcHs59+laXANJc9kU
aqfv78mFnaxIj13OLcalkqbiHc5oEiJI7vnftFAKAwz89HrmsZum84SKFOJNZ/40
Uj1sFFcajON4AjciW+yV7MNXRRuwSh2DyQ5pVlHM0NKAUkGGvX1XAkH/XhwPB0KA
rBvqm54lPygDxJg/C7N7jOcI4gCQFent9HqaMNnLsBhAJWVx54JQyqF4gVimF8Bi
GpEOjx1o/Lu+J3KfYRI1TRs+lxp/GVBKoHdvakEqFSdgIUmnpGwpZIizhPnYfpcV
9t05uF+J5yZ13Z2T3SjPTBJaL37mCe5wznvfq3g0LsvDutkAbkwXXjozC1vZLHUo
SXBbFG310Pq7YS0u+fEikWWe4aEKWK1mGcGugLPtfVfhShJDGNf/uAEabU4eci/O
nS0Lrwf1A7NDE4ed8apOtgZY+AdJDWkd19tNm5AXr73I5UH4/MrxLa1EBGY/ZxOK
FvnYRerQgWgXXdYl6zYlirsiiFLCRJtYD1fH8S4aZz97+RoQ6H/mVPYxKYjC/N1n
WE+TiT3pUP0Zg3M13JTfajujFG3r3PTXYUyt1ZGbJm1W/ViK6it0VbuRq4oAlbO2
pYjuTu21jsoIVftcWaceJheZjdaXiqkU9KuIr3xl2w22N6COFZLhUc0OHb/uaRZu
Iq/SvPw0FF0e4rgPIQf1eth0gv/K9vZFY9WYboi0js9CS+4YeeDTinYSSt9RwfsM
Rds/b5oqNkESgLRNQewyAN/QpnainlLRFfKQrxkpD0H28ulJjHHmYzppCsQaOogR
9diT/kUEXGb2QaLASoAPtnSZWvMy2RU/1njZnP7B4dOGYsdIJnEj46adFgtJEaWO
9mNAb52IFA9XrT9/I3JhApZAcOyuzoQgOXZ1dWO0fffct0ZL7ZkcSVka1AH92pY+
WAhMEp3952e0hfu/nULTVRP5AcBZRClqvaMdHgI8hxfpNRuMQhWQ4gfd7WP7dDCZ
WNzIaGsrpnR+Ul2XYmp0GMAJyMa3G/qFzPidMuslee7zr1Vs5V/5QA2o9Gq/NlGX
LcbqhUABhMo7RyQsvmp5sr9eaDdlyp+fdYjU3KXTzDIGbYIL/TwDS7s0EqYZR2dU
1hEOLNBrE9+GUyRS7KSwhFVWQ6XM1E0vFhbO4d0kvKcjYc4K1FQUvy76Vtk2HB4T
h+bDR/7XapYHgFiBIFS9altAsxF+u1jJQNqmItf7t5upu+lDDDWwLxhCGiV15C8o
LPnTGuqc88NI0F5W+TbcNSc8VT1ljIjfz5QVTOMiJBV05g/q/2j12nrPAQ/1QIiE
pjTwP5LXZ8xQSREOYJoFRoTs6I2MvC2zCmb0lmIET6rHanFQxzfk5UJEi5HEJ7Q/
8Ro+zVYDch6h46Vuf0rYTIsgccMNt+0ZVBTygolPJA2xxqAHHt7as0o+0BfoRL1k
RMi6hnjBNmCliqjwS04u0jQQ+4jT2Is6XnKla+Chgdc9Y01xv2eNVUcTFDdbKxG8
+vK4GE09zScsCzrsMbVeEPDaKa53Crqjy7YTDHGvRh4gU7YDxFgFO1JLzN9vxqsi
PUWtlCgc5y/CIDta8oZKUf+YZHf3u7yACAXOfr/aaXHAGHyGqZ2VmU6ZOWUhBlLU
14qsGG7A/Pid70JWb9C+kvRJ9ISobj946bBteNZMJpYHzb5647GaSh1VSOjqa5cs
os0QsyeFW22XFDzhNlUZdouDOfrxQwMs5E9ovCyDOsvZj94/0N6p5oU2Y4U6Efmw
YcD/pSFeCUXSlSxaihPxK19FkWM1qIpOjXf3m1gSCFJ2qnYMGJf/NH2p59ef11/X
ZF3l141PKAtMDRZXu4TfBAm+fpit42iGzFCM2qpr035CABwpzKYnO7/zsTPAsPPK
XkxfnhkRGTkS95gbBKJ3fcsy3zyDctFFziiis+FVEO8SC84ze4mZf+++XzarHqSJ
7TtfhrmE6neSq4YeAzChukQN9uDRNb4QnzdXFJSKRvar9ncWD4mmGqA+/Xl+XbMy
rRwVBQU/4T9LtNIB4aRzn6ub088hXyqUex0NMq2Ze6TB2n96aSkb/eTu7oOy5lDz
6yrMdgarkp+ObuYB66Vh1aV33sAFtFmbCAhKqVNtg/0+65RGUJqu5nlGau+E9tWx
pDtFRSQDfmVOsbi6Vly0IUzI/51B8i2gL9tZuTPTGBm363VFeS5ZcNE8BgcguubS
2jAvBUem7QB1LkabO6IiiCvs/FSIb8d6n01ykcBIq2gyUpQACOQaj3Tss+wFx9iH
5pdq7r5V5fvu2pqjVP84wQ+DjGcEklKDgbB2Gqbt/lrf5h3xW+4AoujEblelZP+D
GNhEiWbzqRxeC+ZV4dSaaHlnUucN/4XOiQtIj+Bt94ugxLVifvr2mT9tQ7r1Net6
Aj8iTAEZ/mwyolaP9kMJPMx7oj1kstvPFqokjHLuGKmbdikerVkONXgwStaR1cGr
DYcqzWNrBibKnOy7SNS+XEHrgKgAssQeYmD9jW0/frzrxtsC9B2/MI4gRzDaBMxF
YZYYZ4sC9V5EHJ/wf8jesAjC1Vw1K633CDktVkAADcTWVrJ3ndveUJ2/AsBnejYM
zbRpOdmuXCpRd19MoTtzwTLg9NSfvhH+wGAU36m+C2oC/vsGbQ/RpdBjhU5S90lF
TKFGIbIdBQ/lEmy1SMIM0gVAc54XQbax2AJxgHo2ClkBy2TdtoHoQ/L507mecoyI
OanczY4dNwhl2H6hkdpLZ58pOFNdDjMXZ5ONxY+dp2o1cd/z76XQoqpFst7RAdAM
q10Uen4Rfrt0mrktUJbcMiTM/h88tYtWKtzXbmaFsxVn5uPj6dXRcfWnRfV8Sp1W
tf1U+uHRA2PYVv+womTjMPyAUHKyocGCmNbvL/4GDlB5/jirD67Wb8r4PPNozyvG
FhLAFt9FFbkaJBiFUhUrxYfJogEmL1RCX0IWVetB2Dulz+4bCfQWb/dIM0KrihEP
BPBibkOS0AiXcY5PKO0Zn9iUpGQFGPy0nlyeBWjUc+CFhWhDcXFJHsdrnWoTZ6F0
iR5+DgDZWnflvQeW/tv8dbh7nG4czZmettNHW2xTzqHHuQh7crdfdKMlNgRKZTYi
hUOILtqvSsXF3RcHTFVEWFoh43SzMXfovFykv2th+yyCwotMNYbh255PaHEShJCb
G+WYTWkvWkkYbrujHzmSEHx4L78Kj6zHUAmfLR57cbGE0dj8/p7vqj560lFMlmkU
7YqWyrsVbmYGVqeul1h/sABSfV1S6NwkQNi85QjgxAgwpgrq8joSl2D8jM+Zr17G
EBlSW3Wjo6iAF/Gq5p4VUY64jdnGvzjgEfK4jmvo7jtwwDZ51ZKLWMONqVs7hqxK
Yg2qExxdmMyTWnUOsjnUwVT8x8n8SJbebVakJJXg9AjhCaiHFdgV0F8jPJ2HbnWm
8tJbd4mDd1AJf5mNiApbFmepVtBxEnV8tFdU5EFh+n2vp3Nrg9HRlzpyLxINOs8u
BvqFV/WLJcEBNtZHrbJGY8Yy9bdS6JpL9nkveNc1MOIIVmDvlzvNIlyy2xSvfq9o
OxKWbpnpTUuJ5p2tNVtYtxdWXikErJGL7Qe7nzeA3AOAqbOwVCoPVS5Y9uki+Sqw
EN7cK9pFI0T2OHNqP2ENkZyeTQhuFn7ixaQ0EqbHIqOG5zrE+9Z4eEfSjWAyZyw5
iQgeJrjFuO3a1AvNKELtYWl+2tv7ogWN7CPYLhLTUwYJSXCZSG0MKMpnIYmtxhuF
F34ulJM0ou0MTn7kZybKhc3UF76s2Z8r+OE0IQLwW5+dcnYbEzD+1kKgs+0CaOqK
32awK4lIkUFvSb8CbkZfzA0wfu5NBKFKsEFPsqXH9RK3nY5yAzfyDpRtfdcOQ/FS
ZcnPvR99Eoq1BsfwXsdB5UXYdD+zxgmMKnlP/qoStV7C8g7e3vqzKuL/HwTZJAJ7
srm2QVpXe6zGk4u9lQWFWqKb8DZ2pKKecKu1WGfJGQsKKatQPeZCd9MckpRGgDI6
CldBEAG4LDvu4oUQA5dOwQ686pr7sE3xyB1m044LaEFoM28KWGjEZLeZI34sKKPt
IdlUF5dQ4qCiiZRCjpDxmpBxPCvpgrS9hJzGT6J5QOIhVdJWPT9l9FPNHQE5jGul
5BTVQkGVVKq0PG8nEoDcu7YWHltoD0JabryuADiPJOdw2xDLwL8h8/rLYTzOM1LM
daqp4EcJb+rxD6VqXtCVEariS5LhwQOhMp6lzfmYU+5i9Oo80HZ9CMYAIKFMN/bJ
0UpUQjfNeCzgHu5j3LkEHmskrnFsq+64D65CjxC0zgP5uXBzeMXDCy9dxDeozqdS
5Pdfaf92jKJlNe545ftta/xw637lXFkzKytCsihJqh3yUYvg8Dfxc9EuQHabg/0c
s5p9FyiTTaZnUnt9dSPFujKAkm5bfiRImCGERDn/UOJ2aNvwYkES6GAGQQpO8P9f
MhQZXPkG/9oTtAzKHwAJTgdpf7LQFCAB2Q9wJr85Dn7r7PaiizcuizN29B/YsX44
0dt4utltYdzxdJ4GWW+G1caAmr2NMpZLiPerKNmH8DkWug100sVb7kX9a2AiLiPl
krWT3m26xe2zGoR/fzlX+MKkpB7SmH2mU1XajeHvKHvXrLMasIKwQ9EAxmdVobdS
P3idlTI6HVHoPZ53lhEsQKGxRaMdxiZFCsqno2Bhnv6wfZPvQd6vRbAXoE1y9WRK
ZgvHX4wOJbHVC7352whNJjVCih3vZStf40JYoJivAKkrGQqZfdWM6M7vsC5/5nYI
ikFss7w+ACr1ZKynsXgMUcm6TUBV5LfrNnrc9PPEcRicrQc5H9EAASVaubIQnAym
sUpgISLnGJnj4o0DrHChkg/1rBFgMvYxZ5Y19LhSTxXaBUB5/lR/SgdE85Agubpl
496NO7V5BVc7jTEBqDJaRokX10NKL1jnnzcB/jk5XaxIhTLexCjmPOWgYLBch4jB
TXuMHFl3LUUcDYR1nii+X2dh8DALFGVQdy8eo235TLoBLvftiAziDtlq3DCfp6sI
V3DSLOCHlgw7ID0T7tetlN0M2anb96MYBPmKdLIY3RtkaGsIIHM9v3Ywj9uM/a4R
RsLuSLpDB926EkgwNbdAoiClYU0CoSD369iSLLmk4OjC1YYjOEkEBlp/7hcKiLHM
FxhXWbnRHIR+3+0R66CNk0gAYdO6ow0lwyX0UsM+lXJxPJnaEbZEvd2YESYyHJy5
AglnNEtIF1PjjWUfq44jHAuW7hlcS63B87KWQcV41jCRxORLVpHvmU+ca2VbmwaH
JXQtoi/55s+WIfECMCJLZV5DI/TkNE4hsitC7jYpiw0u7L0O6sEv1JNcc6dvhX5n
c3EziGR+pBx4HkSf7MDSCl9SNd+oHhbhfVAX0vKO2FtFr2KcQ8MKoGs38agRf3DZ
Cq7VRcgT7BrifPyy3QQZZDDjVGrbAd9xpz3F7l511e1+taf4iLviFQ8igjJfbv3N
329PAoQl1RVQfCde7FcnYevU7uAmgEd/T/AKY7oK9xoyuxwTUqNyAYIYt2gs8xrQ
2kkM6TzF2bBNqESQMR6r8lnK6fmlIO0XvWQjy5TQ7nnVqq3DpWCEK9mnbTGGLCzL
WFzyTmvRBOallHDBySI/XwtKXsyWnGczbRaluUtz2yb3Mf/y+LKtAzxEnY+12Kl0
3fdCESrx45mDdIXA7bqFciAaYUDT2LpzGQlB7dvy9ew7VKxd2vtvsYvIR2r718yK
IWywmJcqweVnnUohO4EHS2eE+nhI2ke7IQlLihLwB+uQOpYQUd4QNPHGC8QfDcH+
GOGmaBWh0mUw0PHeeoTYfwJE9UYCcFLKBNR55O2MbJR7VI34jojZey70qE/Rsoro
cwuc7sXkn0FvHB7S8zGx+cbVWm6RuZ9V6/s19Z054QSYbM9i4BNJPcXpKTY6DB0p
ADM0Y3iY+rP3KZ62/WxMLG6RKyX74uVQYdLQ26dD0ZYB//iv5MjrmW40rLt20ra8
LQH52suoCgqxrqujPzPCGsF+GV9v1TGcNq+k2aC2BO+mrwf/Mq7gzcuZhmF8dil+
pxeMsUN7tOxIs9pAMf3L6/Q1lHgcQY6HpdztRnNy/pTAkHLCbzYSxmzcMSy44dLt
NHOL7/hAjzl0Jr6nnPm+2/SltaV9tQNV0moStmw/Jr+0+1HIRq8hQxrPEbORKiDQ
dZajoPMQFCwTRxpwTzvTbEMIP2fwVqySMAsWflcStoU6rcYPuWMVOG0zpnx0cJiQ
dAGfkNjTuTxzvlYfwq7a2Do5uTd5CT07BfpcLo7/Gk/PNO/33X+lLpDsas1wwa9Q
c4XxdQ/LV89dbRNVgx6XHD+xc5ITMxw+GezYOa8g+QiuJR62uLraulTcQDWKjacD
gbx8Ugxr5aBWm8eIsAwkRfEwd1jjsI217ddcbEFNopWnyjbu32ul5fU+0dJ4kstm
drZAAeyfb0nMwrx481YohkJb2IRmZAgUGYc/NulMKlukA9B8Aciqvcbj8tsZvotU
F03ZdhKwd8CV/bD8hljgWtfyFioHalNDs9XVIXMFAZDTHHfGN/FNE2bzSmrv/qTo
sCmadS+rM1g3etnr1mRyVTJvIQYDZC30Ri230/rMMLiMqrM1C4L1wfcRCpQhMbaq
WKZRwfehvWMVdCmcl/ymbEgeq/FQ8sqOE8Z0AakmM4yZq96PPcr1Io8h/PGutStV
uH6dxI3U4gSoXDExDwYEy4ljxcOB7t/82eN1qWUPO1rHNsYJVT+R6biGF6ufES8U
wmSWPDDWjTJd6F/qXAlTtEqKIGwmYRDein8coNWbeeNF9esais/jMmBqTGZ8q210
vxj9gmJfBmvjHXxjc6yqhmbvnZgKANSVHvLwFLEbmmmoRAy8K+RiWDlQNZOMvBKK
wTIMGa/p2/k2CXUgstCBb8d4uyJxmOybECNVBoBW7UT+WvAtiXzzplL3bs3v9qg4
fkMWa76Zq+0kM+eqF2rBLXpQlZm1cznLKMzEEhOr1MNFalUcNjBkONHuFmz2IaJg
6x420v/Boh1XMfOu2f4p+KH68zPtfQtOEdBJOLhTKpA/9A3yVe5vfma8yNioTRsj
0h+itN5CqyD1U1yGSyfllXbLrwQfu/dktd1LlCnc7ud9eYxmYMXd8y5lnCJWsk73
iIbVljCEav4tBEAEpyMf8QtihWEO0wF0gW+zByrKUEJqo4LHH/VHeKDn0DyxJ2Vu
ZAs8c1begOM83pN7UPdx3PurguhDE2h1/WitYnNWEJUFGMlY1xKuEcR90LaYdpQT
YKHSJ/GPETfu36Aw7PMSV3bSK6srrAs826fx+wHjuS3otb//DUpx8oAm5SemQOPZ
DGVtg7AAPD1kXtGA6MHWhR9eUydinl/TesSnhzKd9+urT2HH4JMRw9waWKQOOeqI
jbr5xU27qeL4zKt0E3SARIN04m6Jw9sGllmQYLUK+PpKaaOaLAdiRa+MrPtO1jRL
hdzJITy1vI0GIz4YuSd3OeQcERwoICEAxeufafUJ+9JBzx0isRQ8PMn/ffAprQ65
Gzn+z21bexs5P3888zmpBqsMRB/+5FCmtai2K0ZkzarERSkOvViotT/L1tDq0Ct6
hh5nVyvVv0P3mv97+5U9b9535kHL03IYrHZ83uJf5ZO8ucMmBbEnYJTkwCe6lw1X
qh0Rq+oRVrld8UbF3WMJVs4NhCp+smsOIRtJhSb1WG1+99+suHcykxYFZtbu10xR
JdFX0A5jfjLuvFxU63yG7enyJt2a2s3rktUr+1luSNVZ861lYgHWncD+u0OaHJi+
evouAw68VKO0yigPeoCUzOFjEJsmXn9vArnA+zjiQ7i0TfafVjBz28iX+bY9rUJj
soyLMU9iANtBcCjmbWask4jmYN3VkhBMyN26ZfFiGdOfBnB1tmfEhzjzXMD2dd0A
ar+yhpgxLMlGjiw5CzYPtVDleDyUj0bPm3RS0jInbioZKM+Ed9ZxONrixF5Levq8
WBVQUkWSH++8l0L4+nHrbnz+BHfSFAyKjfhiKu/LiASOWE/nJHHWpKLfcRW3cmQK
I0/8iFXdU+aNm/whioI32Fs0dLbQq9zCQQvInwV+MaBi2d8xu970YJIuGxddgIpP
MPRdKzmjUkNQYNdBdqQJwxAXDcZppG2fUNDHDims3BDtndP8aBgNYCezhxVns+1o
RPoO2MdnEhn4tg3m5bj8uggxIqTjCbuC11lmJfM1Nqt+UKqaFfiimvfzNbkXGZX4
Nr9eqsMWzcyTCg8jQ6RMdpHw+KJzZIFjYmYfldYpmX1UsebxM0MOSZWB37oPn7sF
Irj+C0pMgR4CoIPUpyXQ4tvTUzbkJQR/NJHyhT5zTG9SY37D4JpGznIybChfaMIi
hW9CtfqrQllOTyul1RuE1rp2YZFN/0md2azTTlFZmLEAzUaF0jpxkp7dYLSeITe4
cFHspzniMQDYZTRZx2fAM/YvRGqOKtjvDb8dIGY6ve3vQppVMYJndemljfbFSPut
+p29NLroEP5TRv/JLJSNmVqFXglXwRmzp7yMZ5p+XhuXh58GGExwkhuoLny1Ir3Y
MN72MW6diAOuDa6Rp2SHJjQp7SP0A94YQuUSepgL0xfgh1i9aD5yMiqk9LTVo2BG
lWHxV5wgpvS/+nbNhTUavnyBJEItezWshehK/IW6NCgGQN82/X17RHE1WeoeQjsv
p8Fm7d6zJ/il/8gtu5XJ0hdm6uCRXpcqNc8rzXFZit03FJhUBPnpMY/qm+v67VRm
iqPlf6lM4lNpPv+DvW/0F+y8A/4ZwT2q5Utx/CzpC3U0mYhDLZcWBTo7vInjJb15
Dfsy8xI6VIjvlfLj7oNS1lWxYrGRjPcbvPL6A6/yeK6BE4uCXgLWIfeNK6Hh5CDP
/HJYKxtZzpXpZYjOf8ICm8XqF2pVXVBfCFbhWeXOJvuFgKKIhbiNy36DoMg9kjV1
DBo//ihbr80Yt8TREw6trpRWRRINuV6cFlP/7fljJy/WkPHc6yoH7vLI2RugTjYj
AmyWTZyTGs6fxb7WVdZvPD7DdkPKXcwXxVlDFoEiOJ7/IrUG9MFUDGEpx7PtpS1J
WtCCUm3G0PmQwgvG3S14F8oUjAWjgKeaXI10FA9QvplvOJ1eluuAhXkiSsdDkaU6
CZOWhw3Obhq47v1qwUnDAfEWQXF+TKD9pCk6xXmcG+DpKyD1IBNgi9UTXydqpk3O
zpQHjROyMZjgcbpOOyt5zJfrWmY7ZdsdyWXQXXSWnYZHr7CoV/WqqaR6RG5UZt7Z
EYlAc25Fk6POkWFsPnEozkSOMQARdSDH+iwaENIT/oATEj9LZm2OAcVYDL66jnkH
Wa+BcS1pisUaTT8ls/Tmkhmbg2Ex0ulUla2TTJDqJ71cVPmJXtfO4oW0yQEPvAjd
6appAtD8S/bVjSx1cXh8G7N5/jM0nqsG8LdK7O631fti9UdUYDJph59wjVHIeHOj
Hv36G5f9leEbjAL9jUaZPwHVTloc6atis1EavgZ3R3SqpmPFPAd4kVPUWEZ8Z1Yp
ieDn3lZidw5K/s9R816jEUrPFq0Q2ty1A8V5wiNMpkHYyp9UIZXeYSn2Rw77FZdx
QFALn2q1AmkFQH7/RwOPvcCPsBGnYtDq0YCupDGj6l9EY3tRPSJkhjlZKCFOrXbk
aNWxsZbcYguWOKchIiOzB4uhDZvaK8P8WLS6GS8PFpbqd2jY+yym90+hzDiIAqj6
NWQ2DQjo49F9uxE1qjuNwI4rVdt7oTaPFjD80xK7waLfhGrja2vbxaiwU044gKcA
7ncOr3enSO0/jFzdeZsVoE9wwoXvSZlJsjAgvKaFRESkWd5X6oZhUBvMp+lru7Up
9f4L9aQo7pDsELPYYQll17nYjGhHSa36f8MfHNLCn+vPLJ2qJmNy3UtjFhzE0cHb
XeGTwvwwJeXssrfEpNUY2GLy40Bb4fzKBN0fqlugYAHaF/Tf5FK2nfm23tSh5KcT
zQDVdo2HteGb0z7W/JG/ALESqtOOEvLvRRAqVCZOrXOxEa66S2ejOrOdmWhUzMIb
2CE1xTpSUFIooLk7vSUT2Wcy3JOMdxaujnTFSBfusegsLiB2AfIYykFMXlKdL3dy
1H5YygEVKyd2IcwRBjjvwytjPmOsLR+Ak/PyR8Oa0DuHnIcVI0u3qaIpSB8w1FiO
OKOguLIqnaAcjXvVfPTncps2iBmpHtnuzvevKDECsmHvPAgvjTr2CuXSoloT4U5N
nznFhjgEycLY503GvqW1JTfTlyfJQ7MKDutY0LDcPJq2wveaQy/5zuJZtaKfvmkR
YzHi0L8RTfqmLGduXkSetxd4s6uIEv8lAlIPzYcmfWpu0DanxIYFNTnwevuNLQSy
CmZ/YP98gvNpD/jML6qt6Dr87O6YREY6jmHld5ruZJ/ay/sWz5iD9gr/BKylNaB8
f4hRjBZclBSnPS9dQvagqb0SKcPZU00qVAi6T3ncWj1TZE3JLVdkBB9apoTQhOGg
Q8gL7SunvufcgjU3aABb8XpderUfyQM0m4s6K/ShWhcCih6bEuighDhVlTYyEgYM
svs+WrfmRak0umB0svvoOV16YUCcHzRshFxkWzwyEDfm5UPgEG+PI/f5sF2GWGsr
B12pJuUUHBkrKIuOLAnD2d9Kh1WNjD4C+bWGtFUCvZ7MTACeKlG/U0Mi6/C75S6i
SOsQMWBpATnGvgDAtVg697W4kAbjp+Z3OsdCVgfqZAib3EzrKSxmGW0pBA3v0H61
rVSQtGjGENr5DBMDj8ZarWBBjK4YXak0bS4/oQFWkd18TEJPQxSlnFFdhlaDgZO7
NcwMCVsLLIrDDd/50dkhQYbyv39uPzFRO63rV98QBrkhSjM9JUy7wHa0wUoa2mYy
4yWhCrbMcTsHRmei/0llOtlD3TnfOlp8Qsn3l6/GiRFHMEkb7uOHmMN+hyAZgUtm
IugbdHDmhdDQpVrn7vtrAoKUr1v6VHcOv0p4jwUJGjnAlTdl3hnbomwPEpxcLZio
/Z20XRi5uY8QUeccJiDP+RB/z1pDwA9ZqGPEQui/YWhQ4Pm4SerMb7g2TOMFX2qk
zYwJ8FABdThsPFyYRf2Qp09WaKNV+N5AqeKXxPLE0hvtqPPTZymGWERv24zwm4NR
ayC5QOOX3NCAVKiSHm8f/jQingweKOWrwEBQTT/XodEiBSpbL6CuUtbzjHVRrVh6
iJL9PxmwGeqWt+uzGqWFbJATqbYlCKHtMAVQVoPaMXmpXkk5+fDveeX3AGYdC8Hc
W4yVYJLdnQ/t1yEKILUM8SQGfC9PmWeuXwdGu0Z3ZAUnhbnp7l4LQzmmduXMRitt
VzmynRd0S0U0ljwIauQjFR59M7JyoLs1tCGlIsDk+cDFPtHk1UB0AQwkyI/OxAZx
jyzBeN39XskY9/BtasfH25A0gilSFm/9xUajh0WtgUrE7khYvipFcwtwZ/a1xPJS
TsAgSjHSCm7de2qdqp5Fohf67ZYg3Zts5ocWvLEoCUcfqfgxTOoq8Ho+vDt4uOHe
DCz/Me7pTluqTQasClE4mOX6bu1s9JOWF2xKPsJLlPyqpluFZZB8GVAYCR9wJ1UR
znaFmk2mjee5iECy0HFYHqNGPAx1wo96FpyGa8aC/Fx9ntXalZBW1E8L233Outxh
C9V2vNdtpwzFn9KepzYKqvRPpUsM9a0hUF18QEh/hR1PeCrEl/IPUxhVK4jhb98l
KMC0u6n41AoQr//zjLLpSsXFPctp7oZDlH7l5JHEDWlNeEmJwZHIFfpqZ8JxUeeC
BVgnNxTvrchvfuNW3lUnQx9zaEptVouBqHW1hxN2W0m8NPTodU3av5xqOYkydl6q
j/b+Uhe94qVixEsItr6DLHhd/U3afUsOmNcBkr8esxmdLfRRpx0+CqSfMSgiylE4
3nuf3I4+INgnmmbAGQPr9ppvZcHE3wkd1Y1z2ZX3xwaGDXpRm+cBYDq9w0IMjv4f
aUoNk2QXGgGq6B6f1JPHbZ0dwDjICUsUCUYzTeD4fu7ouikss0yf0aI5E1fM5xCv
uOu6krpDlK680oiV5xx8M8XEnmXn0kem6W8sg9TWvsHg/YFs7TcsSXItvHQ6Tx4S
m6gnkBTjMX0IANktoklofLMVHhQ0bjJhHZE4wPQpgwcIczex1oaNtArt84+jahGs
2VbzU7K1GJeppSYFnmbnTMPZxMlsBjlCqwIAfI70mQvciMEVkTJ5Qngh3JU5jThZ
s3IA+zoIq3qtcwbFFxBNatRKysN+fLcvCm+8+CrIT+vI/prwmYvNgruBxbQFaRYh
s6MCO9ZtTAMLcyyIYQcJDFK5lfG5l87mZI41cBNfwP+nLmAnl0FxwKQDyGxu8ez+
3YjWK2UQPQVpdU9PxZSlaO0CwLpTztfS1RHAfA+6O8GCMpCeqWlVHgeYmfQo/euC
nl4KICzQbasWMgMpxMpyZhaFAqtYTZP303YxGGquSWKUXVtx6ApAmK6x3bmMYiJ5
xrPN0KugAAbnAgNk+XIyJeqIi843wJs9UhluopD/V74r7yuXEi5PLSKp0JN4vKnR
0w0Wwn7KihmzdBTlQc37iRBUhcJMCulk5fd+CQIBt8VPOs3VX88azNhRTeSk8Yuk
uFN/T1lgUS5qSRnIHYqQ5ra4B0bgZaixLVQEV34eDoSTTrxdlNmUNiFjdq/vl56J
xS12yFJjPFmlDR4/b+4GcilTRXx1CIT55on77qNsKEwVTvYFyrlKzIhlUxEyfpzf
Q9ukwkm1G8loO7kBSFOhi6Zes902+5rsisSBZb+Lt/rD9cLCfW6XHNleAu6D6k2P
P9I11lx9jPmlqBk0xERL7MD0L919czBlmGtOQVX4HqnNy4U0zbIG3D1qWzXqMy62
//h6T8yeIRxftYe4A4qABtowzktZoyVBPAPMizaHRt+JMpRj7OjP1Yrk8xhc5Uqw
ecedmIxYPCFDDOfV0dch9p0sjF+Ua74AIub5g3vh9dbfdq3SGu7DcRHcnWcQR3dd
ehriuL0N4p/pXMK0merFaRXw6IVAmFB8sTZwG+ioKQKKOnpiHcpSXv/P8cM0LZO7
yuaP7LIoKpap4x6EjDRB2gBw6Samz/SaY1XFPl2dTB+bUBocO2cw6oYbiADsKhUe
wyxoKbqfdAxnDWlHOQLOB/8HqPKKh8RN8Knk8kal26DfqhAHUKrtlCWsAQjGkyvo
CD8dN5XAahRG+4hBo/AmkaDZQ2oK34Fk3ZoeVNjanEDkV1i8jo/NHHXf5ECRmKaX
+gu/6iRG+2eNpJm/H2I9Zb4z8BTAKGeVWPvEH6jez9bJLn1VDgZOofLZHBa7TVaL
QqU/b3lLa1eSuVps+13Vv8WbzvVff+3YjoX/ylERQg52rvj471YkyKbQIbXxQJmf
Be4vh0r8MfXrx1Z+kfyXn2B36Gqt6iXheyyaPqOH2girshvkOBzrsoK//tU2Ltr6
W/TIhKR2FM/ztbLE7vDbs8URnlq2W4/Yw0LaxMjWOWQ7/O5ES7PFtt2PIjCTPiR3
q05RfqkowtB3QyemYyy5nrkuuYavRk3EImGBpONf4a+JMFAsHsFd5F7DylLYle8/
YVS0goWbaBhTnsycovDpI4MgPflgD7mkoIejwMTaTG+1rewUHNPePoOVO45rMJOS
du84isPLBsWdFh2DcBjLW4xza0z6hKHAFBlQt7ZE+hwU+PORuMp+92k7RWdyB/+i
igQbm97zztHTpR33SYfK43+MZ3Z4XiD8ZTpcvrJppBDzA+OHPrNZvQbV2USsYQTP
14Z85gBdCMTvABeOkTMM4Fz66+kMafL89NYeHrACVw0fztKklLCx8GBSENAz2zaK
Fhsq2kEjSXvdZl7kMysA5Umi2QByoVJWOijwucuf/IGYxo2j31N1Ec/w8DnMn8Ep
tA8hcPmePx4nC/EFx1q9UHUX+PxxPowTZaE8PHBZyz1tH5w+yj3qGdhPHkGHrwOs
65iCfB2eB6j6je6wQ0dGF6cRnCji4jUOZatfeV8hztdhE0oEaLd4XYo4LKPsbUYZ
doliqx1aUMjG+8Uf0gDofis19fXQIyTKYc9a7lSsILLUwBTvWuDB0Sicxqb1GXgw
V7sTsCIjs4D9IhKnJDajaKzegbiRNdyp+WMoxFBWu+g/bkFlTJnqS2Az4hynldG2
pKLlDxkm8waLxVL6AiPKXQDqEOXH6/mDVxvjvE40BYYx0t9y9dI47U/Feqrw+f3T
vQyHRVVWoIpKdWK5zHVYqOfmyyr5s7Ywm96clU/mPCVDsZRtq41yuwrNb/wW1ztS
l7qTsNlypcyVetZfDINPORiX6MJ6JLKSX9l9PcNr7w4zIv5JMy01dMjF3ifcF+3/
twguwKjkjZCEuSzMhfp/8+lMEe0ZzvQOxcUWCDdEtyztuRQfb75brWpFM/cKx7O7
o264h0peRj+1xpg1uca5x/5P2AiMyFu2S98tlAeOARhIzz/em8+4V8y3xt9EI2A1
TepY88mPbmg3Ka/+pG6Wosy2mKBb+k5a5IRzI4uC3BwkyhmDjnlgytwKEMKPC0er
Jv+mWnYM4wbRuVfzujDUa+eD0qtHzHpZqeqWGVMgb1P6Zskk8fLNnqSZxS52gW5F
RvCQZi9iibxS9Z5vFr1jCVjX+eDI3/G9Y6NANSVPyYkFdsmtyeh8e2obOuZrB2wq
tlK1qrlPH447oiCWsj4VWXdzA6jYqFBhjoO1ad9JIBRW3kHScbMy+c0w+L697c8E
Es1d2+FxhAFN0latIyprgRRKxw+pv7t1JvCwQQ+vXpf8absCbsnlre4BJUZcCkgW
2Cw4BP9G7bBeAgSbSuDzSMpf6xNWV6UvyrpYB2X8yFTjrgEUIFbfLJn38KQUxQFv
Qk3BgdJmxExYAt1gQ0rrX9xoeBInlAI0zdZPxcQo8gmmszpdDDWYPEkz0KXWL1BS
ooV82Wm22nJsIBc/HLeTw3bwAF1AOHZAlqGnIV+Aa9zzHGTIJC7qvoia+FGi0KoA
q2ddiIWVq3l9sS7NXFt9HvVJpeeDnwRDtLNsU7JIIXuIOVEZo1Vh+2ywuu9uCSHJ
x9k0+IiMUjpohqJyTEjNrHrcY3JGZm90PCvvHo+pturJ4h+PLWAGxkHed0XpAXh1
yusK0Qkz4ruhF0vEWiBNELqkJRiogI+EkaRqHRPTzQ9yBo9g9VYcJmc+qDxMdyp6
iH0rB6RIOnKGDIZf1ARY6yC+0Su422r1lb149QFLM30mqqbQk1oGSDf4UvFQ0zPG
uwBLwPrwVisjgTmKnHLD+GOR9SnEtNB47AiLTaTcDSPGJZ0zQknv0YEFCjNdjkGL
rWZcet73mxsbTXJ60tDrIWvckIiMCdkWxxZ9y9KyocRW/qwmBcKWMtAmlo/FDQD8
mzLlK5xPmGDTzw5kMa1dy2Dh3iknqKwZBJ9y8nj/i3TaRi2XbPyazuB03jowXkXX
7WGw026Hp95dYuSnGzTZrW4XD/h2DCC9fLujYXDAJlg3U15zVzRHFtg9uEIruizo
6ERcS+7EU8PFq32sqTzPxSKSpXAd6abQNdet8k/pj5w/Q4g5C6u3WN0OMZ79N0Mh
zlExqJMXSMODlTZ1rX5pa+MBwN9esZk30DjPUWvaJ2d/dhpNsNNCOiLxnDSDvcHa
KQPWa5B5MlLQkZIQ0BQu/TbsLRV+MRkxPKSbMkddRb9w95unFUEzYGFP6vLjqZPx
EUeBjwU66YudtCQz4OM05nzGcbKNZxbIGvjcniK+22mtfWWs8sB5Muqg9flTcw7N
WE9KTds5uu3Ote7V51FQdLNZRQYIrV/agDX6Zj2SpBz8fK2e1SYDcBfgsB0aDS+0
J21iQvKtuFRt8ijwC+h/BhFKks7GUvCv8FuS4lhvmOpsCiiulUas36nCP3matxWg
bE9A6u1NqIb++uRLHv3MS+XqcKXu32UgpqVWzFAwImwLb1PX1fRLv1D4oPRb8Jg6
cUULZApqG56muwXMtACMzGPFlOxgzsoupurbeN4q+O+KyEhSlBThmp9jKdhDGtJL
qrbqJQ8sSK0eGuhC+ovricVJQykdYUj6EKQfDZqkGOHcNViIO5ussFDUhsHq16r1
zBspesKnNVdyVdJmOQn4h6Tnx2MkZ5sff+M6cvO9Ih8m9F/YUoYR+tDnzfew/5Sr
QEuJvNKKSaDme3BYhIQlY+1ykJh5DtzmEH4BANQnCqIAHxaJqRQDrsDFWbNFMVkI
jk4k8ReZGMvIL/OGw6x74Bt2V/iJ/rXf+QfFsWdQ8hTpfAkFn/uv1EXGD+iASo4b
gHE1FcewpvK7c1bwKWH/ZEFlPtbQGMIus/MJewIX1hWFGfj/TPDOwsHD88zj92Pc
LJ/38r0KumcvS3mel5kO2cY3C6yJGmY+f2DQfzwTONw+PeJBe5/KebRxxoc5zhTh
Feeboj/l4atzhe6aMdrO7z28mCpZdGe8rtsVRXVZN+OXeYWoGtgSZjwSUnrXZNqG
9DykReHPzGAhNvlIKvb8ItAJeFz8hjOMVuW38QGakKq7LDrnO8wVdr5xqGmUWUI0
+1Sem1SDPFxHibdVmNsrpUjvywlPaMtQ8dypSJzYzOwjOkC6rPBeQcBcdm8hgfp6
RBf5WhUTxZA3Zy0T1s79F1xefGdHyN1U3AyB1GV3no9YrJDYy687pIGJG/mcoBx7
uxfE3QC5X9xa9SudHpYwlupjM56NWPTVuSkHgvGZUKkfyvqzRZoQh2IlST+xAix+
4FuZOAdP9Fwi7IKLnEOS0c6fZ5As6b24JXNrvb8eoEo9GfvSGF1Sy55cxrUri6M3
dwPOieBBQwrE8BxiD41whxAUUXsBm0QxblpV1FRyeLQbryuGxPvFrrMYcIMYd9PK
o0/tglHDMGA7EUOmTDeriZ01myL9xUHpde6J4FLRgy9pREepzIByQciyaC1kBrVb
pvRbwObDewhzy3Fb/r0gEABXQ52G++ilpcHHAWabRHi3yfiSEKhcxzJSuX9HmhPU
HYsU13ei2C7Oa5iEGCYOK2D+cIksyMie/OwodMpvgM0OyoK83Is4iX/kSkBmVQgO
RCpuNd17mo1x0UrUv2aVVz6JeDIwI6MP7VH5+Y0VS3LFOY9rpfiRQcOWjqrecosw
YOIhFwXZloW+7ZZxA5WkPyXTk5iNBZdNIbbwYtYZP9lGE+EaWHLTOL/RogsYnitc
Qvp6vzr8W48APp7dfueMVKq2sRfbe1melvZuV792kbwzEpQcl8rYroZCbRiNpxAf
oVIx0FSx1lRJ2/CqOnQhjbayiE8/9wxfSFwIBCPUIC+TwZAcJglVAMZm+DPSbhlw
6USjxbRe4cXteLgCysDJxHW2PkEEBoDdi2KbFyLhe9IsMj7IWz+MnF2Y3lBdqJmF
KX8wr8ipEdpYEcwHEnTx1myZy/6f/27uAecaVhzKkGftoT9Oe7I30AN+d3sH/ZiN
pQtQbn5M+DZdSwnZSIECFibbJZ90oKhPFLJRegSWh7wq5IqxvwIqnHviHlndqyeZ
0Hw4ba+an25a9dmEvPy0dLLXnjBg4KdG5NiweV9DQLfa4TN52k1x0gTMmQfujOEt
2xzHMAEZ/NxxDH4+r9RmcWIGl3ib3VvEi8LV55r9ZltfRxJVmOPGT8GZ8huGHGTS
IxHMfidciLL3oQbryro3SkB5FxXSOwOHp8zwQ1L2kYmwwLEMAAjIehgXWb5I8wKw
GG+Rx1HtgN7ZZUYTJETm104MQkPnePzi66qfattbo64EByxkfYuafV5uAYbsVYOu
3h+aMB3fc0pChYgPNkVWnQVFrAcpgZ4GoCwmONuLYMuYIp8V81eQ223YJJey9ZMA
7Z10qPMxL2TwkIl0MRTsaDImvV5RldhojmB5kB6Qk30j6hKxh+YtXK9FkhrhmDfb
8ih/GbpcqV1DuH7JFxHH0P9Vu5aKoZAUzrlzk9I12crmyWSUbzQ0bQB4tHPsGKdk
M3HnuJNJ26+dPcKl8VaR/AaIv29mSJVYzqt5EByCwQMpHOZlvPMA4YUIKXWFj3B+
YnT2yeGD/E8YE2oSBfWyOuJd2RzBFvvYiasWuAiJT6+vPN03bFdryqXs+zsE7MJP
GCAI29GQvV65stPPWZv/4xZdn8tgLY05skAhIlKx/LB6ym42SfQdPtHU7yt2BTr/
BHN3YqrrOqoqKRMF4znyoJo/QelvOlmuyrdmaes2iO93Gt4Ic5bxb7KZHEDIJk4l
SX/4cyBFmjiSAQpeUWUut4KT8pV+qu7fLDuiqSZSlW0PKIqV2y8WBAlLwQ4E7mcs
T1bn81+4Ym3EFkfVLnspCSLYq1le9XIUrxcSr3476IX/+wk1OI+Urk/xjXuEN1IB
muAW9O6peSQkt+cvyWax91/01BLtWDPJV/tS/O1vrPPI1tuP0OUD+a/0DneQh1I+
mEFrlcOGyWpZaiqO733NcR4zxuaKI8h4vjr9rSCbicxF+MkrupabAtWcTafP8AQ2
BBSWgPy5u8otBBk6mCmAKWHmb87XpDfuOzRik5dktZwlgUAkH/qskF4AFJ3OU4nu
fZtwWpkSDut0Ro+APmqPU81zatGkWeP2funwTCkd7lHPMrdO9iX7/qxlFfh8UpNu
g+BuohbhpBMWQi2tWHEJpzGNIWRjoL8W9LA0ONKxuzrguToPYBMyvx5vcESkPwoz
NxIpA0TMV/dzX49DFpXyGnkc0o5JjzPgxONgCW4W6SPtkf9XNitM40H0Dte8EVm/
viaI6oJXuE+AAI3mi63DZhgWuiJIJ4A+ux0UXR2G/A5XNfIgCjyAhQLO5YUXw8c4
UujrkMiYJewaN6DeDTeIP114+Oy1hMJWwRkSfw7IXCXL5zYlUQvZjV+JKjej7WsR
o+uzmkpf8p+XGp2a7wm4MFpX01I6yKhaydkDfT2ZZm0qDurA5rtNdYgtKruItSOW
MK/8nnHlSnEUa7zhMdL4qLpr6grXQURwb5SEuNosxxa00raQ++ctiSSHsebb5/Vc
GSi0vEFpKfNbwXLqNYV9u/hPl7ZM6x+M6irlDZ1a+awRT18J46cZ8P3st1CRKYnI
+9lshVxnJeE4E5K8Zg4UkmbvGULNvrAvWunQrDAFsleaCwyeFFuKEN5Z+L85UhgK
bZOZ46WVRlp7J8LxZBILGt6QQqYJhdQEmP2gAGPIzsP1ahQo4QXvqIydLbEYQzXk
I8SPy+rq62TQtTx7s8jn7ahSuiAFH+Z2nF8BNBajH/+KvbQSCJw1JzHtlMCyhReR
kdcKl/M9NUnTgvFnprhA0N3I/NLkIrAiB39hwpTAkWpdSmogJvaXvRmW9gBKzghW
TXQQoEiMfVJt7ltjbCDr2iNu5Ki6fhwE2hHdzgNj9m7ZHwbsuq3cS/5brjCSRMru
8p+2TAlVqsGAYPJRKM0GUini41ZwcO4jumz40blVWu47GIQ+Hc1E8J85DGf/fA3Q
3ICEryubkC9HCz2rVq/ib4KErhHwAkOK7huJRvnfWxEuk5nWq0+AQE1w+DIJQb5C
gNCoHhrRIq2IHaDVhxIuCVfFsPOnrfhtsRWusB6jUbt08Ze3SN5gda1Ul0jT8E4h
cGYRvwYzmJUJFduLGedF8I1jWMXsPAENhs3CKQir43NT1PQaJ2hE+cXDEVq+0Ang
cBVhAMSjG8UUMqzTPEDNBfhl4I9z20xEZr8aORQfnFE+hRmRSBD9OpeDsvK+I/sB
bvEktpqhiHo6VjP7vzXP7MXArUpnVSMNMjP4KxzuO9mw3JtdmvGJY0CDW97TYVaZ
bqm+V22HCjiPAdW/SZVPL7ujSEKUnw5d90XhdLvCkG2KDj9QRd+a31Ts2LzQGZ4W
T1TB9p0l32xWnKwnoqKCd+EVbNHIKcFAuqxQzAe99f2ZgJAgUJGQKSkwXIi2bbCz
FccKkl7+Uv5Ugk0xJZwHzhaSJz5ycRWty0nzDyRTh0GkqQA+aiiIhhNEKtGSL/tD
zH58YrjzmYzqCCQpQROoriKPJ+9+COs6iRflHsLgBdeUaTUiOBhPkG80wz9NE7uS
CHt/lLeAQs17sf8zVLutEyLsiJ7OrtY8bJr6dg5x8I0pl0nGdyAidk6BV1fIf7Fy
cMgVzwGUsAZxmEDdzLiT2/vFnOarJ6f6mbo3yxb+pnzmBm9zeUUFe2p8UJZVMccT
I1kmdLZcCuwNeFKkTcD5WEnvIH/kYL3tDLx8fS/6q40gB8yN7HOVtivXTPocnoRQ
m50iRh9fRXxqtDJprrx5zQIvpfFesEz+C/R2tamnQOo+4Tgr2IQOHHvw+xJRZs/M
i+MxbPU7O7fK7ail3LvkhcQiusWfAi30gbQMsZ/kcnLWRCiH9uemI1JKgoy5rctx
FDDZ6vq4B2t77ABTfnqKClMNkmsl5K5Od1QvIVRV65JfGtzaBefRxe9GQkXcXtnA
KGjzm2n2Oi0TYeD/F6JLz+5l/mnOK+tXhBhVzRUT64JSkI3nceEwHbQjBkb7sjc7
nSenTwCPjQRytlVpzq6dMCdlPu+DCgNunoUdRXMZx8uGS+8ejPI8sNfISrEcrwBm
+1t/QTXzlVSlcoZMHmiCO0DUEpYDPq6q5V/CMEBh3Rtt+LsspewhjCRkWmHstFWF
FXF46HGPqb//DxDTad0lyG5mlNkn3YZ7yqmNe8GjZ/Yg2+fCxG7Nc1qjdqUa32JR
d6+wDIsGHYckRv4byKAmefg8mpWwIqqOYDYXtJ9bMa702Zox8zvuT3CMeZIyIlDP
Ozn7LeI10RMW678lNROHNGwjwDx6fFrSDEmmvpGMcl/wUodTA36/WfVLeF4m0OFl
hSXmoLfah1XsrI7+yOa78G1fFZ+O+bFlK4A7zhqwCPW6k5yxwfPIwmrbimrTUF7F
YqBb1LP5D+PDdqWJ0ciKER66l0gI3ICZHtyS1uZVFutf7NsJ8l2EE0jHtGg9ZO8M
jdlo4JYkKjdWtSKBfvy2gneQF7hlft3UpuJM7cRigJcR62b7MYc30IfFoIDf8UYN
S9mtv+akKx3Al06fPJo772d0lMIvUurtW5MdHt1CjhsdOkCNPBBvt1wvqLpMZyvM
rhx3cPUHAWNV2brOS+akP2M1RBAfL77PjknwxwJN6SVNpxxoOcdvIQNt8vznGROW
7rkgm6SCvgTtXYNnxxp+vsN+1TwdF4h8PXqO467P5SI0HSg+czNUf9/RFDihwtZK
k9Y9QC0ptNpJhy68mtsQUnIfwLIaGiWS+Q25kW8PZZLalOAsPoanIAsvp7CJYscK
0i4b1qOAT2AdF921YLWH7N6rqaHR1TPflAVf42hgVZCBHiUYePcT22VRoA1bJMiI
FEuurFglcMKHcLqZ13/2YZ6kjvaAXx3HYvr5E75Q3fSdJlT9KHSpC1c8CuhuHJgc
sGCIrLsmXzsVD9EMNl0Mfh6IzRdegRq60SzmhNv6nXCiRvmCPbsVFffxhYVfynLa
j1XigF0N1n+LCSjsIwQsTfHR56BGgdp6hAj3GU81rz0Bw+U4mtZJWWsC3Dgz1VcR
bSLsYM2QsQ0ER6sFagWwUh/Q/eAhGzdg4MV4TTop9aOXQlJwX5NPvl7n5+hJZzOv
2YdRngdec6GUF9ZLHAmneDeJKcC4zSsm4cs1voE3TNsKzt1Yu9d7dAYrRCkm3fKh
vdcxZZIz2CA3mJI9gS+xnhfmmQMi1pZ98P4eJLZOhNbNmtRSZUO/Zz/+8l8uoJQG
XSuywf2+okZpTGpayoELgtUNMw1++eibQKJX4SaeCfGq0xzOxzrH1CgRXr/2DLij
TljwfqGLgGcxpB48DgKEoe5eWWaWXR7H535QZeFcCXNzMnkicPsRQ/J0qSYRHR7Q
N8Z724x0LEiJlFvMV/TrOXnBKMwlKxCQcG9XDcEPu8BfaCZ+49hrYof5r9xyYGD8
UecQKRQCylRxKxzmwuQE1mCpUdnNUxCbLSlVNjR8TJCZ+dVeI7fsts/CQRCQB8AX
JHVUzMfTvMo6MWRylHfcv2sewcNQl2sUw3SWls5UCCyaARI9tOeGMwybVwSLGzUf
kbU3LMbYHDaA/eLs6eHGmxAC0UBmZ70IkG7PvO/vUzpLzxMEEYZomWf3JngXIdsc
2VJJdEVAJqX5biyqqZHOJOYBAAqQ5dDzTTaW2gypnv+MCOT5LREqp1y2L4dwSnJ8
1eVs2esbsogIjYAuUEZfGvYpUViFnHzrggPI7nr3MsfD1L+Nrnrb4cpTtpP27S3j
5o0IvH+M5B2Td7wGobNniszgIo/PW3A2LKUrFeggbVj0CQrBZcHG+bgktalqjRZo
kS4QkCTqd9KQXtY4a6Cm8RGyGW9la6j3k4tk2e3WcEh5qo8jryrQZMclDDQ1jo4+
2BuWTcyfqNjvS8i/df0rfMGfkKgI1hY7N2+UtfjbaILRaBylmqTBuG0dlZbfxYex
KIEkhHl1HM9/QoU5LN8GM/9OOGu1GTv+NLNWZXft5K4UmhxlwTe3k8x30ziYQ3Hd
0PfbOpHJAEcMr9IWtwcWnfObhklJIMJxsNX3Mrie12URrxl0CtgnI/DtaNMK7IzH
/SLxyGItCJCVfIOjuHrvk0dkQi1hwWQrxPIlAVObSMvbm8Eh001qCdzVnCUFO/yT
gEmGBQjs3nr901FuuhlLfgOvZDd4+5VFRGLIzPyXbcugyY6vJlucS9DZhBMtgmUc
4PXvP8ZoDw35nKXhwvmXdX+tEjHkCKvERR+8xT/RsEUE1AdriK+9ChPL6mT4Dl6J
hqxKxB3JQgX54jO9Z5QQhvukAZp5XcUvIQJ5lccYZGxQSQjNS9nVkn17okK+ruGk
da9TANstKk2LhaXfzoGqZcJY6NzdnJDr+o78KncYQLZ+8OwzW8wFm/Qc5ZxXvpvC
AaVr7ycyev6UOEnuyZ6p8XA4k3qW9GtFtT6tRLIVdZp20Jby4kSAzuFnawjqZPq1
utXnN4A+4exkGJF1TToaBgNDUDxjK0SZMPSFmhOyQk3ZSQNhvRRzpu+4mL2vSJIZ
KhrwoQvd/iY5v0BS5srqKswr1fPjKrEFFTujyupB3A/e71fnXq+np8nRfvQJXvVA
3eNSdUWZEcAkOOoBkLzyrcgHyqy+wIxfpXOq0ZYe4UHFOWr2Z4065FqZX+1/n9qG
Bkml/A1aLf/8EeOuwEZLy5Uk5JrGXUL5/brnJrRnY68FxkYIZgNJcvhXAFJdDAZV
2xAugytze2mIcFOsu0gM4onmi7KEW6yfzeyvPAa69zU6O4Q2vGEbVgMcfCJmMTfB
ihoVqNmlj9/0lGbZlS4TSogiwPmzRyh6GSif20VAjLyFkjDx9I8spe6tpqSpwnnb
BZOsffM6FriDheNpcDpTMtuUEZVWdWisUezkV2gHsNt2Rg7WeD7nRPWe1DjOnr/B
3ti/Q/qQupiP0vgj80AySo3R3/Q6DI8ZPW9E/PAOQhQnPXfPQ+zkdfOReQsn5pPn
i5A6Y26SIp5Qt5maLA6no6a3PeB2r8bl5SzzT6CzzOjMgs4BNWU6dKeCOu1pVcpw
2rf7ed++a8LU4ZW5zRh+WzaGl3yDuWtoz9TvPOAtYkIEbdcY31rodCq6+FObhgsG
iQ/AR7/w+n3fDbcgClvwHaMJE5f5XbgYWfG6vtHF6uJGPYEGwCYjQolEiEwA/VE+
nGOQI+DKe3sXk5KE+I6OwBPPyxzvCl4zFYU+B4z7V3VcYSE7u9FhBl/ICqLTbPaF
zcr1CRZcaUuEwWYuXwD7pU5HFR+BHRmIrq4G3bo2GflRqjJ9UXZeJNi3xs7QGtOz
+703ktxsL5Vl1bdhFL9uB/ZgFx6zut4NO9KywitWlslJtc1fxPOOBFqt1saksMso
kTPtngdtMfnsz1+2UmWhwEcvk3R3iWtsQgEFcv5x6qfSVqFdtcDoQEKyl/+75Y4t
Pj2p5ftB7eDXmQs/NVjPJ9cVhcW5uG2NA+zliOjtyjMJhOPRQohHoLz7Se+q6u77
b1oQ8V9v641qDoELi8uNx01Qla0H6/KIsszQa29tLdrTUvu9BnGNJQGslPiXxeoQ
dlaQuG9tFIkSnlpIRpVCKZiyczF8g1eYMD/AQx34mKpBxG9OXjT5C2JEiF+XKzce
d0t7czL0YtmgEcX50MGmdudhoqcP7GXRpVblOro5AIaiBzywLWUyooEHYZyeKTAP
SIOdecc3zyXjFmIx2pcuetQKB6h+kM9SdPeT2maUBUe0DZ3mXVh6YomkbR+H4oBe
igWUbPgc2BP4BMVhN3l48OFLMyqbYX1oEM4laL5JkU4mqFV3xfWHD2ztztGKeZUV
lIYceeID3tiIPqatxQwOeaJje2uHgUuDaTyoVznniQZxvZsy+CNZU7cu2qmWZ3Od
kxtT28a/01psAi1GKzJg/6u555mKAU3KtNrAotm5WoPzABlHcZOz1oYxrGBHKXeb
pjXkdIR4kMe0/kJW/YA6ebAurpkBUwfOB+ixoonrKJQni2euYlh5VChD2Qxe7n7A
VGnwcvNXgo3rZkSc463qGodOIElArUooYeSYFjIO4YITpDnUJ/a9mroY9iI3qq+N
zkK4ugBvdVrAHxkUrZ/iL7nwFhne0DlstHOLgKlHvzNDvUa7drJivoMgk7qPqP48
sRfsFauM306xAKnps72kCOTHQmKOk57+K/0/NPcul6RcteOiiHXBnyjhdJHnSlyr
UKqOT1ePL8ynv577R6V11IOzJAEH3kedm7GO8tKlfqXi60ZHWqGHWla0BQlN3Ya/
aUF+JcvVq7LkpEXOa56stO964BnbKwo8FtFLAp8XT0zUUFFziEOyRDmihGxaRiTa
LmAXMgLHRNq1T51UKPIc8Q4puTS/zHwCWz2lSYqcAiUcH0ILNdD5q8MbvnrPYvUB
AtcMyVl6/V4Dru+2SsBdNu/IEzNG9rImjTyH+dsoqpMaglhvEwppgjpThS/ocT/x
koigQIRWw5qqRqsKbmupe6hZF0F4AVWr4hlOuVwRu1uBPZa95mwMYG46Mt4MbvuM
gfh6hxqLYW8D57Jjb7l4+luTAfVAP+y9PTy/5yQ8Ep77+JLWTNVE7cUaTfMoCjTS
qZ5xtTA+upTNbky4nkLKxBie1vabSwNgMADxmgUx+Fer6X/CBwxkGG7Zt0+54BEX
/BQUNf8cMtAJ9yqzqRrOv8CipU5osnvh5EYUWoDmHB0WPPplTTLqxHmPOtMv293x
Q4FqaSaIBSacn9BfdxBasMEUPhmnQmugU68BLtjpd09+Aw5mewego+hOw3wwdERP
mMXqsCJdMYhsDhMocZWsxe+7S/0cS1tfgbtMpevePpx+5KZmO7iIV8dzSp9FpIWQ
CrPTJZPZQv1fbvgzeahWrUKwoigu4zFDoOTfbO2bA+FHaN+X174zJyVEU9hTipa9
gPatHtOPig29r4E6cz0BEhq1s7oqsfgt/WB191LycKFfVW5rwkFsRZph+E/Asmxp
o5A+Tl5grI7y2dXzFCJxctlv/OhydrDf8trzS4XNIAONC5UPYi17zHY8LTEIdkyJ
Ibv9lkt6d2PWwFxWO+xvfu6jsuEec2n7eACnmdj4cEHGduhPbHRAFG3YUNgsfD3X
2/TMQEV/BwTdSjqf1Sv+ETK6i2KNJBNcDaPI2C1KKL6nc8k+9OlKOAUSXwc0JIMQ
Nl4axdVMM66efKXP7dYK4ZLF9LHzmqTAUBdAD8rNBdXfKxCfYPukikKdlGA4XY+M
dWYnMdZ3tIMbko0bxL9HrUz9oj1Z3p0pbQTVJNcUmaO6gymKnL7bF1MHp331dD8z
Jz3yUocl1BIVsopwN0L1kX+OK5PBR7wpSxAiHpsKJcE+wSUxATLYi32PzOUbjrNv
EKzrVV11bqCq6Jwu8ridyIy3LKcq02lo8VxoKn/QQRSIfAtm8sNOg4+eACdLnItR
3vBC8vzJisDbPXc9OcfJP4hVcY9nmGdtqvMKwa8V6oIfnEuM+gjG67QYVlBwxFhz
zaFfr+AULhjM8J7jOpy8gRiBgmRV9C67W3IbwWGkBDtueUnOCZihM+F1cMLQYGNp
sDiyFD3roPqAMkhFsTLQ7EtF0TbMxZAnHn2ikXfAuum/HiLvCfIMk2RQnbO0aTWF
hKKIJNZhKjSpgAcmCBM/CVnGlRxrUc9tpkKjVVwrXH9OGbSwvjQ5SfEtrbXv93J7
jK6WkMa9nvb5OkC9n5CcwoywvvZY/92PQFp8QZur1BnF4B4sVCce5lpYl3hLLq7X
WqAb+LQ9Vns8a8zLGrpEldvL+M5LjyUqJvTPyXg5gl85PyOm1dlIWcM/3cBzGLL+
zbBBqrl64pyoXHpDn1YT88BS3S+LiuQ9SKEGMCWl2rD3UV7F8aOTIUi3pOOehHVR
jXOmfmp1ycZ8ZWJR3zb8MPO3M5KvDkAtabPsA4sqgJYwZJuN4ZBrVFBCkRIT4bBX
6qiPaRk45C932BdsneqL6U81mTlIF1rRZaqTKYxCSfErzN9/S5XrTqcO0bqEp4o1
RTytP+hj/h3Vk3MWlC62pUABMCbAShkbrr/XwFmjH9DzvxqNpwNQJyIHGQgJAA4+
u9GQPuqDcZ72mHGfRj1dtP4lY+Vg5obz6jfRxiRsBMH46NYZVaSJ806MKxwhcJge
T4cob+CNoU/QwOxh56ZQgXQyJbvz6rr3xluw2PgxtzAbqC6g2LrS64gYpqluk7oY
zy3IQZJrvpCepAunUrQejHqZu8cKa07Ajd5o95Gf0G3sAmaOHYbTyExTuIPDiFkb
TL6ZsDMig/pWZ+N2aVWGZ2cWzMowKe1ODOpOmIRCeXMiehQzfMZqdAPNunC2J9Ji
OirANu8x6ABv23VVtAPnnhzvkOn0azFXjtQ+IU6OGEe21y5IIULHqeIUekntcKch
uCZJKvLJtSVIpqJ/5h/S5tvgNaJEjXPuPxrxo5tUjcgPGaoNJbGSuAaKWxJFtblt
Z2ZN30ZuIykKdlNJ8wg18Fr0dhsVe5JNwTjz6Po9+LlugcCQC5mNEAXUrxtoNXC7
B5jZqzNirVBIFp4aYpsIX25E5o5OO2AcUSulv3d7eO1BINbp1bGrjxGWSy7jasbk
kFrcH06sxfTFW2GVfGQ/wfIIskROZqjBn4hfWxRLhsTQNp4QayVWm12XhubF+hn0
XYcOm6G7wPp8QfjrziNbOtpPEDI3ahfcE2zTVjCEubuHHIN2ocUk/DueVOR9YV7n
Ze3gxOLTBPk4f1XwShpAVULSR0TMkAu/O3PanIkaip1n7H1Xh7eWiorXNQIi6DdV
j+6MoG+SBUzXrxVoTtl0f4Cqt+6jOYVCHh4J7K5LDV6ij8h+zkMLnxKp1py9Vtnl
cgYLQoBm6p6hu9FHVVsn1564FcdNliWRKK9ZaiEKC6AerplhcLt59bBs5tqjl6HZ
CjC3peEkVadb28PL0FzG7ns11Ak61ibGi/FaX34n30O8xoEts/lWZLUurVMNJYAH
C+E3p3/AXYR8oHarEkgQbQZx+PbCdemUQs4HN1r9D9JWhwk3cz3WIW4toHzqmw92
Qths60Q9Kjz7ZshtEdcYDh4ifALZ0sdtDd5MVVlnsr6QryQt8PQTni2lKzWdb/S1
8ZR29XSG/hfzHdY+lJOgkV5ysJyb0YFlFJXVJOtUQ5GmbKtEYLdH+usQ9sfydRxS
3ueXX9+vuFyjUbQH/kbeR4fQUfjqQADz0IPrNaXuUYgq6dGbO1PyKUhTDalLfQLh
ri9p8yvFYI51edtzGZ6HzFn/OIeEEwk9HFlPFrMjUsZB4d5sPXEpRlMWkzn3ts42
ZYzzTdYWdoSjIo1XXDL9n9CpwChwkgelM/YTLVuEUnNY0q8FEk9drhFCy79UhRN2
NA1u5BO+NAzDFU4yUPGgh0Rgr1wm5xwcAPCCgj4mRzYPZryIB1xz/P/k1AywSXWy
zH9RgiDvIdlNChB/5Ri2pAOYjPLcg/Rx+SD3kszGBV0cZ4b3OAGUGlt0luLmqVD1
dV2njvPLMBkxypyw0RBP/ylIt+jSt+73pvvkB67HHUBGejBMd9ay13mxXq+88YD1
7dM/z6V+MS+Hp95PXijQ8rJ2SlVphIzpN0erwUMGylDXYJMTebWdJw0AhpX8wE6w
411JfMQl94HAxqG7QCfC5Zcs92fDOzN6H5guo1cqLKn34E3eDpi1gCenarupfdIn
aGPrTwlpH4bZKPVcQhaluH3242apThKD70CpYcKMxMLTXk5+fNo5p0xnJOMtuBr/
xnMryRSrrA4epgnPp1q7ZYRJGCrHlqHnHa7CDYjtb7HnuHHSVDQoJvEPGDdsp5IM
RnR0/gZ4TuOJRa/ziJQqv1EhXwRBfh1RhNiZKfQHJc21cCTrk5efenO4fbvel+zL
nEO/+NLPcL8Dcgq2Q1/VIsSn6iVXThBrTL0dSukxgIA4a9MBPH5lcQH22h3afXl5
m5qS3maz7sCcJlNHnxt6MndSkdMzkU06mBd9Btc0wXtTIa88RYyH6K3eS1prTymS
wDpwAxHUVt3PCgWlb8gdReotJeOX32+SRYfBxkNdkVEB/Uzg2OhqOHNuUKh0eVX4
nqIxoUF/XwQ8kOubb9bWfe33yRB09qrt/4dQufUL3ymfPMXZLhAe/VheKzpVOYx5
05YWp7fTzYy1i2z+/JJyVCameZtcKDgSjoHSutebgIy5HPtHHRQWEtuUKocnJ8Wo
ilFdGS8zzmBxrb12ciI7i7HpqZ7wJlR0t4Ykv38SKS/SGkgE7HktSl9xe+Xc61qZ
g0D2QrNbtVks1/W9nSGia/jvZE5t92s8ftnyBfRZ6FT6rd2oReoq6/RbEICMdFYg
RNqc8vUtqevIj88LvMXLaTARCeMaKIwbPjeT1MXBacU7yMVAxBXL5NL2+jCc1oAr
vuW0a8rBrup2SBHebjN1xufaNbwvJHzfaxIQwT01vlHAhE0QQF2Q3bT1WTkQD+TT
b6ttg0c2E5Qvv8NzKgmzfuAbhp2MvqFwy7dScEIWzFU=
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgChinch.vhd
`protect end_protected