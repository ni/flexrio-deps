`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10GXbr/0ybS3CmweZF54Xqu32Puqrh4zc9PwKiB6yJ1VO
EXiufIOHmt8d8C87HIXb8+Cg9uHbJ19OOp+2Ulu9NxESIeCZCETypEml4ZEBBk7N
etu+PGyCU5MmpjXXPCfM1xJ6AccrUxY7fynPszCrICSUET+7Tib93QcQAs+UiqXn
4O8iVzCHvZP+Yba1nm1P1x9djHldAePKl2SLlECVTWBMnez3agZFx4jwXx5D532/
RC0wY3Y911uD/ky6KHBShD9r6dPpMl451MU4rhM/QJyK5nMC2i4ZAK7bjW0Sqfxi
DxKKwiZg9KXDq7MQvx2zZoF54DuS7/m8CuTK7OfnOy6UjrKEkG1YN7at7fZF7N6z
0A4vE/MaTXhBZhGPbX4LKOLOJfZ7Cpg9ydcW5VK2v7MkU14nHUreMBtxnhm4J1YS
aPnnl428VbwRHjDTqljqeQefg7Aom+SGd6h3H0jfnStj1pVXvGPDNOVFawvmXqCF
dsyIZ6kS7R7rL23mKmsqWHHB9NFpE9uWx3r+XckJtJ+XpyMnjPjqy9dImV7DUnWU
EWhMKA5IaRKb7uvhzHKwHFjCsGdoBwqestuRTNtUQGDqVrMGoMP3rs3DLPwzpcV4
ChimpxN253qALuaHuyd1YO1eIFCHuNpr9enLkiNJ8AT0q+6Pue0zMBRYTDzzN0UM
WvU3vQlBVMMarsInH9itatI7olhDzaePiLXTWo8gaggLL4TA399QLN7XweWi+WBe
9jalbrRDycWAcB/oWhDCGFSOKLK/VrNRq8sl94gpswzq2AkMGQSUXzWI0NWz0v4L
tg3MGMfjzk7d+wFxJr5+utxjNXyrKeJZQd77+K5Tbj2D0Ay2zdimgVZAcfQjXJH6
lMfvJ3zAVjVRQdZa7HxCiepTp/HvK00PpUij9ghlp7tssUg6pi7Pir0bt0hsfI1s
rbcSv4jJTJ/jaIBwyYvZxx7C+DnATY+0HmgL10EIx3E06v2UtpBBciAiw4IWQsX8
CRyNwAUCMg4G/LosnE0hZiv0vDFzqpAxj6/gJU7ky6cQG40gtPSIrnjKsPj0IqxA
ql4PVeo+qVsTOSKyU/SybGJJioQqhlvoc8eZlq0oGTNgumer9gpsh1W/2AQCvZa0
colgX/srOz6v5z0dhfXtqxApthF3J1bAVvGaRSx/6CUKccFcDNPQtPLa12rOaxUf
6vIq0qhH2AgIl/wzyItfg22CNVGM51UiUMZTtB2eGLEIDu1vaIj8uAo7FjU/LGKp
hsi0qqoY5HHc67+JCnlyS4Vb0WSp53BBL067aiXX74WJq3rTEFe9RsRZgL5NQXwY
YFhVS8oiWnrI6IGsQ+r7tgqhy5cuj5BZmj3KbvazzvkyW0aJCdWJ67BHsQnmawy+
AgUte0saapR6p37hkAs6mnAyvaSm9AybfBp43DTNOf0csVb0lYYQcV0pdedtAfr4
aIM6Lah+xYengG2xWy5JoU37Ql+EuRZMm9N6odoW+bmzR+8RCMQQJoGHjkQyYBwW
21qHN2JNzEMuQAK4KyHLFKOdaRcqR9H86F+G1pt8xfyRbkoSh5M5TM2D5fDJp0x/
JWiEl1PN9jVLvlPMs3Mv1VJD+FZuOzCiSOQqgyMrxLAGzGQ+OjVOEvn7ZnRI55i3
CdSrZuPydiASMmzRXTHC8woQBlspdm2ECv7H4G7f8C5EE/coOpnhs6g+D5pqN1Ut
xYqyelKxxnnxMX+eATeXIPlnUKBxlSqKOIljCYUOWhL2f6NJYbh2hGeL68MuC90e
4UO7MJuDrz3lZE8lX9l0WcvW0TaI7qy/aywIKdVb/N9xNzvMdosQFcZRqOfpRtQY
tIGK8mEXg11yu/XqGAmD0LUmJ5ZzHX6JmuiW+msA0e5z5eGAZHj93gPPmLaBJdnp
qizB6xJb2dXASscszLdFC3Q6d7k+KWoYyXAb4uDq7KRWxbW1nxEjYPQnkEU6VDEc
6/visB0FFJJlA3BZVz7qKmvUWlTuiGO3DMtYWGqG3xFc7SiucNeXPEyOPT3Sviy+
ly5NuMkb9SDZRw4j+i5mEQuLcbzfMI+6OUrDYvK11bgkkgakPDIxsTjfp5Prjnbm
7EU0xhJbKsSCW6StG7O3nnYyQ/ZUQg7KTUdx2AeP/OweRd+rbhMNfMKh58rtnxkC
8ZvyP8CLZcMAWKWYOE1VmbDNs4lpW8QBpfJrEcAiFZALt4mjaAdZjvvXzYrBW3wD
jVdsXNLn5iOBg9X59tR45uCq3LgE7WodpWNrLwUrAKRAevaur9GzQ/8yN3mfORqf
uVKlicpUEcCDgZdHK991lS0eCucz4pEqxD3Bc/f+XQVuIw4lteNmSMrheKpX1KLV
SIuTQ5Ue2w2iCi+jtlg0vzsyEDjfICqe+k375AXsvX5Rf6NuAARHTy82WfWvdQtO
96HiOyx+xJd0nHpWMunhKRXkQTISNuOXeN9gE1QIiGpCiC99H6r4ASzMq4fu36VW
mPAhMF8kfY18WF8wNoJV9iGTjL6xEapndMOb4NN90tvFswcT31AwdiSx5+4xeglh
lqP9vM3W2CGPxGhzDwZOs54xTxES+5/BuEsQ1XmRpeRpwvxuHrh9Ez0rYWkI2GcE
OtDc25GAZOn9sqPNFJ6YO8zeyqrJhAFLRlXvjrbEI4wkf1v+LL4b6pXfBwQqX6Zj
2N39wD7ctYNpaJoiZzRsDjCt1DSK/Fuj2wfmETom9h299KWNU6eKjEYC3ogexhDI
cSEEsrSXPwIA45rrdD9okow6fRRKkJkKtE4e76AfjiXQ2GvTARMZRXubzroMme6s
eU+foBfC64LHbFIjIHxYPr4J+s2MjPsVr2IwiKwBAQ8zHpdt/PpglMUa79QLvvMx
0VbHY9hQ5+HHO/cj8vaEr4MqMgHormkKAA6rXp+GvnI75fQQxKkMoniLaFpwJIv9
EcvAVMH/BBI6cq/wPwrb4mobz/KcLeGKr0lWfRcPGGE4+PeKH2lnQ16zg9tTnMA3
f+BG43hszNd60bzy9nOy7WxgsIY4Eu3kUPREjUkPZcLLJHoCyfDBOzyHwP+sAhmj
srICVwkVRB0LzRgZkYFlxL77rvy7iXNilFZMjt8xUA8430QyhsmPYqIIqf//rnmW
Hbt3q3xP4UN2GnNFCMpdxY0Z0Q51uApNA3TXLXNsAmJNokmR7x5RKZTcpw9eocgH
VQpw2OJv859FTTnAS/KSUy0f4T2aeIJUF9pzy3dkFUf2w0hraAn2T91nDRFSbiyv
GeLN0P3FIC4F7GT1p72dJNLsA4NrmxheONmX6IBssg8ssqMpPjknxNBdJxnYpubr
Ihcrg+lDQditXSt+eH8GGqVWmAjObS/C7GF73P4eNK0fwhbInsQiLQycFymbgiV2
eS7MKCRt3fRnjxINbMde3Kd6f4ktR0ol/02c2/N26xVg/OOBV80VGlK9O/3A6Hu3
MVV9Gf2MwrpGrzHIOowHzyacRAJTRV31RBMWPbyQqMLSGNGj8a+ZGm+LqBWb5vBV
BKsqomxmkxsuYomssiF2J49Rzp2hVjuXfq5mwMHGD+enCs5J89++ELb7ZtzCr/1F
sLFpe82XXN15JZ3owLFPWTjoQRIqb73eS9qANyikcSJHuZ54+SW/VZNMTxVjXG/U
FRTyNEHYWvrOSSwgAUtLW5Ag30l0itSOBafdQtqPDCZdlz6QjDrnZQDTnmpFRtj/
pbKfeTlJdUaAW6hLUVK1TfS9+58rgoVdNakqdYKpKnbpFUKzTLv6HRZjHq11jE/x
oz8GQ0pf6I3mRIc3dHE6tBt7rGZ5MGdTYapPFN+71X6vU8Ec75Cr2oFiJ7o7pl8r
jcL0lJ2a9dOsdyC8jGryfyoIRIgHxmsUfOSB/3dNkEA3FDOPTgimpj7idjxhQwc8
TyXIoGeGBFyysLKN4XZ5EyUr1EUxJRiIlC0Ik7zPEXlY24MqGYOaCY03pAWhLV4u
+I79mYfcu6nQvy2dYD8lb74xQzFgc3FbbeJtnIaf6BKu81m1lvaNpKO6SQpCmJeD
VKM8zFRmBiSWr8t+1hGmQyXkCPIJ+v/Bmy5NPfl5Y6clhVoBwAz0PD5nxVKkF+f1
KCeswCVNTh9TT7SzApnI6NcKdVsj1QgrafVUZWOkOtVXYZvvQGuBhMJ5n7c2OvYC
Qsy3vqvRpb3Bw24ks7gX64FLkknq/iTjdIFoOJ/hrt1e7CWlRIyH3oNuxFqlpfGv
F8s87uP33vaU8dnxVjzDorG8WNSAMIMGOVNvHO7ATuNmv5Vl5g6BAFu/JBU1YxMt
NzJi0rZkpFfCH+XjyFwigRxqN3jvqEFBAce3jhGB9x0VWMEUQrMB/Wtmp+ALRpcI
hciEuEKBdiNNXLy2aAl6YiTlbJHsG0LrmBFCh9rXh9LVGFM8OiWCaG9M7kuLEHrc
Sm+ELD+F61ON6rLu3LKY07ptA+nbi0u3ZQUFJl0dzQE5fVjf/zUpOZgmAMGKHtCM
GfT0+UN6Nplr3UyLG22tUTtH1h5N0p9Sc7iEhwezGjm3ht+rWc2omHFkvq6I8ost
VX6KVkDS1EMmQXhqbiWRBjhds3o/1slhsN42BqjyEjB3A8M+jxzaKhFipQnxvl3+
XPZOL6PtUmQFfa31MLM3rYWERxeU6Yal9ThVfuHIWS7weXirZOOxJL4jWTNTnMDe
xdhQF5529Vxyji2vREkJaufXQURfrf4UF5yom1A6Z4o9xupKyLp8joWMWfIij3vG
IAgCOSMlvsgQJa6RSKx1Sn0etdGZqQRm8XoUggKZmwluY5kriiLxUsOeomG3sWIP
B7FQlyXqsGxFyUegPhwnlVGVxug5JJLxmPy6fUC6eoRIfNRzQHRDY5nZm7YtdCLK
/Ab8y62Cx8uWCLmosS5T2wk1pF8LtZzwUykT5J5yAK39X5COOz5mrXSDd6elJTra
GBN2Ho09MlYOO4kt8rdDg+gWMqu3x0wiRhS4Jh81xasu/h1cwZehiDsvsRONxIAA
s8V2w+BHhAWdtFqp4n42M8t55peM6bpvAAscvGbCYST2/x/n+U82wjbTnpuxhY1/
pI8T393MUR32Klr8euUDw+FIkzyviJ0Gr5pFki1ilKD/5HjwclE019MUIL8sWscq
zYtyOQjpnQjy1EhLobtD4i/Vjug1/w663eTXQsx6Zq/FpL0BmIuDWHLnmw8DmY4y
khlD/cD/kBcvgi6IpMVyepHMRorTIBfM1yGzExGACrhjNr7nY93oS7k5cuX7yvBN
kENPL2fkJ4TJBvLqCnCKZ8l76xq0FXZROXQfxevCaX4Uq/COr/uMzakBFBn9g3Al
eSU13KQ2mc2ZKNmRkxZweap5dksfdTYr+A46hXyKt/APjxV+/dq8GYYi0sPKrDTL
BFnvyJo3DwMmQKnImG7yWOS5pwS7FLuR0LrJwXXsWFUsfl1EWN0rTe6i8domyAsr
jY+xNYSW8F0vJniN/P5PPw0ktIx/+nPZh13GoF0Rd20fY8IZijUp0u0amJm7mg3f
sqQo+0sAXKnHL4Ul6FnMe96D8NqYPAkot5zyO4LT3i27Tt3ZG8KFNOpUXcnFRaH6
DcpeOVf/I9jFNO8cC2aH+i4OtpCZru/DwzIkiafN3W2fsuKdnAhHXauAA9UlzyB4
saeAEU5jvM5gd2ck/K6sneq73ayBRIsOekPbgRFDd29RhwaMxhmgmCyJAqjXlSv/
CckfNjP6AVF3Ziqx/vW1ZFwV0CBUpQ2fOJZ7NVQDwDUXGsN8jyAMM4RPvI4at1kF
f73BxYaEgAKObEqsPjANBCXmpD+9gp2szqQn5siwLr91zN1Rnx9yofEXd1W7eUoJ
/T8W8IKTDZi2z0QWO4BftFRWFopWs1fzYiia5fJCq7hYmdQnfKU0DIjlqtrbsP0u
rjMXZiNO01NX/0ORid9kwVLzkS4WLv/dKd1lVunhUMMlHKUTXGDXut3zkOTC0/oN
vNF6BWepgWIdLFwe9UZY/0XHlrJBFT1b9Sw8zc65jK2JbhHIPDq1o1lC+P5kR7vJ
2m3FwYovsX1UzGxTPIiMibRJt0oW7H/XzbCMcZnhgVKU6ycgBnCXIkRirhnvlLls
J3VHuh7xS7V6sFpsz+cK8pVnoFi7JmKII7eeL7zNiz8ndHZj5e3Ov/FrAb7kzgEx
OAjNa4IlHrqa8zR70VMEjTwkQ5zpsIu0bpRyrd1xtLsFHoUKFOt1Wbn0lxUU62hP
oXh+HYqKVBhSv6anJKfVGb9mekEHjvwnqc/uAM6TGX1BHFC4604nkJ+xES3Sfb/w
oY9lactarU0yTkqAaKPtPseHY6/h0p+LJHhtxxtmNoXhFtDuzrrdrbCAjEye0Zmg
uFZH3OiOzhqQSXvuYKICj7FpRznQv6OuKkg8WGqOMEWbqpApMz9+OharG7AJdlVy
r0A/QfIKf5h+xmfqkx6H/7sBhVQKQD+91Jog45VHSDAa76o+KA0qgEtJ4bOkfp0y
WUOBAYxQMpV/8CJ+7ypSJ3UVMTekHLIhxO/WZcVMGpsrXA3ctSWq5SLkrBaKOJld
mZdPt4PtQ9rlVY0I23t4RMCwzVAIoZCOskfMs/41cLWr8q4Z+H+c9BnO0Thcbt5R
UtLuvg+gPOLDeL0JkDIjEhxXSp8tMv9GqUAomoYbZOCvgyzzhaK55F+FqBBdBQVz
i1iT4cWvIk9yNfKmx5423/Lp1p+lZ3+vman/xivNDb3D0NNy068WjBaeuGazMXpy
9TEJEOKC2k0jGmud4qqmPMVoiFSA8LooLxBPQzAri1NxELh0K0X09oC+NzRxRmJu
HfMhY7U1OwnpkVScgf4pKlSlmt5+cYxH16qpvSESZ9xHEHCDQ3eLKs44jtnsqQjV
BX0ftvZ06vvalFtPGxN34f9FFvTh2ORtlAq6gDfQ5t68K4An+C4lrfWi0S+h7n3i
MP46E2fZiQC5D9xWGLRP4WoUOC2DiI4SJKOyGZXVccheTOEXyzXFaLOJpRKQvAPJ
EXm5e88cg96lkxybX43LcKFgSaCRR03oem0ItwcIR+d2LeA4KkFmcd6NeBq6HoPS
zD58HL0XmecnqaF7vG4dyAd3oIYtK9MEjuCS+tLZJAbyE+d/QDPucw33KNgCHb7B
E8cUC/7bwNSxJsNioJmelCtWqaviVCsNTz09wDUAi2Ua62Tb0aeCMW/K8ya18r3g
m4SttI14u/YMDMotFkeN39OiNOm5UDjjsb3pIZWKvDx8GvrTUJb9sBshSrgPiLby
Xp864bBQ9Aygd5p58m7wy7Z9mC2p3FEdXf/tYyjnn4SrJefoUtM2TverTPEO/o37
ShEIDqscNcERZu2it/DgGwwMuH0j13gA2vHuoT+vwEmsET/2/atsgpWQlBOTAyF2
wXgioq9KttvYBd4UJlblvnvDF1hKCnCYlJKp5nNiCU94q6cnZxN2kRT9qnP7h28j
bGRbqhg/TLSvnK0xw8lIU02SDFHfwR12Ljlc+F2oDTGBzpjNUDHW03Y/bj7dmk/K
rznDKSOP99bUWjiyI0VUfO14Sq3FiUarYigN7/CQRmoZYJQ9vJv6gJnchbwDHnpY
eLYaSzSC7DYWZZZV9/c+FaYUp7CtntOdoH0EF4xkPiCmXJKykMIVnTmzxFdDivkm
vFnPccyP1aYKa+OO+Ox7EhswKQD8hHrlM3LUo64/pXrzA1Mr5mRaTw1XlwFaWroL
Kj4XK23wD2kvMpDGatMGPX1E2U00raueLXha5JMYdPWkX+h/18R9CUY5c+qzb8BZ
UQjIDgaVV/60jP/EZ4OugTUxrhmNZSvASFTyKRIQuxomY+FYOFguMw1roDb8T6fj
DHXBVxuWIbHSqaLcoU2yNs0DHCG8AUHULMHxflcBU86ZHCvP9/yYRv2l1rUeRl5e
Ucwm5dbhP7acY32PDrSFLPikw2lV9XIgBiazukZK+d1iyNALiMPpdk7nT7Lch0N+
jPqE1d160JK/I665eIie4ABX84fSrNx+eeuHZ1Ng/oenoQKq6QJM7FNJ/2rwXJKx
X63eC5AFpC4WmiTEDtlfU8bwE+qPO3M2qw/9PQTg9OgR01MF+zLrpWsXaWTOWKQH
n00IV7b+SRYtWKFYt2ved0sWBrWVSOuZ7He/GXuDZrPMp/O9vDxW197wuu/dctP5
v5MFvOeJjH7RBXPAqX4PHfc2HNQsaqk7mzMSvDhgtI/4eUs1KSZLzwsSdpBdNtQF
dpy6SlmsHNPmDUkFqzCxi+WSMuJZVzJb5nUtJ8TLddzGa8Tkgs5LFi+xMsc1YbJ0
jgO1KLteR5N9PS7/EMqP3srB5kTYNDVw3t5/U3Zvt38D3H2DUDmNqOFM7SB+NwFV
zzmhLYIihZTiWmifBZBqko0jaqdcC8t53qAos02Uz9MCUGpY/jOzQIb2z+bwq4l5
KS4OBB0pQw6dARY3jrq+b7AIqUaXmPqRL0LTrGe/f2AIE4MtvYg2JTtAyroNIke7
uIJ/m8lAef8/foNRitryEdGw9+5P9lpjX10xwcylWKKcbbtvmx5HZlfUCfI7GLVe
fPY5yeFtJISvsbm2KrzFp7gdPyAVyAUdDG4a22LAKsZSFRHuVjKrN9mriSi3W/9u
AWTEZabfVoL8cAjh6TBbdFqdml255O5wtytfKNGB49gTrH/OItnS95JheOANQ4nh
Z/BWgQTRoyEEpJTiddi0QR4Yo16ugBSt4iuCIkWfIz/QByjP5PYB897a3R3kTcAn
vIrLMId7ENFSOCKuH7v+ofhMmxvuwamXvJB0eUzMeSHPQMCqzoI1njn9pw4t0LvW
FEZHU5H+jUCEs1jrDYkwR7XkGowm+8qhQ1BPEJk7ZIy8ghHH60kVXT+cyuuXyOdk
o32WiRtOiYyIer37UaiThGh1t7myMN/irYRaVEaLgr15dbbB6syA2Ipq5tQrjAMS
1QY8V/nyQmuO/nSdqpXg+Oz0z6xA5wen+zqcTCKxdleolx021ejWT41jXZU29Ums
wp479mq/WIZbYt4zU047iaOE83ucwv/dZ9UOduyspcb363HagzPM9naAhvbyAM3P
qYGnTBrNGRiogahgdj+duNRyXW02/vmN8l5fyxRJBsRSyL7cow9JagvEg1wTSrOj
E8mQmu9pRq6vcHadplFvmbDfIGNfGWBww75+z6BHFpPwgIka55CvPJg3H9hc7bhy
zhHCz/Le/0BH00FXW1ifl7lGhJeDKFrDMSehazHN+Ok6o2/wlzmayNnLlupErhoQ
fB1/dYD7nKQ7fF66SebfIUnlR8MuaZ7x/wAYD07vL7o7WXb+1Lcvk5zH8q4BLgM+
J3INu3qiD1LH9v2BQ0Kj04qGWY8Xr2qrh/UoS6Oy/d+cBG8+g5RwykDjvxCg8owW
ooHuhjwhnacbAqlRRGrCNOMmj47n2WIgTYYRP8tjpE1qeRLvDtgXnQe19Z3r8JGF
fkEUenRfjtYzDbjmej7SoiFk/sAJvhrYeeJ085LUX5iGp3UQNhzeB5aQXDKlTZLz
C429iNZGDwFzTIbhcima6aokMpHcYhsAL8zzbcD8Xe9XS5xoRABh91JWjw0Ldggi
KLPgdrI5EI4sSdtgJOWePwFuQiSr/swS/BlWUGHjfv5ZD+j+krkrDtnLNy3Z0C+V
bSl9A97W/gXcIYDlkKkmKyiORiba5rUZcGHwpy8AZGceArjFO0oucNGesMLTsAwb
H7JYK+OZBMWiPzUdZZfpm5FvmuK76QI8jRjRhcSAehlEXpwnSQU2i4txuMb+c7tc
4FNrkZ02Xkldv9Y80NrmDumIDk8hY7kW7U588jgDiI0WkeLyUhJGavVPOl1g1O6K
ggjmOMgR4seLJxVqSUBGnsg2DITEmoV/F4qTUhNxUtIm2LdcRDZ6S/K2DMqbs2Eg
Fof3rqnMl6tHRketMoLn9PNzJJNVEMh9I13f5tvtlMBgn3PmDRrUsnHGPsfwb4md
aq477zX7B586U5o84Ts9juHRmHhBNT71NGf4yWigtBcpKK7mfKQ6uv3itGM+EC5Q
H0n41YuavyF9sC2oVOfi4Iy2q73wNwDN9dBa38Aqm2yGPgCbZQ4j85PMRC+7E2Dk
zM+nMcerkkjNRvYO/e6aAMR/NBuUjDOaTYC70BDbLDA1VzfkhM2fk04oy9nsvlpJ
wUSd8EL7mlRYhhea3e50wLF/NxgLw3fwKWX92iFbRAUQPPhNXetvxExm2YoE5N0R
gJQmgiuJFSLwvWEQZ9ITUuLUFw5/kL7VKsRslnRyjMXE8z4Ds3P3yWTHeAacAWL3
dXTjSw1zoPicPdzmHxoAGueQd6xl+vUWVoPahxnX+Fu0QpWI3u9alO9Q2OF5bIgJ
1j9kxoJHTlI9tHgUOy5l12DOjMlNL6HzMJ8t7tefjA/tcLeZdJHxObsRxXkqUTDo
FxhWUC7utJcREwSEjVtZKI3/qz+TBZ/ayS0mfgG1UpKSjBeVAfqQqsgeejc63VXV
E/Hm0NGevzASDmdu4ekIILJZKMd9iLley6T/6dCzqRfhx53ablMWUv2foV5tl4tM
SZhNfhy0wGstqnNRZf6qceDfQXieX93kZzn7KQZkam927gtzRrv9JL3hMoZgXHbb
fbEB8kv4+Om2HPDF7Zh51LgBXjYRLK1DE6jTc1XYkwNVi1/vICK0AmgleJCE9jvf
aFW+Hb4NeJ3ecjFzuR7scGFhyPSiIb54tR3eanM+8OnbYxmQr3u3kC3+eupcclpP
hHDrqdytoezSRpn1tVth3bhL913jQ0Z3QZ8T8L3Pi66XgUEgjOmjJc/YuAKkiAId
AUZHEfadg2j9NMABF2OO+Wetax6iFAqjClIyYLEAQyiOp/K57n3U6EFvFuQo4a1M
hBbr7TqIK2f8qEKOeHgu68Vr2wALYL2sI86WDQekWwK/CH4NDC6udWGCaXlHngQ9
N1P/6tAfCDzVfV6M+NgcqaFbPy/HTJuTD9aBpibiEV/dqCqmF1MhOVMmF6VS7F7E
a7yFOePjJhydv9Y5eeETwtBQThaZOHRjwZB+2cA6M1t83KSAVWvP0HpARGXiYUD/
MnOBMWPHtxMc1Zrzm7F/SHoWjuFQIgCmwLXWV7AKKiyuy3+Xhnwdqw+CmU5zT8d1
T5/GrMBbUGGm/SK3yXkEcGHD8WPoyn/WJCCAzopmQ3POnGICI/I8KHGp5ykgpK9V
hQLAJwx7LS1AaWVQo7QQyqf6YYzpVhKvf6a31gwoA8bq39RlDIGyXwXaZ+cdj6yr
EKmUpQdjugYiPQ2l0gYOzfD322B2F7OkBh6OFHzd6XKlvi4cWgg9cyhk8xlhLjVM
FprexrNNHqRRW68GKL5o+dk8BI2LM2pne7jbYrvfY4k6DSWEkXt7qcY5leqxxnly
kGPjAygbfjUX/MJ1eCMDAyup1PWa2hJvLlr5gqWBq1RShAq2cTFXsoyhuwS8DAES
tOWRt+KaBjJgMk1UB3WfNdVF6yhbil4Zl4Zj8jWT333xJrjM4WeKiCvjVzYAWBf3
f6Fkde/1Gd02QMcEhMAA9vLpc8PB6QOetWjsviDf/hX8FD+x397XLzlAu+wz1R1a
mlpByg7jvPVQWMdP9r7+UzwgDINARQSYAs/0ZQ4/be14Zudi26oJSIISpPEG1HKl
+ORkLcUaWpXIVmtfGcb1/tqTfjKaC02ciEt16JY6Hx+c/eiK4IfVaqnZ6ua4HZ5B
FPL6WdcZyCQ19ZyOnEergiY77ogt8EFhYrNisUkUsiIC6n4XZi0U+JxJb/tDrNEE
2n6+aOxFDvKn2WmzpxTkSceFa8n7yQsLtv4PkWFWIloRLpj3jWmoMqR5Q1tERsLq
6w7KXLDHL2mhOCHRM/HAloamrLWiuyHlzhgC1NqB4I0iRQ27SOWGUDEkVbWXg4l7
bd+9yvT7r16rxtceUPtDYvhy3DqkpCRmxR9rjjw0I6+RPH+ekd2snAvK8v4HSO0p
lc4JSGOIqDvP5o5sPZ/VmUBVXwmf86Isyb1lhMmfea06sjc5dkvec5vXM7nvDPg+
J0VYx9NE+7YfGSE74+w0YxwvgpNacLrSIaQeBEB6TViJ8jffUDJiWnOuCzB8//ex
z9JR0EQ5tLKCFPtAqkiCq+/s030tfdUQOoJNC9XMC4Y7craFd3YEN8z0xkPxNhY4
3c5X/JM1w/DhUeSY/J8xTM/e5/rv1iTAGzluLFqXVJu7NtkYqPagGQ0paZjAKHzv
mjpPK9YxTQnBu+/QZQfQkl0vrwxNMiCOces9d+X81d9u5SnqI7jAw6wQMPUDVOMU
ucpDulgMawsH5uLo3pXfBgz0ZtJyIZWfPm/15P/P3x54ZdDdvvaKyJb6dBt0qsW1
jwR5mpVv5MkfU6de7g6qF8iWkCqoc0X5QidGysQR9Cxh7F3Bsbc0z2OBNaMUgq2I
JOauqd/kpaIWXzTUb5evDRfPYXQjpY5rkZLFrrsvc/Tv2KWwJpsbRHyXhCxRh3ku
PvdSZU7XP45kMrKU5gvs99tU3wCHjBtLQFZDe00OxaC0g3y119HWCWoipjjp1q9b
r1ZNG4kJ96Ptb92C8601TNzObpo3QwsDNb2+YKLuenlzs9qSu5Uu5wgqvh9e8SKW
2SAIkHM7OU+LpBh11HB7BD5JNmb+OVZOOUwbiaWJopB4pSpHF2b4hoTXLX/AXoLL
MnSyyDi2ojtf5u35TppJN113B1JrCk643uTvlSoesP5hGO+CWHOAh0xXd+KKoWCA
IuWFSZm6bagffERnKhXdHsib+FxIrKrzjt9MGplG+/6mS3S3nCZH4cfrpmh/JNoA
1Ajtvk1rMlNPf31XrUuTgIRN6ljjUgqq4i1pExHaBZQ6NFvEXXcBoAY9v3ggn3lS
fnUvmTl5aOLmgPTuN3GEG8BD2F8HKuDGMaL2kUv1IQ+Keqj8OpCyvP3g4N585vIW
tszzstbx9jk2Nai53XzjIQi2qeJU1bYco7tTsJSgCXQYalidDqDdMXVatkcQPp/7
YGNeG0CyQbu56i7qLjhIiqtYKZsf0q98nC3KV1/kFHmg2t6V/vLSq8UfwP1rLjJm
BYvCy1RHalNcLJw1WbobkdPTS/7PpacRyuqueJLQtnuVXmpgMc0GDNChNmzRhJpL
dBeviaCoNZtjGshnnRop8ZXOPXdSdT06bQUt8Y/+TLOKfXWWEOyVebxpor5MVxKr
5WnPslT6AOczdSqYcsi9Uv1naUiZLmxK5jdBG5jzsNTGKIdi+15KZRnXe4C49t24
JuW6qX5eJA2ApA1tvAPJpfqtXk3WpY0WehQm31CWbPN8H+oFnQtiIYPLT/0BFd5c
bwpWaRL5Pw6PRuZoyVNR1tCqiPl8ZqZmeAy9ktNWYj05oz3SqI4DmH1n/xWzexWq
JJ/WY32kFFKwUbx8FgbwG7v+2WYg9ymXk9/+BBUCeo4OjJQph035r4wqNxeGz2fD
zgUQYE8RalySb38sl1Ain9T1oUZGAlOhl7wkqwdThVDE/YKQWB56Juh1Nq8TpEg1
4MVRisQf8q1Y407l+p/0yktsIwPgg2Vj7OYkCvkSYmIRoaciYijSu6hDgMsUckZV
dWGPrHgnZHnLIrRuxwvurpB0U37lrqLebVSB6mrh9SkY87Nl2aUJRQgAQqzBr+pX
vorAtJ0+BvvMDUaWnLCJPgwJi+tsZZq214Wak75ed+yXu/Xmnz+nfcOjPasvGGeM
cBKuOvQF0XgzZKrExeHhoRHY5e08YXKSWx3d9oWUpdqL9nGCmnLFLmLde2ogrU8I
LqpCK5hjRm2hIxAcc2QxQJ92utAhrdmj4rERRBTlCFk02XYVpY66gi6eyU/aDOhD
qJG1VokHFehqiAOjduXaEQi2hC06xupgJEUo75JTaU9W5L4Hq9ZaQP9KzfNSIy/y
mI6F4Hds5csXihMRDzgv8zSWudTSF3ivmsaW5Wfx1Np13enCXGiTTEWgSCEvE7YB
/6BtV8x1hUWFDmgwFDeB5lZSOHEpVqt1Z0uf8M/vz+ODvN4WZY2LbbaTXX+coJl5
k7052lANIMbl0WQtjmqIBKpV3m39V5hkGXUQyS37RX9ADNRnWiLyVKFt49HzJGgm
UIXocWlbKCw7nepOm4SM9nwhB8LfkDdW+yVDVBaRRbazecUS4qAI2tiijjzCVQRO
/UFXosn6CcP9Ps9l372APRjT+bQUksO/qT3PeyhMsYlDA6uUYLZNi7qwOC6SAzV7
Xl3ka6WrnNrG7PXa0Do3ZC8dyJtqh1PgSpuul+KMJoCNNoqwEmjla52+JomS9FBu
WcBdtqDWmblM53358eXyUszkhsRG5zPQVjAmIEGjjEeC5Q2RFMbnooxApDHlwQ3x
buDSG+8r2B0sB9m6vcYELT6SbBofp/0nhXvwXys1xf4/P00Jf4+D8XxoHiSELHR+
g5AbS3HeCc6bF+4RSaMKf9MpXHsRy/u3os4s0jbRvspaqNbavTQq2Bl6UUPfr7w8
oEHJBP4V13rZqWxhBH59JtfchlXAFYh9hv5cVQ7LnnftxDZOwElB5MdunvAtbjwu
TAtaLFf4lmVsTwHukZ6yC507X27XjhGhLFhEcxuFiArZGnNUqUG1l+DQNaLohWzL
gTgNIIBx7r0yKWfZs2Kg2rDhtJQ/mJ0rAkXc+In/J/78/Et5EvqPaLLcQbCAWc9t
p8YVePJPCcWJphwvS42BM9BdAoF0m1/JUxHzuJvs23EtgDozaVkLwNSurGA9s4ka
PBWvDrizvwvN069xbc6Tp/DKj48afB1IFiX2GD3SRH0f3SABu00gx/gQAzP6NUWT
bK5rhDRTvr5ft/Vz96YrhUE5taD11eeR0IO+8hKViogW3iiRf6q8+iivvJX1GmGF
SW9mz7jnIl+YmLXHop1PIyf0vL3SiYemhmdwaFBWChwI2/Pq0SQjtk5u31ibYvWK
2+nZ0jDAoWvu9XNON5C3Y7k6Hy+gCgmwjy8Pp17FafAiuqm+g7WwcIfE9k3wVIuQ
KseE5BacBXZvKRYfGRVsaHHn9A9lM1Nmg5/h14U5yjR52/8PVOnO3x8P9cW9Z9rl
OElhTPvBNXBWsKGbfG+D7P3q2mV4gUzt1HuGt43QyScASYKS6v2zu3kRo6eqsvRf
Oa78jIopAVTnFtB9cQlAnHmhnAo9iPAi/rZkKkeo4uLnzITRLmqcvEcXeSS3uxGj
1fBCzfklZDdSZzMynixipFvN8E7sI0/iBZ2s4PyvzddcWtps/bHx3Qn3TqdeHUDS
QTk+2pX5z4mf7JaMOkw3nf8H1GC1sAkzzTk11qu/Pak+k8Cv2GSvdJP/hXr/xG+8
h0jQUCXEDV/vATXsRHuE/4fXfhx1uCETgxU8UoxwFkHK9STix/ObYmmf2OnMg2y8
1SdxxpRgJ5IZZes3PmUoEJz5w7/ukgLQ+wXqLXTLVwbUzJQqE7T7yLti1WEF/nS5
iAjFp7+z80M5tedEoVD8Jmmwm0XsXtRqJrYFk07ah9a6X9nHVqpR/4QUrRArRoY7
Asb1Agnf4uZafFdr8lb9/Zh5vHz+0n2q3yVJiwP6CUbVaa1Wa4Ii7gvnF2qMt9EW
8IeEFs5pirhKkiqHYI8/cKrjCteRo1QCYD99dj9EPljN8wSKZqBq6y7fKXpjrVRT
3XG0eEqVjHGk2j8guhT8mhIHAXNc1c87yeT1b61qTmVPXdNeiNnWXuze9RuwqVLS
LaKd/y0TW+B+Q+ZknG+FRsYTPCcOBZ8OzZERTiJcyF4edNR/uUfRlStzfpysuJBO
u5b8QKDuSjwkIDf2MC4iRLE8oWKq3Z2zyPvL0JtlpndYRHweMIClFSRj+WWtoDeP
CQoXaUpncBZ2dFIyZxgBJBjgylj0vB65Pv8w9QRb+IbZJzloDlzQzhxc+fdZcX7f
cmpdsV9CHv3CHUD2rOUGtHFpKH7w3DDH3dhxF4v/z5MXMudAxZBfGwzhXKA7O66x
afFit1iE12F0bgn3Ps5Yvz/7tEz1uZxa6+u4YRYEcAyzAyco8TbB4tkGLNUyDmxL
JN0mjdyc5TGLXf1E0NIlKnh2VdETKwgn465h4qZo+LZwpfpmeQQRP+rUB/O8t5N0
aKg6QTvyop7wahJJ6iHGcEVzCTcU4/lTKALVp9HAraAcz9TiU2UgdGVPVWNmdfqg
DmT1juLXZPGCNB/+BUkd9Nqm96a5mNgOwCN5c+eMm2z6l+TePR68glinfHpRMFoQ
roh4rcbL39ClXq7Iw91mc64dn9NNCa7NGFVUxUrn65GdZHJrKVh7B4Os7pN1XBgR
ueyBZtm8DMtw30bi+RFJ5RLHbx9qU4iF0jpFbhM0pBTYsDZKXQiv6VUnup3qQEmc
XQl5CU0YsD929ADQyo+zq24U8fOUMShknwQaVIbzto1yLQrBuYnbgY6R0WEgC8w8
5rLKT3U83f28uqlB04HBfKI1FPO+6JcBHWAhnekMg2spQJ8XpLdgNpjlqA+n4kPt
Pgp6tvoKmuP3ohlW+ionza6C1DJsCaDHCHMvKtApJ30rtvdDExkfGOUZTcIwaXhX
JyJXpdaMxIleRALA7FXSErbBmoX6vDaiSeuWKVUYppoWzqAQLTL9MXWPiHML+uza
rrFCQ/qPiFB2/Jax0BIM1jxX7bCIzPNZXZs1A6l0KXCM2N1+pbqlrGuihuPwKyOb
ixFiBmcoJfgrst5Q1tD9SEVpCbeyZndRngAJwJv/VTDB6HYOYgwpy5uhPJwET6As
WiMWoFxt0jWl0fox4CEI4+ZjrHjjfFzFl6Kzp6ecz5AbCAX05UmoruYoj7m5Ln3l
rAKatvZ5VolF8myrys2FbXxEdwBQxwe6Ha9R3d2tDChl72T/pGeVMur0pGY6AZHs
txHXASJOvFLQzYimlYRn04gv+S79TXJ5eFU1P6V1P5XyDSa9gX/Hnr/Em9wti+uS
WaHacoYX2/qU6iTffO89RWLmqYgFCx5SXS6wiL04B3kVRrIqh/o97xk5USaYu/3b
+6hDsPoR4QzEke7czSjMjztnXWPkN/dF1C4QcoD6rpqhmdPRUeJmU8kDpm8XPMar
cCYjBndNLWYODTvdjVxCiIrEiEy4/Dv6mMGcU9eumrvCslY0+Z0e7PDfCjmC/daQ
LNX0FTsAnEC9TldGA28APuXxGTN5jtmYBo+yHg6fZSyoPWi0H07Ci7PXxccq0Ie9
YQLeBblxYMCGoEaBZnM/LAKLIzSFQtWAAd1fRSN2aZGDYUbaPzuhr41w7xH90Ho9
JRQR7xhHQVpdAUTj+QqXMH/4F2cjqhDVriHlDAE7B0A5Rc33Bg9mzuiKnaTzPxAi
qqUNDk6rePAvBgeLpQHsJAni7xg0mwCp6V6gjZv/iVCd2WUFTuQ8dXCTUV1u8t/T
XvxfJD6saud7H3XMR6qpXdPcjpydD4+sCgvklg7z4u19JbgAkEm09/qexuAGrZpX
2Y4WruNuo9FxpM1zw5tXt3K0ctJC+omEIoAHll/R2JF1ukZsRgtgKs6BNeCKbX+2
Xx6Bq1b5ZhBZp5dXsqpwZ3HgMw6VeAis9ZT3wTC37BVpJndlVS+bDvXTsdcwIxo3
2eqV/We8IVjW9YppnIZKQaTFFhHEzgGkS50wxqNogTQRp5z2st2WS9HLrkMk9EVj
KeqmGXghiRxUyV9vWU/qUve13jV4ApLdycJsOAqe9guuC7PW4X0xpUGYlAHgNoks
YXT0I8zDRfth5KNGXUR0zptO6lmm+rkOFLvepSq5nQniI9AeoHwBOtd/S2P2KHGl
OAv05yxWnooMGnCKGS7lv8Pjyi87xXvfgxTORAPbQITSbMBJKCccRJUoactnypaJ
geIU4M+Mdl/p4T7B/yP4ZMlY/LNwN6uKCY0dKw+jCvpmAhxsnY8fLouaIQTbZNiL
2MBQjZeDU0Ag/hVPUmpjz0jM3oE2hMRIba2Y+aiH90KcT0O2t2t7W2/ghx0RUisE
aZcfK1HztWO9nHHDH+thKprkOM9oXjHLo4RIMNk4rsnSzysUPMgamqefJZOgf+Sw
7ClcocdROfxW4f3baff7VLfykd7/UAM1imlVwmgV7lB5Ake+ERtlsyUSmwDmZb7e
1rNWOkuuB4NAHcsXYcwx8X2b8WZN8WkVZsKWiWRm2Rffjb4q3TU/tZG4fuGIMTgT
fLjSUSdKD6pON5rxLbWOEqK+KVLj5KhjoaBLmwQBX+bEPpqSngPDv/eVyf/uDKFs
SrHfhPtDD3HWdhDRYXB69YtaqxbqdH+Dv05B8qvCTc2M4ox49uBafruoJz1F8Bck
lrDVbxtPs4aSePadCjuifqyJ0C2zPeKomynDR6Ci0eY9IhbB8EQdipNgcdWrVa+c
gqfbwtLKZ3SmUggSPiiWzJG6atpfIYaOmHVEFwNEOEI7VqpuTqr0bwQEHTetx8+p
JqkUiatADgIgTv9d9vXwv7vkp5Fj4coREgArfiMpMaQ5kjFKeuRgABj3x4kdSTLg
KqQXf40SFxyFXDvDTjeSiBBemsao9EmN7bA4yCTrRVHLeYpyztCfR7KRK7jtpcmb
7W+203+GihV4iM/tdQxLSH9pmpanua4Hc0oYMfBQjx+70dyjem6j8ovKBUaJDBkW
StLDqX2TleBFw2NY41v8AE1rx7zK9JGE1zK5xkUnZcPkhCceYRB9/1sk3pWIMq0d
9Fr1BQwuouQJFZwoQaA8taevGPf3LvgqUA1uzre1DK0PQY63/u5lV7T0ZbdrQNue
rnH8rpGaN3Z7jxNJGKw5OluiJenHGYVHyie8gkIx49gt5FD/uGUXkZXczxMu3uD7
6WWkFoZF6gkrrTVtXYamOvjFqANy/l3Gf3D2Ne54hg8k2XvDKoxuKVZDoABVtVOW
HMh4FXzEfURPxiG/kFN4AI7a0t+c2RjrZBJENJ49vtK4RZuLupbHx0bAD8pPHYZH
o0tJaTSbBpcov87F0NWNbJ/RhuLqbcKwKTh97YqyXGEVq8Lg8WS2o87loXQYT7Lx
T+bGR/Yl3AHhZ+fs0Cw/pBkhSj8cH64TgHbja0LVD3J5lhzw9I9VO0ysN2CFQBzh
E408NN1SU2eFhbPPwD6uM/sFnlxwxBJeZtyQeG5NQzd2AL2/gI5/pP+LyxxsK/kN
30P6uWlp2FaRuQQ4hPA10LwGMglyUzNc3tBrpzIc0XDsz3UEVf3hI3CptpXq7ER8
UOXi/q1QhrUpMZgYLXpf7iF5J1xZNf6VCnFBCeQNio+MsqFNyQkmDxTOI+5hrPpW
x8yksgagqh8ugbcESTGGHKEtTs+6DkJDIDIvwyJNhftLo+u7BNk2g9MOJ1hwWJbH
wNTqirOfyljRvJ23I0bpVrtkPk32P+N6KGzCcY8ZxZjEXNIbR7uEXQ6NLr1nzKMC
0/NMkV1nNa11J7zy7yfDo8hzDr4RazmDOxBAW1sv5WLXG76+B+4XhW/qrUjnjSgG
CTFxJLpNHxZuVTifGHChuBpvKWghAxSFvKZoTqmPYzTKScIH81ntK9Gzo4kltRPT
CfcfNLKrqVb/oVxHFo+Q9mOFY3hn9cSKqGlK5JTOHbuYry6HiWS2fUXslWya2wGA
xsMWUn/kSFQbf/q0yjTBpiGXELMPuJ7OwbGp1VgLhXoL/AWGgRSR+E2REUKZ/NjQ
dskQMGmoXSof86WzQCcvnbHKC+LNgAuY8GfWXGzM34FYjC7qV1R1cE77OjpkyOrE
p4X7PiuMQ3RGg6srbg2a5Rl/ZrB5FDazs8YtWaJAmO92PEwclJrpkKEvTJPt9Fji
nuGcV0A2eaRZwjCeuKmSUf0GYOrzEfoW/kISTKfnSZL5ziZcU8FMkEjGUj6WmSw2
u9gxFBfuxW+28oh8kYhn/OSACHnfRVtcuCYK9/Vv4wS855vYIvtsvGlNBJxu1j1e
iXtCjYaacjRibwKsRkKZ7fEH9nmJmMz1NsmWNFQBlbVq7f3SqzH4t9Ho9+xkfZcw
+KHtH457TXPFr9qAl0sYk2CdNz6ijzvEIcNF6WMCHCNe/9KTNZsS2NqIWp9Uj9wC
nU1iTwPfZfflDmKHyYgYUzbMTtulb3UPbbodznGhOXo+em5FOPnZIfcPCDSQojBt
ZeG2J/ff1jyds3noFSt7drqEUrGa3M/OYhODOLzRRdbzgsTg2aQm9RVTgHOYfXku
G0kgg6ugv2wSDPwES/JhI7T4x1xjzLsJMippflmhdFbEUdglmDigMTLqDmp2MFxd
0LxqmjlGvj8q+zx9wYL5Zhp+nREzLNFIGbpgxu8ocfsVuuIeNZ+ccgSqEPVKVUOx
0J9ZCLvSylH0stB7MVNJYWpURlBzeZQfQ67OKA1oSQfeKPQa9lJILfYGGA5aSYBy
3MfhWjiaOdWWxm3UnBMVX4PFtkaa19ahy9PdO5nx1yaFR8xfSgPM0rKjSJYjyAzx
19+qv7BfeOBpeznTlep9B+OmnZS13AgLNzolQejc2PPaE3upJ5hqvemS83bnEXio
UzqiK0F4wDKbfAuCkQyTzBtLfu+MapGnq+QC/s04PXgwJlv1xHHC5OZGKT5Y3pdg
/KH7tI4TXeKjugKmVw8iCobjmVEjyrUIVUKN/Q1HeUB7CJVcg8SCb12U5OhjN1rc
IbDxhhvGdpvWnI0jsBR8Z+UNnxgLI3iW3Hzswdkp3K14SMq+um8V1McAEqplEuX2
9hkvBw3trQZ+HjiNOl4BkRipQn8W1ZYPX/eL99N0mWTGaTRS5V9Rr2q2YlJi3pit
wxvYyu4cR+Q9k1SD5P4iISHAreBcgQmY81i3Fk4funs3Q3KCOlL2FHfOfB6XOWk5
YnXvmRr1ZpIKOwN7Kf3rJz7G5bdoeFj9XYQ8MKqpSDeiJXksg3EKMpVXLvJqBeBD
3DI98VBbNrBr404v3Jvec0RAiFq4u38QkwuZf9Jvq3t4/Xl9Tti9qaqjm0J4iscG
E6TMqAGnEFz/tqKFw/ei3LaLX5uUVuNTFs5j2YM4xIY6Vt3Rdtu42NKdk3PSuB0A
bG2h80wre7vR+H8xQe+0sAz70ci6za2l6tGQAOF2TcVlLZHOG2rCmmn0YuNfGPVi
6J0kmELIAomEMgmWDaxiwAzX1i4NnqlNenOUDow94q7m01q1GlNiW4IbhPwYIJk9
Z9U/0gQ4s50kPt3HEjXUydPFzrBmeZ8RkqdnHrM2+X1z6EuSwICCZNGFBRV6riQC
nYc8w9luWwxP3SUbvkqT8QbELVy+qHHMu9PoPoQDSxbHVyhzYi2dbKOFoHloCQE7
24Yu1vF5YE0lfC7lpjuMUhmVwcX4Ro5kI9Hn0dSlw2mj6KvwaIwbtDqm/CiXogzG
2eTiVESVl7FmG7ohebhLCo27ymokCAh+yDFsg5spaLNHyvLMKOHO//+BzROZogQf
wx5Fg6udE67tMs1lnb8VD9Kb3UQBi3Ct5J8eVM49jFahA6WVJVG/R9jEpG1Qp/Mj
+tvGE5SUbXawLVh4AtAhzxecv+mZLrbRIg+XLMdjfTEqUzbOFnQujf0ud8/jMOm+
b2VzqV54Dll+azHP0goZkS/oI1VMlcY0Ew4PjeH5vO3fvEzNi7MsO9sFsCKsowDg
MMLQl6T6NYqQJjt8q/8h9mAxcexQn0q+0v72zPSqDMPQ430JDA3dmw/Ewmwt2Y8l
ZWPhRv29ErhOLEWdk/NDaxMlDHaz+sMqImMeQazXmbX6Al2s/hIB/Na1D4pCcQUZ
lr/zthi9UgxQrjSi9PJhZt/eL1EtHGttOOeyHUJeAwCtAratXQESULV9uejNrkdP
TUTLfPauAWhUnrcLXx6G0IgI3dT42cIxl/FOaBerGz9iXcOPheWZApFNxtwJgB9B
YURSC4qtG1eC722CkLdpfDPPwwIebFX9pckbRpRxvxfa4W+AoRWoBICjY6LBVYJp
nP1leJWBXxWE2hko9qsWXdAMaA21Q52mOh9JMi4LUGWIaNQTXUeoLGjwWFlD1EbR
rIYy1NKYoNdHhheCoAsJ8EYHDPlgfmhEvc7dt6BiUwE5WnaV70UCG+oFnv2Bl3Xm
WknAD9FA8pZtSvxiTsCf+xt0zdBSzE6tq/+UWqB5qObUgDcJmOO1PokoDluHXE5+
TmmBZ26g4KGvxxMWV12h6nCEitg5ufpeutF+GKv7/p/NmqDuGHDXAUfyn651W8Xp
562ZmxKTgZrQGk66qCV7g9Kr/gfSF5aGB+4UKXwFwfh/BtTSjuUNSEjFfO3AM3Sw
lnBerO3PZCL1eBBntg074fovWkr5rWKS4kJC0MzXx/MHN6is0tLyWq7rhm4gXlDV
vD4yvmp8/k5Qs8KP7Y4sc7Jw7RZTtfacUKnf/iOo5XG3elD5q33uFQgjqqdU/jyx
jKfyRQmvcJHEuL8U89JIfmI9Mg1zffIhbdUbMCs98BBQRSt6aNYnQHEMnikVU81J
/O8ZBc2YudfV3BCzHribT82Um/9NfznAQ6830Y5N7+/g2FR3vX4AcC+bVpKGXuXz
ytbbIizEJvJZDOE4Ede9vxGQXOiTH5oYIGRNgqXAiWHJ5ltfCaKgjnCej1v0XLaw
bkKuQ7qsOOJVP0j+VUZ3lLg23UJUzLveBiIl9lbYj0sH1PIG7qeh+M5Imvx4LPGu
IFqGcBNVDYawyg1Qw244gUVH2wZMqeTLB5jbOrUDfhY7fVX4Fr+P0I5BIjrMFqbv
XVK0+sXD2LKXA9XN5gn4a2crc+Z/au94ea3UIRcMvbk6pBCeFYYgHwKfd8h5WDsY
qCm/KhP7NZOmmX3PAfjeKYRatdsO7JHvFwamppZdONjZiB5d7dyon5ZQsvqRC7mx
xGrQJcGGtuLHlCh5ZFBJyw8h6MV5v3EswPM1wXpf6HPyTo1ug/PKbFRJwNC1wtP5
DTWitRonc0FOqEcDIrQBPPu1ophVQ3CeRQK/lP3dyFr3VqwlAPcL2a+JlVX4QbFo
OPazPz7WRTLTLe6FeMIbkNwPBw+JspiAFRVaOZc/fmkwLvvHJgNv0ZsCZryUXrwT
TGNBXPOcghCmEVfculthIXzxx/pB1k+0oVOi5arWTqodq3RYjLaAg+ZFj1Ac7FQA
nkGPBeHti4IbOdUhzSmuqNgCU7I+/TC1oFhu8dUvQR2/1jdUK8FnNWkpzY9/yWcK
BgGYYPF/3wembM503L0t/eqQOIV4KD4XVUnrqgAYuT8POUn1Y2xTfNFJMlixjClr
cHN3N/mKegTB1mEJrZRhbAOMlSQw1SmgH7FwXcO9b7xGl/rNx03TsFPdC8Rway6S
9BDIc7DBg+AhhlQkBF1Zjjafp1P5BL2trWGnAQ7gg2BWNj8AlBWV8xRb0JaMX/rj
8u4NCt6/LPH+rhwVIqSL7pmiqCbVhpc/GRyqtEjzOkS6i3TNNGxfA38YRBj6CzzB
9b8sE56tVUDa1Rn+ae6NsXzKVNUOKoyv7GfFMaKysVhaYJg+lp8uNzdm5l3RX7JK
zRn9RRmxLyACtpxdYpXSFCSE8wps6wokUnekrD7U5TNM6BqElnEQG9u45ni8jlhW
aSVerzIN464fHkyH4LBxpKy3OAYNCsclSIyqZTgT66fCP2wC2oWbGxBCWz8oKKCm
oa32wYRI3hsZUA0N/xKHuRZpOWfvdMVuP6Kqvh838U9ofSJeA7wCXF1Onf6zRrVq
p6pIP4VKKRML4k1GuTnRO0fk1GYeTLwp2ff9DnM5rc4ecoXT9iv2DJfZOFSpz2KT
KfucH2fRqibBEnPkWD6G9rhulvbhMfk38Vsdj5/qFjWqBBYruxUOpSbGjq59+7nO
T+R7+NENO98Lrzg+ePMLzkcE/8Hpjx5gFKcbzF4G1OYcxXaV1ECHohk8g8V7zRVJ
B4GHz1LG0MvuFNV3Vhce7qdqKyHGIh1iHm9tmurIafFqffr3t/6DAD3h+H27itka
BycIIkwLvLXreNW3M14d/CnBUBlsoXFrz+TqTPIHpHYFiprPRLhtnKnd+I86n0CQ
LG381qCiurW0I5D2uQf7OmD6mHChpdFk/PBvm/nJVEmnOHCnbf8lTq8ZWzvKBoVO
SwkZCXbmNEK8xpO1RWcsDNVEi5ptdRb1hpmL3Pqq5n11upv5k6Xbkj/3WcfVt7x+
Hm7uy2vOumZrU9ouOfHnptW9Kkmathuyg3x0z0rdDtfm2888VRe/eF35QzD5BpFL
hNSFwYlB08gRTAGgVr/Q6qUB6SMpUQEs4p5x9kCmZVyd1QRuOy1IfO3kUfhbkrHs
/FjZM5OjhuAFg3OtB66ppOJzX2ng5TLrZbz6gFkn2aTmgSM8nkoOUCBuz3l3jSP0
DBxCQgoih5ovhaxZh/r6AHUoJSxUBr3mxfYQEc3cIOZweNcPfgm3+3bdrHz1cQrH
bTkP0i8xN2BJ2dR+dhf5L8iuJIvHo3KuRZUXwXcwmnBz7fO+lPPvoG9UE515BNxc
jN92E+Br279u/tteFs8tMSOxVHp7Lf0JXFwvtGDuaQHNYivxyycS6xZu7fzCDZ8J
mh7aol193NztKGXQCIHbZYc+keyL32t91isrg8CpclxNoN8DE+Knx54bMeeKhy8A
0So5d5BR116/3EIqelFxsTbYkOm9GpjAUSLyDQNPS8pbqTwFQM2Q8deiJ34AUqrW
rnt8kr5O2V/yER1IFRRS/zw3LRyGA+Hzlzfeo02a5IlUuKlzBDuHBZlrDhFyhZL2
OMk4qOBOyNigvM8HUHpqoHlO+RjJsMvWeSAQRgxQ3aCd8k8A0Pemu/knTyf4gEf2
SdPsUcmJqlUTADUEXIcW6xtkVDPu79IVI/Pm4UUNyVYHPUn1WWs+/uOtHINFz3Nr
+J08y+5wIpLHHGgWxii6681Hec+sv65htHDgVcDl+kXfoj4/kxo/dfoowT6+y+wV
qzkvp92IVVK1GFna/9XCeoousCbmG05R+4eCBse9prK/2PEos4k5SJwmdAalvkWz
1K2pwdLfaGTrs2iFG4U2N0oUZJc3KjDqWi2mAe2Y6V6t26NBE1jMIf6d3wd7ETOm
KrSKo02IDEyxVhnoXF/jlpwNeM7qNh/YOhRyVGN3BfCf6A5N3HrUoBfvQsB2C867
NWAfk0bDnnDAcE8eVY6kmwYvvehA60Df6fdDDKbhoa1PWx+Czagv8T3WsETwwrDj
pVMIXcaTfAyBj3vklOcd0mdbC/iPFzE1L5lyOXWii4dEmTSZnnPb/3M9Ax00AGcR
wX4FD8+JMf5IhPflTznFBqs2YuHTe3vzFOtgnSQYU0WuU/tYkYvZr6W2npkBvS6f
m6n1GHQPllzv1CXIsM6m1NezSDmOSGJnyQjtSsgggcgETiltS0Y/Zaw6DekmRgZe
qPxgo63ejyU2imrCXjn1bwdmNf3bd/yS9cMbjHZlRy0T+gd4klvh32VMxuBA8Zw+
GVzufXAvEiQsun+HGXRY1ndL+ziuu9tRKIqpBOii1tWDcRru2Qfu14Dd7cfGHGVL
ECL29JDvR6OqrChlqROwqmJzQhOu6j5qkaR/EkYs1qRq61tGpkTHD0oOzKKypXD2
4VmAeefYye9lv31/gQx8pjE4rnD/bwxV6sVS2d4AtEJ1Dxg9TuPqdMGcHtfObtdL
g3K8gXueRnUAyOF5O+w9N6Dcooh5/G88hPX1gVMFIqZ286XNjIgPW2N+VCSShRgH
EqIxaz5L3vgTdi6/e6QUynap5vWKMMqM9eEjSXCGfNGwPq5b3Up84VJwaPQ4Y8mg
Ut8GNOTBM9VRTI91iPAJbCVH25BkobpWNL0Yky4IxrknPlDkuQTsmVH/RBsXO1XY
HY+PJewF2i0h+wgQ8ucQzFyIToS7GeFai/19eOM3zF/tt+TWe425nBeeXAv6ruDV
qfGZITYcw90/BUMEjsCbC6EAxg4NZP6uFbzQB68kBCkyL6LWmQwo7AJ67Or0u00l
nZwsvSWZPhvdLUvyOnRieASP2roxtQ0h4gxIW/Nx0LDAgPTOm+XNt3bzF+dT/Ohp
XtKb2l97wnkhyRiS8iMT2LJ48VkpxD1ArWGMjEsTENVN4YPF/jk447YtQPRzIZPj
upNCWtqu8ubMfxvLPojVroYT7nJfKJmGl3B0fmewZmJ2RY7vSq3jFO/JFtSk2IZL
tvHJImNGthbifB+WgcBiE3dmjApm2f3SBAia4FMjVvdaNhlumPRgecGdrsAZ6G55
cxQuCqBwF5tWLRJ88VEHy+nbB+XcHM1YTRZLuHvFO6we0OOVYhlV3udux/ZabMrl
`protect end_protected