`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
5UzYaoC3tfpGCmdkAmjlgsmaFvl45qUiO7pZH8R6GSiiVi7yq/KhNfySpb73DJcm
2IlNVg1EiaTij4cmwYlMi78l8HGIqeesgOW9xbcFFxIpFNzO3jT4WOAKcbQ8jGWQ
KAbz0B9NF0sZp8L+DVHqgZmrRn42aXP5q6qBkUBn0Ngyy4Nd0QjSbdkAb0m0w/JD
sQTUzxg/l1IPiquS6ihfwATiGieEL8DnWBFqrRof5c+fV8+xmcZ6+3/EcVYKcD/X
sT0RUTrA/em3DfOhf1b1Tz21BhhZjP+tCEvkj+Q/lJOF/Bq0cFh6RrMy2nofD+5z
KSVUnuSCU46whFv9fEk1uJcAZXLsDFPoakHO4wFhoThUbYguEYVMRACGcyz/oosF
I/eQJinTaOk2bI+/eYT+bvyy/zvIlkpkbg2oNcfeXXcyFrz4HOx1Jwokvv1hrsPV
FeeJbYgHJMI3SomuWZ2+DRl1pZ+YDW3N5yLTMd5xRuevG6jpFwU3zFFY3dkLq/xZ
go+OqHnlv57t9+ykcWh5Q1CHKo9KsFq1OvNdVbThVqUQVk8HG6KErXOCtI/cE0mo
eC1mA78Xi8mr9lpHpPtQyaFkksQBpEXANhuyp+9uNi8SqTUf12tIr+H12oKMKUJA
ssokfdHlEXGalKrcH72drxL2f+Tt6NIlaBwf+rzJ7sMLqef+/zcmnIIzgd4auEl9
WALW+G8ouCYcQb6owvWg6W5jBuPCGZgwmQWd1pQNswBCAz7z5mbbnpDjifSTMKXm
w3gkda4DA0kKiXgWtv5Q3Za/P0YVpxp/4972rpbX3V/e3AI55eZKPMY+TwtOxehK
gwibQ4AemkAHmtxLA9FMOW6z39n+wQW5rL0UTo35xU7Fy517CpIL5DlblbFCBLJv
nj6xU1mxaUanqJ3eqFKv/3ie4NBxZcjPGSRjkK/0ZuG6flWzAjNNEpzlFBMf3vGg
Anz0JxuzIVMYb+h/Osq1JR4ovJhKw7zFx4ZHufiNbPrGnlpiA92wCAzFPxRyt4cN
GHrGgqCiJKM+oyI/AkvpvdnZ8Emz0oTJspfSLVghcFFNiGDmLUK+/b+eEiT80jvV
sHzPfqD5NL/Cl3L86O/OWOzbPYxFCXzIfgVoVcfre+d2K5SXaWE3YTig/gqPV19O
I4mRJtXEmOJBa40f/BVE9eyBJ1+9FO2V8Gy6AOYw+vU4yb+BiSrstNOeubw+Y4Vu
p7Z7GLOR6VsX72Fxpgjo6Jlmtf8Ei+xDnyDyjw3uD76jnubFydBhtL/GjC8p0YiW
XhUCO7tKL6l3cMpqvPTbuBw+f1UPmnh/fuH3BI35VGOiJjWgst0CqySfJNMFMA/U
0ZWWwaaSJdzQHBiqg+BXeD+WOdX3FdbI1+EvMF5DjZqkYQo9ItKxFxozFSxPJuV0
XH4R5FjTQ721wkd0CKXzmj280yE69CNE2X1nSH3nJItp4rGB+x8vXU4zqamx7NN2
GLVifG3lMuQqbrKyZK2GTos1WxwtWy/DLt2EFUnqBN3lPlRo+dhN5aG6Q92CjA/s
pgE5ZZabYe5ezfuvqXlVSv7maFw9TgMdaN60hsiAvLN4GeW36f992d+lRIb+nHLQ
yv2bptZV0GgimruPJhN2m0bkCzbXE/0+42IU8soM/SUjJXFTMRXgHTaMbBI/CMFP
0bXh6D/II+uIs8mvJ6yOifrRy3mUEPD7zjAvrmq5BuE4slhwc481YqRFSU/5b9M8
//KTtHu20JQO5oTz/EUJZV60WHRqczy9n3ZkBZOrZ5NrYPDY+yQm0bBDZnNCRWF0
r59A59IhLKKDB5w//I99vK69/OCgLx4x91ES2QV/CwY6F0oXkg9q4Etv+Z0Tshhb
Fpu9q1hYST4Y617EioxgLIDE+nJuPrL1IHe2K+52QTyJ2dx1F73BhFDI8GESZE4F
ram+NkPEl/EMp9Aq73KYPc+m2evvqPrdHcHjmoi1/mj9wNgn1vHdTGarN0jU6J+1
h10ucRFXJKP7QGEUK2Es3RvSvx7uIXuQKvRGC1Krt3p1aCRnHzZaLTri88SAndMS
WsdJT6D5sw2VBhPEO0ZNKXrVJEgJXwhdejTcXYLSaAX2z+gr3beb9UVlSsxs4Jmg
U6r1RSRYdnsaUzmQQEgR9m4ZyXt86OLtIf0COoNrF163uIC5nRqjMyQYQyAT0+IS
hOFY6NJpTtRmQvp8DilgaoFJ8K7ocMSpVn3EulBa20l+FqcARLnaAgtphhvDsce6
UzCVAw5JfTwVIIobrV+aqbrVhc3IEiHSnNEFXbqJKEfdO6bpfF1ztIw8iMPEuvpj
OprpMbcKX1zuPd45RhecXgwunUD1qU4klA/dKSkEuSCoOiCiIkfif/jSNn+XD247
9GBZaKKfrlm5EYiMxWVeAtKfFrlsxR+O6US9mZp1IUXjQU+wfw4xHrws0fvliQco
Y2b5AIy1JdBFg8N2ggYJY5it+a8uvyFZuhRwyrIVq4g1lhIn2AMuANQye7TmtdnF
LWqtsDnCrSLHqM/RnClnDPQzldw7xcG64EpJ82Hvj/XoQhpKQul58eC2RDEHx8hg
wSXUE9KLxKMH3Os1tA1PbjC7ZG5cF6/DN2PmJiWq+BpZP0FxtfZFwqNce6joKXOy
+P10aWqTBy8v3+2myHpXmeEwzJ4MkW6G8y1PXlEnzbBbOSzsUXk5mP7H2iLRda58
WnPlczFE1AEeMkDxBoLOBkIHv2H0lFH9oAZH+3fQHunsIvvfFGt34WyfsJR/Sy5m
9BAFbPitGh+8Q/XA/1j9x8b+4OSREsw9dt+s9Fxnxjs2fqF0Y895gbEo4pV49trE
MuZlP30OuZNVG824uzwwyqqR/XQUPjA+a70JBzY64Uy60kCkQRqOP8hMrE9XBDQP
EJhISSN1023rH0PAVAzfXUZuf7SpHoTcWe+QxIju1oG95dXtdO1qi0B987EiV6Tw
oukL9Wk4tq/DdG8UU32xPIvAmX2Veq2imQbjPbhZcoXcLuEefvJirPKYPNtJBL0E
QqUnKn9mScn+zDlSxXz688hUCB2QmqgY4phAFx3CIrRist5fElogBuwsq9aiSVZP
YwVwac0IH8j47JHO8bt5GWMZR6L8QDoBRhLf9vZ+cNPcNdZiYOpBXn90qeUs7pGM
cdy81f6MKcq3fPGND/xEUDLotyRRsa32OjUA9PV16vRkQv7hiYxyM6suznWI2Nsg
uNhgv4/W56fYW+08xZvONPHBQTmwUv6WxS0XkWy6gHjiVmUdPYG5m3M/HCpELxlD
nc1HFbLfDcWkzYjLlbwdDarqn7d7KCxLWMMVVm0Z9IUOFsDChctRLUtFZVgTr9JH
xK3YAgpX/ccZEwDG00EPD0C12VHQ0WzthlbuQ/H9yuYZfRlgSNCZY/fQZloCptSN
fw8DMDIM+gH/H8p8hUIf/Zs8X0BsW11JbA6w57TVgP30gDskC/aMrWGTxlLZydFb
cdhXBhjk5QoGQPD+sZtQHZN94r7NarqcFB8xTGaBU4BNRLhdHD98FhJ/bJZUolmC
p3hqxJ3AQcdC46NeVv8eTZiF7WCrxL7zvaRn6hmMCcC6AK3IjaQT1+WM8IWFHhwC
2E76JHGq/qZikMmEuPEMlCroqL9gw+HuKtmzLdp9G16tv8IVLYGGGnqxZppQVCrd
0Un5CjCTkfIGfC4l9vw3zbqyVNomKXU+eEAKFbl8te9pz6I2os+cPg/7kuHVF1qf
Bo6x1639+x+uAoIAR1Sfgeeu4V+UohgKsY9NaLv03IUQPNrTPtUQioSqZrBYBCPp
5AmPi/NE+lnfAVHzVciPsUUe0ikVaTeaykM7+gHDMlnjAxTJ71mb2W4xdaUzLqju
pVQmKjlj5niCB7eR3e6zB+/y9kVOgwQusjHaQs4lBJGr4agfKcuB25iSVLfcTbvh
JSQoxzDoeKlTs/lPagtcCsnfTlvpQNALX0Xz+czz+QAAjS+wzZZ3cTZXy2cIQUKL
2zn5XF6zJFigdqUbYEi5gKzxJNtk4wgZVklcM9xNbimGh8/7PFo6Ijt9sK4jLvtC
RSeLxyK3LYh7bA8hPZQNPm82n/3ncYJnnvrigHEIco8+t6JJMmTu/ydZtt22wHRN
gs50MhIvXEmxa/2pMIzM58C3+A36Cx6ZUY4AEAkAP6PMAUlto5MMvn+kKBnDsWae
9+FkkkTHt5cef5tCApCaUK2zhiQBEHagUKCfOJgYWPkR0HfC0yVYalRPztqNFSus
MmGurvZXojMFjtqv3DlmZja2foBZMCKTdzECop6w1yLZk6c2+F7Ejh5J+/BYbaIK
ix0+m7H+i1HrCqSPlK+q7nJzKwzfZyrb/BAzlEbgEerVCHbDbhCMHVR7Xzn/Iehz
lFf8Zegqx3AFCcnbLzdiNQ4IbEDcxNNv1mCwfRyqR/JYqUqGjRTUWa5wz6/0cX74
p2pFEDYafGTW1Amrpn43E4LedFc4W2hwHKsU3qMMPi94CStGn9wPO5NXILokK9vY
89eXKuy4SJNqYGgpURGhQ86xSs6MYVc7++sm1JuQxmPswVSK44tgvFaSxr7Zj3Bq
LUGAZk9MIdFX7FsEX1knLQOwfRX+vwVQjirdw+QACnkYezzptcJ6AUQDzxQBk2O9
VEtKiMz89O0tgQoGVO0quVXbFj6cUcjEqoiqB25AokIX1OehssJdz0H8tny0D+Jn
gsifpvyP3V7MeQ3HKJMCJaRODLIPbWUPr2NYKSfHNQ/MNPggClIFpIvVp7VnHJR7
Ljq5794KL4Gr65I7K+GgqDRaq2IDsmqs0ehN7x5gD1yQmyLv92dMQu1dPiO+C5iX
WyBBLDQS1sWb6L5QfXILxR/7AaTHmVNdj5KaAOJFK0J4HIPOUjlAPzX4AFWSJLpb
4pneJbJ95Zo1xv3goQD67+EKR9OCI0ZattYvGGWB87lJMqO7HAh+acDY2GUKngmL
5KH4vJbWvDm0OhBZmdVItS3lhashGBpy+z+phh5MUEIZSes2DgCqkmTMFOzGALRq
iFqrcau5lj/gPIjF8GQaxmxkIAaLioD2ZGb1hwVg7Z6WkZqmOsc0nlJkngpxqo8b
Z8Aq9B/xtIZRk+4YYrV/sVTXJvqLvu8o6KbcrA54BTy2amJ2X1+JcnE/aNo2VW5u
rzrvS+6fWhzDCNCm39m2hRUey/zgWDvT/yxBYCsRMYoXJupUVqUDhRAhhri76334
nSZMlg7dJutnI5Sm/lB3vuh7aWEYDSGs+jseWZy0+5aQzwrqQJ6As0SUMRIT8ILM
qhIYTMUcpq+KQ+OzSgcjjO+tHFIHwdvjJU2AnuwxtWRjF+cJcZDOcBxlcIQM+a+I
MraHKrUBfUvlWAzl4Mijvc2W32iV39pIua2RuTA1lACS47fNUUM7JXgEguKr7Nwc
ERIq8wDvubRs2Xqk+S4CDh/cjjJLW4Sf0N/W/A8s76yWWc9GGhcqijSlKmNdIh4h
59HEizOGAttZYmqpkwMuBeCXMyt9FXrsOAeEkRwEVhbGeGbyYB7l9Ge7sgH0tT+C
LBey+levn/KR/d6MNp+Aig3ylvMtmWKgKT+u3nOXlr7raEFcUcgD3gCRKdOonLib
/xY0NYB/ZrySLND5Eeit+fwiHMI+Hz9GdWXq7j7++9XsAjdQtxqns9XnM56k2cnf
cMyJCxSIET1L26LaHOJOQ+n383esPB5AFZM72sXfV/j0bTbg7KZEwQ9eO0tEPvZC
zoTEn2trGoJMW/mltUcuUTCY2+ZJue4Pxal61g5rUfddfNobkZiIGZ+AxFAYp0Iw
OnASmOm42Wyoe7XEyhMyPt57lUpBPCbeBvd5GoD5xyj8l/AXXkwTo5owIva3dMLN
pgb37l+RTj57BSw8q5Nghm+b08A3Mhpkt4sBbxtw1SE1Y/jIcrWpbHcUKv8Pg+eG
J/T5Zoip4E5s7vzvK6QgwPhRPcccom0CxCrpIJNXhcCTSfq8tTO6I+Pa0IwwOpbr
ABHpvjCHAs1n8EuJ77X6KVVNAG/u7RfkWRfG5wiNNoBeQvsEdvRwcOkVBdCOKkNr
0w6nru8foSwSQwZgg0juQ7QIM9fm6aWpSTF1xo21DnF1X8waXavVr1+jRGCd4atV
8HkK1rOoQTSTz5wAK8NQ4HY6Q2qFzxPtYlBBz7fDy6VqYuBsjFPE7MOEpmHwX0t5
MyRbhZxrFeyiCr8gMTad7LufeY+3o1LhknbG6DmQ55tese8EQdPqtFPYRoQMJzs2
wfA/aTIhLjfe3/+2lU39jgL7SkkvdnjYQ2kR/yCSSCsKVlJPCXYu86M8Utqxxp7t
fI+NA7IXOEAbDiLab23Ozo7zLjT8l+DvFdkcYMGn7XFpc1JGfopKwB5KxJXNWi5n
pnTzP3PU7XyOBHjHvKbwlK8mtf3xa7bGlX/btYACJy0c1VLEHpidxQI17zH+Z7pu
UN0m8JVVMHYHwojyeMGgHpmEvDF/tO6W1RFeVROhYGxwTkPtVzu1xQGMmjUeFDRI
5yYi5g/OoAM075bbQfZfg5hZ9DV5/7KRGI1pJqAuOV8zr/O5rywQ1rVg/k3dysxU
sHgKVADLRWVA54M4go1uzbWXZRyBDAsmbMPdilSrXHmacxVwP52DAcN7GXij/vE1
w/hOyuayUZkpIkitwJZTwbIhW0QdRFui7RQOCJd2k4+L0WpRnwDc+dTjm8cyx6aQ
OnezrtZznVXmeY1U3o+0wKSJA8+2zln9fAWkmPXUDwYs2INZJuopS60ryNyQWel6
iQKXwe8sfVhk6hB8+yN4RxXVjfSIlC24uvEEkHXqq0CStlKjQ0DV84eXnYB/vs4L
WchrhggjOmFzrGIewVrik0NLQdwq06cYSzz7SVsbZpnAKEKHV/h8xN7vaJNLBrzy
Ch54oK0A5oeMCqVxGyeKPC1SB+H18GPqXhyBYXGsOSfT3QHEaTLytxMIZfI1Zs9h
S9iK9yzv4JODhgfJdRYAu6kbwQBQ8qSWdeb0BGzdrTYYt08bvhnIKV+vUzQOEdDc
t2OcP4kKMpv4+xgPgoUUDui5ER7tp4PaY9d+l+aojulujV9dnmNeNiOZKiDwhjKO
jbSi38/r+wvXWsPSo3s3YO4S3cNIsLpkw8SYhZ7JcTPUQcRkFhAA0ptvgapj+7rd
eQhrgklmM9r8/VQuRnldHbZ1G/FHALZwAv+cseWL7/8X+Pkhdu2QRlk3ReESVj1/
uIg5HYJXD/J2np/cVtuXm908WXiwIaVk5bZ/Z0HfP0KfPIZYtLvQjlI9k6r4q+Ou
nIOoiaPGADl+8lfryC7lEHM/PmXWJBBZnLRukk5slNX8eeJC2F2Ie1jn9CSkgkaw
rzq5YnNugNcWMhLSqirQokWAQBIFnCFddi2NFp4D1ep+2LtRuKeiS7iH7yoHMEWu
R2XUbwhoEcnuT9ReoccROVn/1kq0kgQ+dl/BuEx6rBJV+MaLjqhoxBbUfTsct4cM
yDxT/Y32ohqGwz9eq7tTazqvnKEBA2mVPup8j/ztDita2ApEiv7QFkXiD7V8yzhr
gGCoAg30/nxanWqccjyvQGX5Hnei+4loe1Cnxa4CHZjgNrdItskiwTJ5a96AddcM
J+WcqOWuyVSxQBW3fkbGqdQSj9RXvTYPHv8A71H3pKp1keuCnmqGSkeB4vz3AmYT
oMvde3aU9QK8W2iQZfAOQII02cTlkcQSh+tkTHweDTZBy4I7mJAGmZWtWBh4QG50
017Yr4wsBbHo4weStv2pNw38vPKo9CyOj3LGH1L/k1DOO9e9HPiUfCfHkwli+GVq
qUDf6T+gMAE/FacLX/fSf5kCPnHX1l0FcWFB2giJKs1FMcJ/mOyUnih8kK/smBRC
hwinnr5v2WPnlPSgYon3cdD4RTt7uArFumZEyC4TQgXC8aBBUPRnTE5cb5mrVXDk
zqiUs5yeZQLCndoFS5m8dxNJvFUqBlonhoMAJfOsP4djo5ddU/EVoKrFRkdHMA1B
KW1o4KLHDjg08Rq5A0LE1b5KosjnnB8uU3stsx0k1Pw4zGWO160/cEHa2YL4Ih1A
ygK90eU4+//5lMWGKmfsXfwZGp9UNpLZKW35/g0y2XzG1VZSMklrZ3w05y3/6uGO
EXEbo8AJN7TEYNpXP8gMo6OIcCaTdU7R5wjoFMMiI9sCELJTp+UOEFMGJnjpnC9N
84TIoO9JmC0pOQyBVt1j9rkSkIA+m/GNZsjK+/newc6uUnUTnScBb/CXqyEDXG7g
oVSVA5Cjgpa5yoKo2VNOYkwnDhf5OOyczbrcIgTMAb6i89Vq3DToy2OmKcTYDsEi
jo2ADuw+BQk2Rr7EGTPOeBow23cp5Ayz9J0B8uUyUxoejZS31OwBJJ7qukVShXwf
dBO+wTIj3G42dRh6wGbJwIx8P2F5MM51zJtfQ10rOgVHUAi6LPAX7L81muTzsE34
msyPOsBd5ZcLW4vgzePsxWoGGIm4eVCV2YSbN/GyvNOLRq4LDRBwSQ08TAe/76wz
klPI2Fh0Sru+gnP/cY8mtxtGm8gdJprHI+5rXksMeHcUGfTTYo6Mlj/Fjie4HYXn
Itih4hnqWUkvFFOwmzZ+h2i57LjZLe/XcLx+VSRIeZoZKvyKks+P8lbOuqiaRCEp
/jiZ+Uvht/Od2rTf7zqHcoz9JgM7eaImLZrciF2Db47o0vkdz7A7ON8rnWJaTBmu
N5TgEffEwyQg/h94x1RojyUQNg5n13MqB3S/WNG/7k22xcsPIfaHA/lgWlBCFALV
0ZNddGSPlAhhnnYQEh7/d6C8LjKFBx5yNQ44QTaCKE46NlCoPJVV6SAklJzNudBa
V1xpyLgY7Ybzk/6C0OlD8aO6W9gqBW45/RmT0QEKUWeGKZnNFl3p9LN8sd/z7LBF
l9ff0Cd3bAAXLFnhQ5oYPXqsHyPpDCCzzUUnb+O2aLyJl8ADIKQpH0oKET3G1POF
VfTcFriHbjr+2RUtkTAZDfBKyv/PxZT9KIwvxHgoKYiNg6FD0v27pT6B9KdmTSNl
c+any5dVdRNjHiHYZ71VwR0uL7mhqwsFyELCsD1traZXXg5pfms3szuRJaEiGLmH
W2igeT2FVfXX8HRoKOkekC2cNA/YfHxnuHW5dXMpHs96n8Jo34SUJErZrboqHfpC
tIPuVtg52PjwwPhYOAGv85Ur3+YS5Wg+uUKuhJ1SQWJSFPs1am/ukGYzbGFigMXq
XN1cJTs4j5IAhy09rBJ/li4ywfrX6ym6F6wnekqUYJKK7SI7x/lQOSmFwrj3fLl4
xTVtDmDzwfaGyAKyj/z10RkZ6DmwTVYoiCiocBsCMmTiIvSmuljgGu+ihs3Yxvpq
Zh4c9sOpnDE335P++kzt7Vr1hLlEolFJ2JXMfurHAGDsqFz5UR31CAlF39PvW0ym
sflOF2MTP8A4Coj0+bVqfX+w+Niq1dxNedVO+Pal+E+NthMjDaDZHH24hh0EewRb
iiRJ+3e15KDfp1wXBIEruMRWRDEy4oli5+M6zEBjkZ9M2nmZPdzHGq2NWAeaqva4
bTGv0dJi3T+mM+rh3KRHsDMEziMsWHY0bSjswWbGuSOkQdWnWxRgSqpV7ZNg05gQ
QmC3B2RX6IpfeE7nfbp9bmEMcu7NRlFRpdAQRpo1DbroOTNCyroDHoRkBXqnobMz
eis8CgGB1qCMKm9KOSG28val2T8S3UEGKbA2Vqc8dAbSOVj9/v0EE3bPGbCoSLU5
bawFf4JGDcTZV7wjATWQ5Q6Mqp9Pv9IpjAFlOdcBDxE+nuwQGnUrKzkxeUizDzCV
xqYPi9oq5FjgH0g6mScb0a8LSUW6JMRGIX12Zo0LBN+Qz3rzhFflwUrYpgqGfSLQ
7+5BZMFTG06wivfC4Xtp+w6wWWQUPbjhiXygznBd1gvtrzNWIDDfL+/4bq6OASxi
guUsiKSsrhQF5ZuK4rzSNg+PkWC2VK2er3CK6XK0zKAW8ZsQdm3Sx4ZaG5YJUE8F
IhrBKu2lcr+Ka3O5A4oqu5LJiS34chD1FS3aE+kraFex6ifG9xVUPWkUpn7SkEFK
rCdEG3sQKGbHHX23oOy3jr4muBv2CRCaZqP9TyhLwZijELkQo/5b54Wyjf6JS6z/
VrhfaZHbui3ujzzjhVQAOeTEly7qhR6tbO9+QdFGxdRlNtwVdHWkHVgAIna8LCCT
mgm0j8FbL0ETJQOwtADxjGusdRE3HaJGf3vpjm+G03+OiVFkdtRB++loLOcSl7/T
Jn0p45aiBQzw1ON2/KzFFyex884KCdiNNJh/DSXvT1MKJhoSEmznrOAtFzQytWg7
Y8biLUn7D3rL9dNYs8LX81nC2U0OsLLtISSfEwbtRfkNByHp1GyoXVBxc+TvtNZ7
LPUp2ZNUpyL6SlhQicrSS/e/qH02AkOzes0ViZn/y6qEfQcyy9e9Bm6nJORpNk91
WlpfYzGeOJxYMtl+nleD5epiENohLVnrzVyWmCNw66gmNOk4CMHZUamDoKq6gtsk
Eql0nq9CB8UkStXs1SwRd2QdRnC7lYbdCylnRlJ8n2AUcALnIoWj7Z+4u6flVhb8
482afIOA1AWi997OZF74sq8evIKGw2EkVYITFmEHHJ8T9yGSiZnzVEsOdiq5EBXK
2w0w2vNFEZofmTSf5qUKLfLTadGNMFlmJmk8IfOfwMa6862VclmCBFMZdRGGV2es
VRNdflEIzI+svluDKjEDMOTUG0XZbVA/tHTG6BUJ2z5rlova0jwKqzff+Fy/4Pu0
V7uMwDxF5mwje4ntontUD+KtypYp9JXR+LaErajj5t+gIu1kxfeBWUCichczuI46
OjoM5yLaNnqiQgmvKIzeUs4Jt5wnTlctwRmS5nY/dGdPp0oaLSKFulXrjVfs52pV
kWIDv/lhSAu6LIy+cSSxqEqkDy+kHMhTvQXb1PdFMWLiozLJrRZCxwt4y+n6+pEu
NkuxJdOmusRujMSyEK7hhSVXVE3YmvpeYJpcqvNzPsUoKO0E+ZNuAxZWjEgBxqkm
CSkKNmAMmaG+4DQUoRr7HKIyrkrcOGee73QQq3ZrA2NH6/WJTwzN2I0UnHtMHL2B
SJPN+67Z3E4v+nE7LQco52E7lfc7Fl7fPCnBxTSOcSznU5B5ukpEMHIcmdAVcHdA
0POB+uPu4U774PyUjJHHoIzYl80ryZ160hPW2YyU+3imh6YioLqW72y99cwUv/ic
w9LRky+qRxIr3f9I7KTczU1i9mpmnCPxt8UOExYip5GuOVsmv9Dn1VOoguDnChnR
tYZTUBniIQn82YSfRUccLxU/rTBw9ufqrWh5u0lwsolNcbNgo7aJNLamKyfdWg1X
7Q1sbDIodFuPMvaAoSC8Z8mBmz3VcH+cK93ui0TvUR8WUreg/3sE7Sobx1qhAjdO
abw/S+TX/v25eq/bQTkO2wRt1z+1vq9jgv875zTkp/E4cVScaVAkXz67H9dw2tVj
bCP8JFKLPZXpg5TjSYilTpiq8yI0f9k2izvAkRcvNUwG0H9D/xLHkfwXnLc6dku1
RB+VC0dlyBW9zeWwEGfcQ6LJqIzpcWNuzlbYZbn3TE/dfQl1rD0ldfDoPfXj/VCE
p4JkoP/PJs5KqDck7Hz6DMY3Q3ZNu1q5cWOmC+48wmWSvgBfrbdOU1KarUmyGH7m
MUQDfapeEIw4/wEdl0GbHGkr5oCbmpLcmeR6k0dfnpoEwC59q3Fb9qcIAunpzjlv
KFKBI0pdm3Q/jpIwgYGuw4w0wLVZjw93jEOiXONwhEJnVKq39S+kBGRcj+DfaRxm
99eifXE9EN9oSJE/F0mhikJfxJ8hffoKiGZSSehp/pJ2l37urvZv/ATd5x8dpCS3
86d31L2/Ekxm+x1LuarEZzqDW9d+ZzTFozjtwbT/CL0AokRmwJdXSFreevQVo67Y
2yO5BBqQKL19pqGd4Or0RVtB0S+kUoiRbqiJrNKs3nRi/HH7nh8tSY0DL55Zx0zj
tAsnb4TGlt3Zgwfg2wQhbnw2iqJYeuVEEKHRdK6Nb855BGI0W+Ff8Bb+Y3MltFJq
dNPPSzw/sIeUT0LdfCgXIItAURfG9aJKkFrmKsm90k2YT7urPxSjKkRvc6DS6waZ
8eFiC7+d+18yz6ESxty46E3UWl6Ge8L7bcdYe7GFIa9Xi8C8VETPF2fZqiUg4CTO
PMHIuV4PUfl81kWlnq8L4UnFEkHqbIPdeL+wz/Cx9eDsWw0RPTK3xSozRRolIJn6
7Gy8m/XOCtELbN5JYXP9WTIhQ08b6uBBJzSiBT03TiTsMM9QY+MVH0Ugswe4WnQZ
MXXarv4yTTKVJGWJ5EL+GDhVrj5BtcmSjuVC7K95vq1cxQfW6sK0PqY9OLYyiK+4
5j+b3r7QxGISbKThrzl3IEHJl8WDbQqfluaEW8N9Muo+knTIfYSvkltZ1HOd8hQG
6VTBYWBp65eGw5Wi4TSUH4DjUVj1qOLGN/Q3j8C9IdFsrJtLIkopbnPgsAgmZnw9
pCdwZQsQnTmSSq2FLAmmAeE5dIHEwJwMTueatr/NRV1khTjMmyHyQgWcz4IpAJIb
ZHic+8l5oNLEh9tSpvXKMU4XTe1VhmJtcm/IqP0t9K/LWnzYN+udDrlce9OFFZ+A
OhMg31Mk3HmcAZooeVzZLiAE5wccZMWQNuHuxe0lZCjLrI0oETtcaCW+6PT0TdKO
Rzt469eA8hquZ0l+bR3P/CoQkfP51CQ+KGYVgdttWqrBBzP48MXFK1y01Wyuh5Cx
hU4VHnLN2WnXYKlau4IwZ9FdgcEqR7Fou+0s24+1PFl6jYpSRJeH6wL4N/8ep9Tc
csoPNoszhTyI/mtN2DVnTxJtdKU7IpWxSJTBGdmlA/zPBpfQWWgW0G87RAc5J/Zy
geOzc0JuM2wNAfrz7HdPgOwB54Z0SOgWyITtFl10CCy1fwiotvkq7Hh4jDF1EzGO
vm+FCjLqHwZWk0Gixon0/Ze9WTGt7I1RcOfpzmLN76P5PStgiUAcPmOnvWQGHQkd
Qyaa4AzYrTNnE/iBO6EZmlT+eUBqPM+t7JHsw2rad1O0Zw+CFLIVEj0bDCUht3Bb
n2Mq4AOcoJFebIsymyDJULGcNdtE4FjhKjyMuy1lNSjCSYsxY0vau3uqOxc424pk
yXYUa8oBnTzYAJMT0HLK8iHyGrE9zIkj7zdq++3mquhO3WKmUFBSUfBZXBYZDLNn
6B+LQqS8SfCD9B1IKitjvhUF6K8hZoshFOvXQet3umTwVwfypSwVBV/zZ1Sm6UPP
thLmcZf6aV1AoGLjfnoi0oTo+Je8OufIC1e6d5Y9/wLZqk9q6KoHR4KNS0LUdpKV
383gQGCPDhHW4Gz6b6kM7kdNIPAhY6NGbEcx6X94lpuQHTo6f60fjc3wgzb4LLj1
Jw2LtAvgC7J/rhQJ2l/kWv4hW1BozgFKQSHyY+Bww8QOXWm0gL5ozHTWilidEBH6
eZGfF8zmoGG8woHXmqbhNqUHviCdScLUx0OVwD9F4yIxS96JU10X3Cjw3TD9g5aG
yK4XLLZ7mMkDSqM1P08CJDuLUUMUHz1rHZePUq2VqzrNAnUhBQz5LovsZgZZYctH
Qo27Bu+MKYXd7tOe4XXrtPS3snr9OSp19vRBo+k5KGhKt2Gxyk/hxTDNY8ZpF1+1
oMwcwulaIzJ6mDCVV0KJHeHS7F01fQdnsn9DKKckx3CNn7/7xKLih3EqmVGaErS1
F720UUB8Zg9or6/FmJcvNtmIAI+axnYChwBuRM2uagsucPJLQwnsy/sHCmH/xtB2
8tVr7Pe/MCZa58CXim9yQsILYO3Nfqrf9sHb66/jKIrVRYMj97dAn48LMxZZ/vdC
HhRE8BmwMLoqlYEPhtH8ey06DgfzGrBquu2pCL4ILHKz5RIVvVipZ2KmxlUT5yy4
DyNtlWvrMmLTeVTwN33itglwYn9oZuPDjW2A+5BXiH4zKsIqkVppkfWfNea45h8l
STsUrsf+EgLz7XthHL8NYdYIinPYcoQdnTJVMgA9PlJovm3lnslyp0GHH2YG+uwr
FZPDVNwRjJxnr7RY9INKG+oHPMz+kc/42jIJAt+/nRPieQIPZuQftTj0NLd8EJIJ
lm+H+fH+TXj0JT+k59KSI7+qtpbnRUW+YuK5Wl4pAXi097Ufh1WER0IixRwu+w4k
dnJlDv4wbKPu+EhCj73oThhOREyCOw8ynsVQJFe4by5zaE5PxYbhPZM1kjKw4om2
+5MVtOyk/yE7mwUVDRbJ4NPn1yZHSFxs53BNbXbCEVk8qWzjNA7csJ/QJK+l1UFq
2ZFUpczAQUrPtFPGGTB4FmwdutmGpS4IBKOVVy1pZnQj6zMM1psZbjKOLZOwYkLT
C6g4IfzLiyz1dUnNwkh9C3yvxwLrWtelt+xkuLB3XwuMvMpBkpf0g8M47PKZ4V2M
tPL/7rl8Yy67mQsr4PeTGDB2Aetncp1RI4Gy0fIiQZJDGzzba7bwama6zxCrYuSP
l+XH+WtBz6iOO5sE3hnuFY/7ePaP8q8ugJ0dEIcY77GyGuL4rmHXV+D+RUWlR6lV
AIrG7tguvI1+4bRbL4wLXqOapVkkhWokm4KcnjUUuW/8cbuu3NadU6oUyXj5srcM
k3TpWqDqBFGEES+V5Zv9XimwT8VWRNePDDlNyfdxtARzjjrcY3R48nDz9skGOLCX
9tFlB+E2/hplvpOsKlXRhmkO3jFORfTH47dDDLB/kDNPO0cujGSA1GgrplZ21P2Y
nvpCw7i6v8D6+vCvY3VBTMkoz2UTNulBibgTNNhv0pKF5f2qj7XDugJvi9SRlBpV
48dAX3WMn61EQbJf3nCFtM3YZOMt5Vs5kOetFnosdRUhkrFNJA+1NgFbo/+TLPl/
OmZLZCItosrMNnif0SHdRRqH9cmFZoWSj457uwQsCzEuh6bDHjkYwiPCFF5QIsLa
zN6qhQYxoNnBzbcgvLbMSkSgeGs8bkhL9UaD0WVSg9/LWA/EWiF0Rl7vqzLLv64+
3g64LLynueQDY0A46q5Cr/M1GZup1JewY0TgcRddnNRXSy8PudZQWOWjMNBtO61W
qsYr52EYy/5Bp96/9iC/ProGzJP1K++v7uzqQMJAvSNTBzMAVaqaSlmL1mZG8Zu4
sINVzdJs+fEdXLE42u+OAxN5Ku68ozGEJAnf1x5HhdRLSK5mVhczhyKw6xEAXeO1
3YxUJ/WQ/D26pwqkfINV0qIzpNKBuBcf91Rte1p4oUBXN/B8K9cNc2n73e18v+0E
Ujq5Aw1ITWJOTdFgYi4sHfyGtbRboB8eDQaf9rnHpWYV0d8SFssuDWKkJ6Z2DMRS
MRdIi9JYo+3cgmjJ+sKNKS26uKfgWibCRYXe3jI/5tv/aIDhCzagflsLeByy3MLW
2mgynPwjVv3N4e59rxVugQdVHpY5SJ2MuNOfxtrJ7xGjfskb3T6nt2jEoKBOO1wB
zsm0xGwPFohDslPtWzWdfch/Lf9DTGgPR4PEk2yjpYqytHy1XBAKytz5wJ/2rs3+
frbt/Q8iPxhSm7Tk1pzkAzNTq2oeDuL1ICh3I+bXhM2eZwYFgA6ppi/OmdT0nk3E
KtF2aNbd0AW/OzO8CU11gYLWXvVzzwMd3djqSWNId+0pJsJwDQNao3bZNDiPt416
9560Z9ClwzNqTXBVHyHDaiVRL6CwUOQ1WhuCixtw8As/2kbywqGlwj98yBCbJ7K8
OTAGmQULmyafPivEeH/GNByE7newhUoqZjIMer4dyXI0fAVrg0LMq5bwetvbjuZw
JeesAgoyjExY9LCMytnXZgSDCZLZbhU3T0bzf+iI4s7MfolM7lYwqCpUj4E4ccIH
8+/NdFpKlXvzUbJykae8GS5fZ2fWdOYE2EUn8K4/ZpEzH6XCDSOemdOozaQFvo2T
zXK0RoV4VwboS3flR5MoOtn0r8zIgy9Dc6CUU7l88V20sHxuYjf/fouuKSFv74Jd
Uvz0kgptjSBpQEznCD806b7MW3cImw5i2enJI7E8JlXbpPNjz7OFx8ja9Ucearof
BVDene4EEv38UgPxyLBOl71PpSDfHRXYhyz6qj3lNk4fFGvOahDRoVUmjasNG+6b
8R/cqnA5MroKhi1Zx98hm2Vap7GHCP7gCWij9CFfc4Vm2835xgBZGhpnsJxQZhVV
tZ31kBTHZ8pDcVWH7ifXTVi2FyRAyOenZjYoA6wXnQVMOlavdP6oIQFX13corAcA
qKGmchXTxhSf/leTxPrnryz8Elee0j9dHT8zZWoOkCQ4mlsrL86IRbR61BF5rd3s
9Sjvud6AjCAo4UC4mI4woTgJnl2g2wfl9ArQR9ExwpKKOKWzItG/szELatuk1moA
UGTxm3dvras5oGz6Vw6b0DkuWPwe2bDPuYyO4fYbCcWx1NZxMQQ0zlMvLrzIN6c7
iVTl8X9hR1gUk/lK1jY1vjEgfAs9PenMdxAmxBXL0BR9KSrf7ywuMK+d+AT4R3SG
0KGVIjC2JM3DafDhHEySrwBR7ueXUXBRkCoVsjaR25E1+J3oxQQPO9FG7Spr0Flt
NTC2wtn4XzR1/3s27hxlTgB2r6exhwf0wvNcZZFjPGdA4G+jUyYlg840Q0prG+uj
hTQnfOPlHoeIY5m8LzqqNZ+3KSPDL6sU2vmN6nu13+L68AX4Kgnk4QhpZePHefow
P6OJ1GKs0oTB3+fpyTFbD4kaIyf+eCxL/jic34EW25DM5u1PzjtiwXcgXe/cnTV0
6LtTQcoVJO8xUYBq2y+Z04x6W45uJ30Rd/QqDreDsulvt+jYw0h24IgX5Qx1bRs3
/wpPzQMLAEs9AAL/DkZZcdmmYTxi6c8gBc6N8mK7kX4xyrrjMxqaJM0Gzw0LQl1H
2EPVyoTa5TzXQxBfFXS9ZtrEJ4Bk8PDJUoJ9riUXsGeY15KWxzg/7elPvHl/GzXU
8zboPkes7hPFMxif0KKN5JUxa9T1Q41FBT6ejyiDshEsxUWxfdaCxxFVxHUyUmKL
SYkggN5BV0OJONjS/VSVsgc2AxF6zE36L3m4ENjDIrAKlz2gvzM9rrJ8U54+hhI4
3fr1TyEqlWyGd1nNVdhucWYNk5KBz3tUuMv6S5VlFfUHaZ4vWenSExxi1d6v3c8q
4TZmwiq1VWv3XwaQiFfzFCSVTEqFzdh3u9NmZlC6eg91AOAyoBET6BGytdLtbueL
WOgehui/YwaBD/Nv8D9kB2e1j69HAaQmP8PV7ScLccNfT3CK8QLn/tJ8YjDi9Mjm
AT6yKI0ciHPbW95MZD77z9QWvHzALMSKc8KPaNse8oXf7XIy/GOISG3UAbZ7yGDh
N++xVcCiQ8rxN+Joby3aig1uFTbpXW6eNwd6+hN6cvBKKgD0Ns89I+dm49F1jfwj
Mqkfw+AmYzCH3VLe0qO3Rr4ABmqRk/VWpSJw0/vBt2wydaT6Vz6RWnXj2MOPA3H9
QQ7vFVNklEuP/00DACs5Z7X0XVMMMJlkzv01ZGtctfk8tCFhCaFezT1TIIuNAKLc
oBZhC16VcINDTk/D2ktGPpwkM1p7EmY8S52T0nPxdeL9JWSla4rIOXadT268TFoJ
bSksG9wb16blonA9b1bKWQIOj3STXgjBA1OWsFuNXl7mQhZ4PmDqQFM7K+iSzpld
VF93cbV6BuMvBQmxA/MyhbFLT2wk2nhyoDhv6a5w0F10M6yMoWxdgNm1OK7N/0fg
BeE2Xw3M9w2iCngiJCjrny7wHvwYU8AEH65ci4gegI8cvoo8xxX3FmhYOR0cg5e3
tkgPOIu0Guf5ddwAqx6HhxBzWnXIVoJNsdYAib9MPUkDPkKr5L2axRmPn5x3oIha
/zhGx4gCapmZLG47aoskvoeEavwhhYgKoIq4wB7plAKqmFQ4r/bPxohfKR1D/H0w
C3dHO1iaZzhkmlnyq7wtv8XQo3mABN5fIHzoaPKNo8cxLN+dD7QnILIghSxTdRwx
VVnJrrAXG+BUyGYsZ2FdChJDN4/b8y9LtbACkYH6qFlloG9ueTStQe1VVHZf8LT5
yRAubB199sDYXTcgv6PottVuMJk+fzcVt3t0XKdT3RQz9EHJPrFbDCSywQwe6/un
iFfLi2ZXho2+Zrx/mVG6htj8Ibts/V6HirdB8B69tgQwyDLox9cDtMbF5EsciGip
sAL2myMCWtwMB1pmqC6W+pV7G2Q13WHzRmifkrUjInVtiiNmcoZdzDbGnW8tBWqG
wgsvS/GxsRYhworEWcL5Z3xJRNlYLKzi9gdB0dU4l5sRqrWg/gkKU6If4IaYi949
0gGoIDXWB9osuTlCduob1A4EmQUrZGpzzls5ss07vPPWRVeZAJGIeTpG7ct/AKMF
Y44QKybpQGrvP2lb61yKJLUTAkqhKbKrem/U0PF7y4EZMzM2Cx5X4erszgXRFimD
NNerimnhUo98zwLg4ZrBNKRYH6CV0C366kkSP85jKUBqYDc+E5VvaXoTm+t800fZ
FGXgPobWXKImLDtSs9+cUkc0F2p+Sgxeln1dWvIuzQnZ5LVGisjYPs2H9tc/hqSS
m8NNoHRAOYOxAkSHAepNPZ3KEdLKhRlR0mnU9kRfeH6YFv5Bq+lUvCry4Xf9ILVC
sBH07/n6nnAhKgUejhxxKyreQVexH3fFkghdE3I7uGQ8f3UbRB+yMUb5Thn2bPov
CkyaGmkEWL9xQC892rizdk2o2/Xrkf8iXbjoSmv5boblH+FgoAsr6wYxhc6ynG1J
IOveu2tv448IcvEWLANoV7CEU8gHi367bKo4EhmqOueVAjb+XzLF5MyazrPggVaZ
ZdwtW/rLcG/tdPZWW0kFH1LJw2pxyxGq4okyrh7pdL7/J1tWC3H13n8IxyTJwi6n
Nx6pLCPwp7Q69tSygXkpF383l2bDuMOo/mAnofECbNf7u/MZpFemJtGiwryQQ030
8IIBlQIxG+sDHhZo/aOO2KIffI8ZH0nzGORHo7JjTjdBXtY1VWt7gE7q5NK9rTTu
2ZVE6jxYBZ2eE40qIoecdcuhfJyjpSPTs4YtJakkhdkH7mD7/FYwxqFR+Di8Kr3K
qbitQ1jmgCcJIV3wqFrpcPXLb+LttBLXS2ncnSo7e2c1mDNb4VloIBqCIWqhw2xi
ZvDs+pTNBMNsr4tuycZuDAfK9j/wpwIox2GQPxve3MVuJjIsAiCjlQl9e0dEErx8
cpbYDw3I4V32yFVivD5QlhT/CYZMsXzC8x2b41Z1mE0ayGRFpGmCiUNmZl+5Q+IU
JVhoDTh4jT+IE+SBONX1GVXilAHDgQQDG+UclNGVli731MIZS/3ft9a7i5Ub0o/Q
jc4n/5ne976MdvOZdEmPCglh9pJGs8/jpIQUdP/e6VUw2+5ejG/eFAWyrcRzAW+c
4ZLYVmFrPPQbN53nrxMbyuMvrLRsl471n+BZeUunOuwmFJ3LeEFE4udbkQy2NEGT
brhW3t6P+2Z3nXNAyACNKJhR7Y2+2QeXmCOevPNly9YXaWdLBhC9t5kCbODHtggh
Hc3MQjHh7skWepF8Xggtwh6P5M7Y0203rxb+MZCrvB5azjE0+fhpRWmJqiazP/pI
jX1Y0q5yLuxCKtkC/mepZiydxCl9zJRi8K9E6qhdkFepv9HtVp8MW0/rDJ3ai3RA
zjmx+YUE5yhgpTXOUJj14OhqEIU6WVP/q/BZH5r8vmkJJylKtIKXmF5kIDzBO7cl
AMZxqjvEWLBIi0pH+rZBqx4NTRVnVJNFHofUan8+/q9Z55jgTPkVFZ0Lc9ja0xki
eZhrl1tgCa+OT4COmjI/zJG8QkMNzbWs/XOdyPrBbjLHsuvGIeT0fLgDITWDlnM+
HZPO3g4i30M8HOQqapon0ITPtskg0ApdE4ZfVlX7c+akuYYmsQ8hPEa/5hX521zF
6gF/zXRDoRrRs8iACS86+THzYRTafXH4X7cu4qDd6g9NksJkbviJ/hucXqb4JMEo
a9XpGq/TutpzGA9F9GfqDxWf7+NvtH1pEHdR2neW3leli5Azcct7nHgXBdSK9/nJ
Dlq/7SHE0fdgC21Ubr1UsL+i177tTh+wTI3gl1OPTdoJWDNW2mBgxTBidQ8rQDIr
Z45Q5Vc0Qr6aeJTB7unI8+Ua7jS2XWYzJTg9Cxw4067QzdLMiQhGc5i5PTsepvpL
yz4Iac1vaVGyo/i19z5vmUEMUg3unuMR8TrRvp7RQoRskIN2qfUzIIf4ar6POVlL
YD8fGT5PTCHqC5dAa+SgssEjN4/HCyU+CCMSNM01fN4QjRomVDBb/axvlTPgzTxb
c4OMOnNRTLxoZyIcvotRERNex1ksIKzNcvav9nkeHh8TMp+F2UdEhTqkGzHsxqFt
+MWGQvm77M0XQohu6J90OpRnAAk1xRcrOCrheJavFLWZLtiIcpcFGRF3+Y2IB36G
ZZK5WvAPaq9TbXARXle7Jf31iTjgHUabuqEqrNf1mbqj1VP0wxVOlYA4jpbJWNQ4
L6beCagBGCVnjLP5/GgLsHhcFBuNg/bmU3EscGNzx6uYqlkXV+TiBFrkD6QujSj0
/7QjElp0/Z+RNjgSZZRnm/f4DQybiL4cbHIb9YCOwZ87T7z8YOSZcwaBUtfYMNXg
5BLnvVlJ9CVxeXGtcYlJZ3/HNReN2YeZxvIMUzvt1q2ZGN4JPPyN0ZpLrJ8Qi+yM
4K0f97DTk/Eslbta08aXWvF4qvnwF3+RXfln0QAbA/R1TE6AwD2ba3B3uaROgdYL
LVuWkKXXsFbJpJNFhAqSdb66y1PL06yo0viFodFZaVypGbaXEPZOmW+5SH/bT7bV
jwE2uwi12FL6I6nEfEoxER1pYxR0tm209Pnug9SQnhu2wJFp3ROIQtn1DXp4JfUR
lz2gEw7WvG0EqnrqbgLky4LKhSnk4F+O2TMUKnWTRJB0DMeUBmZZKepxTY2dCZud
D2lddFV/h/MvSXTlfUQL1pNhMjE4n4tKb+Q6yetqeJ/z/pKvz8Q/sL3veU4d4JFS
I0ys/crgajSxPoE+d72hvOwQvYd2dPR4uebQCoqZwoVz97p/F0/e135GJM40NCKZ
FrH7SU4P7XgwgiCENKbvqvL3uT/zHhk+cGhXztRStn3n9JeIW6TljQ6sywJjtPkM
25nQrXP6kjA1qqm7K7xyqVV74G5RkcDYlm8KB9CNw/AAvYXGjER09apWKryArVTh
SPAmX6Jdxy7J7s7xk6xzsyD60yPVW+Pj1ks4MXs+Jq+qTNs08k2uH167QMmonctY
4tuODjibzARRId8vGQ0Ylyb0dD7SJzxBjw+G3c1OJNmlRkeiyot9EBuzFjLg2/GE
hh7AgWHPWeo0XYFETplR6yEQZ6DDk636vr9HVTRfxyOll9YKD7wuSHTyZVq7Nenh
hqk8w6ic6Lc92zDdhEhC6EWB2Xwb+qKQ69lrk03o6DV6z2kvtWxiWyi8mLEguxoI
IyEsntA7JMIrWyCBtJ6Z02aD7wHzxDIyibZUFLXC6vHV4Ps6lwy4G1uggv+G9H7B
KPZzSwlA2wXN4UZeB/M0vEyrvxJVC7laIRIKYaLirruQGqkGiPgbU7zIXlEB9/ZS
hBrMr7dZlEcCZK0qGsgwaVEzE3SQtNx+hLr6x3OXJJjxCfRlN9ABAUQ0wPbum+mN
xTsFXX7Tv22pHGQ+5gs0jtd/lYD22gy6b6Q9HrKO5Qq0yEdYbNMeKe8qLiBkh2X3
ML6ROX1MxTshRa03NYZ9FQ/wwTgeogRNOqRkAsc9qvz+0JUNBgI7MZNkcuPyUmWR
AHg7T2DnoGvxykQTQPFbfbDUToICDcoBKIPRtVF4aRYXts1WlyOrndQBXewh/ixN
zXXVZ9fMLlITQtD5aXjUlqyaN8wxA/oHaPUZQuZLpeI0LULVRaytutmvtHV3p1aj
ugAlLlFU0Bt32cwA/5MRSza65xnydkM/hXmaWujQ8mQmitQpzjh9ByDB0g1PT97l
vBCT1PF5Qr16Z16gHR22Bt4EmD9m5GhPK1rbWSGDRxuhYl2ffFx6o9sjrCHti+zH
MBfYI+d2irBDqO/s1dIa/QxvT31laJ8ycfudb/sBTLlgVcdNU35Lusjn38OpsuuR
vfQaCfqW7l76+O+ar7yHmFAN9z6eauel5feINq1ZMwGtiep+0ZOyyg0a5hAWWwYr
co1oQH59vpYQWbGJx4kXjfNNIfyVRXdpc39TtYdbQ5Qu5badxWyGCqzw3RhdsG8x
zm8kLO1GkwXFUkx3erk2dyQULX2bWmviUufxLbeBONcyYEJxctrlNewIdqdt9tsS
2q2keQD4Ro+E8Q91XcsdC9PaDibN7vgMtEbcubUeR//bSm3qVEc2VhSnCK4bkmIM
tLQPasxHJOO5J3tbi9AGlCYw64+ypvdfyMjcQOV4XfOvucNa/TfvsaQex+PXPbn/
rclhJ/HJq+cvFu4SWqM9+MlM8nzmm4KLli+868gFFE15IQntSQmhiuaW14mrvuBC
L5RMHtSukcUHXpj6HWsr0WWmrAeUyit/16Yodv4sz+t2n6K2n+47riRycQaBFT/J
nDBP9A0WSWP1XvETrBu4eRcM4BswBeR+DXdDFebHvdi//5KLcnMqCU8hhasJXDMX
v6vCDHOnpQETxO1KSDNQEKIWDHPy1N3/A/Ir4QhdQ3ENx49g3TqFFCpbqhoCL+J+
DPDSn9WHwHWjLWUmOzvc0kqggDzJ3hJ+fzsBM8TTtmDiad9++jDqhHlorFBI8xZc
vH2+sxQvV+w6Q5tLLTtoiaHb2YHi1Wel49qxQyq76Z330PjGRxleM5+KThGm7YW8
O5/oz7+LxhnVy4EuosTDeoWSPL769mgSPUTgMRoWIRZYoDFRMVgxopLOcoNxpVgM
dH7+KFCMLVqiPFGGoSb0R537in6WYBR92+gz/2Rcjufr3qausqdjOH0RfUyxyVgm
DzF9bbLOy8Px/jl8vZYxp11eMkFayrHDx0GzmFbQZyYwBpWlgB2HfliBDWarpD56
De2aLpULltAwviGBc4JpfA6tRZtV9W8SF8vTabL8KHizWGRHCBc1As6pLuTXH2vy
s8Cc+WMUzyCbVfvxJrAVu7KifJM8OZYkQLctgk6ak1jCpqGLIzkdlmraCarJbgjy
lxfAVeJ2kDnrQZNoaqewlIQD6esBkoi6GqgVPl5kwa8IN05N5TnjdKQpNtRiYzYc
K3r/fQ+0MZdlktHEdmClfqSp5EaY+E8PIgMAjTTfQIi557UXlrCPmKJwQbZirbpi
pDSog47e1GRLQKjJkP/QcZBRWwEHiKGWKs58RboN0JjPeTRwi0AL/glKjneSBcGN
IajOb1exc7M//IPqJHdxVU/j6Pk/I8mqksuchbfZ+Eg5333FwHmawzG+HGBkGbED
c0b8cWAShQGYPpagTZTR2OlPnNaHXYeEZ80wrNf/ZDMT1XgGXx/rKcjG0l7q6lLm
rJ5evfXgmbGuk06khCCsiiQ8H6tlev0rlPBl0kMJ0l2BPqYyGxFo55Cpi9u6XBVj
a2BNO/wPEnGuWPW0zLo2LsV8Y1ClcwJIssrlMNdc2RoKOTcdtBy8dncyhq8Mfth8
2zwuwgaTDeqzBOYYf5D2eFQyQ+gQmj2yOUIpbWXy2h6zjFGPPq3tVwLULk67q8MP
+Jf4xtbsnZfgKoNSGzZi7w9dHHveZY6p3nEBPkx1J1/EYUUq/ECqGW4t5qRbxQ8U
dafPp4RPRNTFCeQk8wx1nq2D+4Jg/Fb9YVbBm5FKHNEtwq/Jf2KQNEGWzohWeLWT
Cn63nKQSRGTr6IFFoWlWtSpzssLjdLLOSW+0zaTQ7OPp46u3EReyF1OHN2SBX5tV
n4bJZsBG+Q7aSoVApRFbrTAaytwc9uL/ZQcX3VZCcG/g8EUjGKWJJzobXMovKAOa
EJHI7XRDPWPmYCYochU6r+RXq53PnUEW2BvyDM26cH3UCwNc1ytZRZBXQT4DmbJV
jufmJWlD4tb1MJ8MUv8maBXT4SBXOf9R3CSKe93aGsCmOaKk+LXNi4JKVFrOPtyP
DKafp3i4godMlI0/ipCFPq+n3YOrMYEd4zwK3rEi8ofbs56XamYN3+36kYcF6AFe
fTysdsgd+gah0lHz9IEtiTqnQX+fjx4LMFPTT6qyfMTakQEQUVnlcvzXEUAsC4vt
hw46p/9fM5Wyt7pcCXX1Xc3fqvoERNr5tG3Vjsel0nx8x+o0oVbMrSCXUvhawv8C
na6zqkxoD6h9zVTRcs2u/FrM34cq73CiCBMCFqE8MRlY+g4HFVeuf1UwTsZiFAWt
WflsAdAdNiqEr8gkW0gGoJ+xPWV2zg98ohLy1bCXXEu79jXHwaBYHqUbb7dETp0Z
KqFnLwIo15NdPQMf8tMaA4mcLRSxxAgTI3QsQeXsi/K1jM2UX73pHDgsp5Lihx0c
hxT+8NcYzfJgUVzyd5qssvE1t7L3H1HDoE6oQtOWy7dHC8P/vA/0WV3GfRVqUcJH
mMN8uT7HSWzVZNUosZkUNwbJsak6lIlXkGX2VzPxcAnbivDYIHxnQ1yWOzH9oOSU
9z4PR9+vUZK/BhNjHAPpIXh1+9WpnOrQ2fhxqGXdHpgHta7d6B77r1FI1Qb44dps
pEDCPRKtiUX8K9Ae26ZJ6Q2grLnZxoHwUMJ58v7S8GtTFwUoplO2qkWLw40vEkqn
EEZDRjedsHw6UHjKTmpdKI5hMLLg+1NvHEOo4bOjpc/kVGKUXnsd5XLHm0W2fwPi
+F1aorbK+XConwyIzUw4GDaFmm4imKFT42qmCQo8g5CfYaOyHGo5j58PxyxaKidv
wySfrZpTFcd8Fgy5keSUo5ZTHXLEHzgELPU3oOSoK8Xd5FWo+wVugtwoZO2XOhTG
2w7FOY3Atw2bJSO8Vc2z8f02/kqL1XpE4rYAOH2fAO2rC8E//r2yExqYa43emZ/A
23Y3daefnUxNIi4AMVj7nznQ2wePbLyYzBNGJf1ygcveZG0Ow5W8bwV1PYDc9PVA
QslcYu7QUAqObIMzRIa0Z2gKbl79jQQUnfg0vs8YZSgdtfJbk/Mxkz690WntBnoy
cGEXX1KfbCkHyZNvFi/u3v1vquxIZNKt2M3ydWLFSMFeN7UZIaEG13sCdP2FspOU
lpd0zqBo5hD52SVjtoPRADT4GmKFgmQhu5LgHUwEC2d0bpHrf1a9RE2zQiQ+OiB/
n1nXILw+tRes/lva5nxvkPLrzs4ryG+Y1K0iGX/Snx3g8CSnjvjqrbpZ1uCsBx4Y
v8MOvrtuPIUXDtl/7MB0yMwArjf27X9BuaZNYmQgw2mq06gMmNtyMShio4FfgBwt
ubIcYDY8kL46J2KzHrRAxMcOHunGEp/Gxyh4jFc0N0Kj+1GK8DnQwin/dZcXGcOH
eAL2uKsUxlpV70ShnptuVxuBxgGLL3q4EpHpBGM9fwVCjHexGAIpd8k4W+4WaMuL
gpyJcT7fmnOsiT9ugfpJuxOvhuregVFY4A+rduMGZ4KM/EkJ0tpp7YCS6bbWUe3z
N3bh83g563Z4YsYJw5+a4LT6LghV2snuAvXRY0XPKKqRtQxZxZJtNmEEcDGMrzs5
jKTlixbH4teI8/AIIH6cWHi61xKdyg05+t0eawzeiOvWvMh+5veQzl0FHQm1AaDH
NA4r5Cqr4eY4dR+G8bwAG/K542GJYIJqL4700p32My+PgCxYjVzrT+VeFQuxK3jG
PAcgGMfmeIJu6R+XaDWROzxgUfz/Fba0mWnikIMnzk9egYw4DZTGx6+LxZa6Cz0o
PnmZ9RsJmfiAxJUMXSu4ZLRnvpeLQ29+MzLk6c34DZTFJ4LqvyqYq8OsTwKRc4dX
/4MtXh84PK6hG7zY3obYEwo9zFyhVQ1zuH5gqYcldG8Y+0vWXb04twiXCpFl/AJS
rO2FuFXgk1Onf6YwjL4qiDruC1kKKTfbeoQCPLoxm4AqVwiFOgs9KT0p37EbZes+
LRpuimqsLDdMtwuFMz45dUQOknDwn3wvd6cpZOKrp660agVISgaUTQZDaeEDoDkP
iSUrSJq25B6gwOSYqKkHzQDuh9C7A5OMerjPnmn2GyoHpO63qkdjwjwFYuRB6/cg
sGsXYA0E8qTJawzmLTRA8fwWbuA+arPzWwRYqJtINr0rWovDK+py3Vw0CtbrqBty
Slk6Ywwik2C78vJjtSB7DRt8gt3eK8+Z/oT6VyE8I9ivuRqMPH6HEnGnCCxgYNlT
8LLZa38k/YDLQlSAoc7R5TiaNeLXoPonOtvDghuQlsw8HVCtXCUBgNqZi9r8/+5f
tOmnxv4Qp/MdgqPlSk//SsmdbQFjqB+wwDgC1xQ22WKkav90/FStvYTE0JN9uham
p4Yf8YOwmi7Wt5DD2GcNa/fm6GqsRxPGiq5cXGxSqWyMe3qdcgeL+lV505oLpKMe
DVWu87yHh4g58dVpGrovCf4sUqT9ZjSDJb3IOcVKX/4Nhk8ndp7GyZPbySTK1Jpq
TtCPBW0+i7FCjUw16FCR5YdwuqKFsUqSYzHOPM++SR2mHqK99ailuiWhhJoImbu+
8NE9gdKjPYDqQfjKpmfGGILhf1bS/CsVTf2eA/uiia8zbh4Kq3NexdkWf7iIg1Kv
yGg9NDBqIln6ig61oIGRZLTICCYvpvczQOVWPwreWjHFeqmDk+tDs6wM9VyiuicR
Ymo5hbUXtQDuFbv4XEZYvC12SIz3zzG7+Qz+8oL57AnuqywhRFwAvE8YTOVK7KeJ
PgBz8tXM8Ecoi1HDKuVZpMlGUxw6Qvr4AkaeX4WPNMo3nr6C5IVaTZTiFEaL6/vC
AK87l33ZVR9hbXlLTQMcsamt+UlwxASIi7A3lNY2cJKzkPtXxXv6Ka14RW6MsiY6
8hSSnG8Cv7KOebmmQrX+Y/zgBmKFIGY7GblfcGq1ae/xPzsW7TX5qLAe36de3HNW
pMlcBlaEylPSPhowfU77kViVOYWDZgx9NvxT08tMC3o+AK812J6NXhDxlMuY98A1
DLzOo8kLoB56Whu5dbhmgkHOSThwA2NHLoXxL43WgA9zgObeL0eMj3JL3VMqAtq8
46HdkoHmCz79BCkgE1l2TZ5ZEyegQDhFXaYFmjQDqsSjRZKF+O6+zXQny+qSdg2h
Bm+DTZYLVeYXLXW98U94B9XMPw1TDoASlTQUChVOvLTmrqWiw7fejy+4wJhH3qZM
2kOMMtNNobCnC7BT1o9j7qU3cyCT995nfoKIZ6+fKC46Cn5jgy/XJ6E5uDY0BAqL
QdwmUvLmgJLCmdmUdYsg+HyxPMEGQJxFGhnCRutCb1Am4k8DEZDrxN+4sqHV5Lx9
jJXaPJRZm1k9im84Np5D/JgOLWhma/ZD7AMCtxeA8zwh0rrcaPe0jbptnIL/f4PD
shxJ3rDv700IHPnyJK9ZDFLsxR+fcdy1nElOmt4layhytjdD2v3IXr7sG+Cf6Ygx
HjNa4Lf3Frym34kQBx6IF17Yez4SI45d4aYVrxKt2BFp22Z4Mx6txuLv986qPTwA
jeECLaEIQnewiYBQop4idWF9ULnWRaNfHzV/kdpuM/42mhr0gTfnpca1XMjqn2Fh
CanmrbDWiBeN6WhUcRkJS/RVJZU0DEgSHZHwNrLa3dtf8KuXf1NR5QLCZ/4PZleb
IKKv0JqhyiBkRi3dEzv/Y2G6UWNkXBFOl5Z2NBfV+cBbHLoYQ8dgCliYByDPD56O
k+/v3IxD2hZx+E+S9J6h5RGJPrloS42k+KcRLyDaG9eb77jFFFA1riLM9VpeAWy9
a+cErhFLJOKlN/AqGcy5qWSuLkqGl/sameLCE1ha/RN0Q7WCc8k7axE7l26GGp1B
bKxpfJaPQAiebTYhhojaCmigrT7EsMxd/FTju1egMR5W+A/eMnpDI+4ZYcwTWGxy
esZFZOqO0fk9XId3F67HB55tRM/iqjPm8zh9QmlIsA3M3trbFWEng/2dMn8KSJnL
j84BiHPApjrOT5eh1uDkpIioZZAMyDxi9QNAgX55D15Sd6gOHHsYJ0TTgsly4eCL
lsXJeZQd4IRc3XEWamcmFIxMwVfjmUb9dmlfFZr7LVXND60zfTeX1hYGV5O7tKjY
ovd+xO2Aa+hvYS+7jmXAS+t47693mAm0vRCTWg7l5pMwWS5e79p7mRC9yUrTimeB
RS7G552jEZtzPPaOxzg8nXQTSykMQD9OR8BrGYpIUbguAUQaLCtB/eHkJlqsuWc9
9ut4AhPL7kdeyOgzIUU96vzJhLWVPOzTviMexcFtK1mqAJB4lpy3Fq0g8u+tLihV
9hTiFusB8u/0DRlT9xV3qH9yn5EmX5bSY5c7TsZ9C9zL7t6k4re6iCt7Lg3HQrkq
LpXTriNn/yg8fXCTCsDNoWvNOpNp/YK2ax2j47X+iJBio2LqS2inj/rv9m6pwGOg
7MnIeV0IPZuAnXg/8qQWf7jZT5iPaHr9OG3bJ03PSJNor0dQpf4Fg405IEObsbG1
oojOBsrUpzbAX8hCVOdNm7pDVEIYryyKfwY96taeeh3pbOdOVH13nPt85m0fHNO9
wrFILM/7Sjcq8l9xLSSLX/QQBAlz+TD38y7D60YUBNBfK8SelIyad7BIvSB2qiQG
GlUxPUvR90GQdIC2lKC5liYRYQYaLAfq+6fAuVCn+KDkXS1jURcrRCLLKnD98H/1
Cu9tbArA3TbhWuw2rblK1u+ke6xo7hejHz8f3q5KrVLZHAPgBY8OQikWXJ3g0ANo
/ukiTIZql3yhvE0ItXMhHHtdUq2VWDutbNRegdvDh2z1xHCHDJpoHkdAFfA7EWIl
k8iZhFUrNxr/EJkYjBR7QYxWOroj4+BBEkYCYVipIYIzXAlQGTpcivv5Jdp6vSp8
gUqNeM/qR+nRGGy0nIx60DB04vK1zRGUyQPKnyR3+RG5OhlOA+BWPrEYqe+Lyzkq
o4uqRUdB/jjCrPoQtS1mF67OxWlaDXAg2Y4qcj7e0XlOLqVhQZ6i7mzr8i3MW6Am
rIvEZqJZViadj3BceFVOVu1lFklTfjee27VnwMzinZtWooO3vqLAiBm6tmacwXET
uEfvr5M+dopiV4wUf6tgJNg2Ut+djgWc+h4H0VQAi62x4+5Fbh4VtEJ2CienwbPo
W0UKBGaOFmeoWbivGPlUiwKsJWYyGt/kuteScTs7f017/YB08aYn90YefHcApGA9
ps6+b7Tk8D4wpKvNfcd8xdqivgrrEQZalmfqhmVqgLvIIxjyCS27LTSm6E91G6Xl
A1pDConVgrRi6FyExyye30meIpg3fwhJEgFADiiiSXBzmguf6oRN8AJtztoMI2VA
unAy8bAhR2YUJb5moU8I74TUVHK2BEqY2BkpxysprLusFBCF57s/LvEUTK1s5pIP
DGHQ4xND4EllmvXjmohEbaWo2YKuJ7VPfcC1EvgX6QNxsCWVDV9FNAzrUHA5PeSI
oyM6HWbXKHaJs+MSEXnmB9DK5axtxUvjIEvmvuwkr+TifWIc72i2Hr5/crOPQMdN
QsYek/2I1VnyEq+N3AuIQi0z9csAv5I481ZzEZ5Co1LANP/spcviqkZ6qZbePAyH
n0FKeWCma8QHmc8lCLL7MXEFigr8iIwrddTGgTgehYEh1mrNpwRm0mDl9MSmzqtL
tU6XB2z3wdrFjsymXm9GhBwVmj2c9mAL8bhFHHB4m3hVMVfRzlNSx3oez0s5TKhG
skqyYMP194VFUvYczk6wYSdN7Dt065H9nRYAwo7EuOzOtSJdA/Dmn7UW7mDVVZkP
sNzgXLXoThnfSvrKj5pzJT1tpYUIJJgw2L7/XGIzLTwwHLlwQKfN32WcnUYqb4R2
llk/Wz4b1XsJ+tebSVrvI67wa78I3G9wzSq1ZUDuLHwWpo4cu1v8IUeYT30wsYMT
TsuktlwSv/qg5EQwUqorLx8xnRXrnodDW/T7oqStZprxQqGT8RZUnxb2MAqV3bUv
IRm/VatVEHVwRYJCoWLDGvkjJvWPaH6+ZVG1RS3dHUeSXcVbQ67KAfjAavOqlXLq
KOzYkwzeCo50vdYyom7atERI6ocb4D6PqM8/d6gDr+UiyPHyLX1InfFGgnD6Kg2R
jG/mAmJJVU3/iDndTfOdbUBwWFPmBj03YEVnPC/TDySM8Erya1DN+p61U9qDXi51
weZgKhcM/1lzypp6ABl6pB0g/AYMfdg47YU6gRgY3goW2qsXNoF3XD5cMe79AU+4
T7OUFPPvoRsdTZtgNkKLSZ0qvd0BcGP9KvFc1sHFEERT5ThfQmxSoJFFIdbOGc2B
P5JOSNop9/rwmWf9pCRu4yGNfwxlai/HMPgStFQ3DMtDOQDd+a8b2c76SW4ZzX5q
GdJqw83yjVRR8F10N9p89GUy6p6X+XI7UnxpFV1Sm8zLL4WBcoeqHrLbHdU7ew5m
TEkNRdl08dxIEmFXtNhkY2pm0SSoz+L8ExNIfIeARnokjjQDLk71Ie7Ha7koAilP
LBjreeQ9cUAGnV3+oIHqsrOIouga1s2nHxkjqpuKU6wsV9ybbQ4XjJe2M7UqRL7L
SGCO6DSB+ACSpvVueA4gc/SrZpJ6CW9gZlNu6oXJlbSHA7MHvZbpOhpP9F7lQQkd
kp8jzw3kXnEaI7CYYSTMhEs9RANUjuB7eSskHNgBsN7oLtikP6h41ln4DZUHk7Lw
r0kPmtv18m7E6grSlfD5FHj0MlICTgG6TkHRpproCCU5hWTnsOZqL/ZNxKsaIRIi
Gz3VwpcjQD0STrhfro+VdnS6Peh6oTb13SE1L8KteA5p9v6o6O70H/P01u1XGqI3
l7VneWuOVY+We/WlD1uQ1M7XFhj8W16hwh/I+woXm1bybqdkHyTSlwYPNkVM/cCc
j8yz+CNvUrgxJvJjMZW4NSc6JOgFxXgD/G/l7X1JLYDj6qJggZHdoDuyuFXzkRoG
5Lr1Zfg2sz+8cR03wYxQQLqYAhqf/+xQcpaCluQpfslAsJWhB9a4yv/yQrm4UK9x
sqU1x02dfR6O6XRXMs91XJIvSJ1Bso76TOqdMG8KhQ0M8QmR51RYJ4VFXBQFGrUG
x/V85KbL4xqXnKaL9tlWdVWBLAaUDeWSi7ILiDnQVFsuupDCq6vGdSv6IF1lywML
miS8V4n9/4QgqSqZwXpxqp/ACKpO6SQWGIALTwtJiDevNz8X1gRRw1L9hOHqVjX6
bbYFAOllI/nZZHXdQ47P/TSoVD2QP2y4h/RTnDDdqYfaSrBIJdRNevkODlKEMfCl
03eC85gmATsav01l33e63JhwHZbR6gsDvlkDO7kmEkMXQ3QYtpddhgwDrhIOTVUg
yCAVBA0qxqWEQmxowjGs19D/Oto16TUaaIn7Gy3Oe9AERk6nylPnDBJhno+FHQdN
kYN9dtIDsjxWyMeNCsjcAOnUag9aJZR2JSPTQo4vEg/EDqSGPMZLEjAjFLZya8QT
A02vKJmjlvOXDKuOc+GlzPMPy0UtvjxMn4oSzCybN1Yr2labCofcCws4i7QEwHQP
40QroKOZVwWpANwzpzpFy+SejwcfdXy7zSHcC5Uq/5UHuHA5sdpSGkuzOIqYfhpv
0ZhMnIZuN72WrpGsVkqfqu82aud+TXC1S+/tALWES1D77/Drds+Ou5rxHN2vNyCJ
nirrDL2nNAMKPXuzmQqWpI++F30dDSoEJfVUZWbTTqkyxfoIK7+/IVQa62+6maGK
h2xMX+CDWECJ+zakg/idqUvcRdZ2948HhM7mDmfEuCyR8I1T13MI/xsSZYdMHmBK
g6HO268WIRVT22iAP5ZAoj9l1j9nBZn+qe6EyxxsyEsASSDaMlXU5qtVNe/hAXEW
Ldx+WB9HF1A+MrQOBbdJcRMhsI84N3kP4hZswA4EwYxRj+aTl9gEx0z4Hr24zGBq
rhkM93CYHay3gasLc1NaqilV79YgW39byq0sSRUfRW7qrlJjmR0TQSHrn9ZHZBVv
WUjrpocvXV8NGrSMdBr+9Zvd7/Ic3M5vsFvHcWvGyMzS6gxEsZNjNErH6rwjzdqn
Om1BIExlAJeqZNFO0zl2ZA7C2+dM+htFTEJhA89MF8ThXuVaB46EN48/OZSLlLAW
SD7RKZ4RBFjwPCo1EKQ9IQ9Z253BEFW+rBROmeE74KgVPsgDxzzLftPT92QlNVIz
iyO3hfHF3Cvha4A5lCMufjL1/DZaxsaeU9Qe8DR8diGDZKdLd4YHQHEOxbv4fN1m
mlFziQd4/MgkdQxqn7Da0PAv/2Jnl0XwFVF/29oAE+GWg1nQKxTA386Qd5xczS3K
P6LaQU09ukyZDIrLwsNvAVvOmNcM1+iEuP7920rCweblWoVQH+f2/hmXVUNChVxp
c+VYgxYxsz2YeIlUjbgeiGCyrTyy84PRqquiZk7O6LpaU+GP9mGaFj8unQlZ48vU
vPPIVbGUo3aC57gqeP+ibrZYCfwzho+b5/+SGb2jE4dS/dMuklzkdVed0MjlIT2j
GuGsM9qnYP9HARwWJ/3Vn0vkC7+z73dOvK+Sr3apu0eTmA2yVfEQZow3aFwQm9RY
dX20TAsn/J+1NxiGIsMDQ/ZpYbuvrptYCBO98J8c8vDkRkmBq/cDTXhgMPN2nDsn
2r9mjfntqsXTh13bhU1jtR95hC7Ia3C1YiRQRqgSAJhe2dl80q/8us0kgrSHghSM
bzip9MxN10gRdOfRH2L5hajdxSSEwUv9ZTLvvrVfJh8KDzse8l1GWkJLat+MnW8e
eNKr5x3RQyXifQH+LYZJEZowWQWfJVPJn0I8oV17q+IPFlKDiSys+a5GI8wnqO44
lnQRpDpu4Zi4GKI2KyJ6r+UpuhbxIFnzJ7yysisQZtLKau3O/sFAW1MMUto2Qjhe
n5wm3qp/BBMuXWCu4ZxtV9t01NrOJGknNm1hMLKSuz2S4X4OI7qx9axwM9+Vj96V
aaynUbMuUidKqVp0ktRmaEsLCCTMVL8cwykqmgUSradNMp2RyWFMTkgiFsSijSiZ
trUCZpv8ZZS+WYUFvehEKIPonNoIlF4TRpuht0Yats4QlIeqdWVA/pR7Y0hASZBX
xF+eKBfuLv6TU16Si5Txfd2fJNggE0iD7eim2yOhZHzWbhrQSqHE66ydEzYuIGPM
ApFBoio3oZ2mk2+HrxxGjqUIgSTRG+gkHqToliK3GVA1CdKYMnGTczev2oRpwEJD
oIU7rxPM2uDE84tZa0Y3xLJN8Apcht565RMOD4Rq8zMmG5we2ZvSPiTmMmWxITJs
JPpXL0fRT00wkR6SBOBqk1XHW2PwU2hs+7o7DiZLqKFn3FWEDnbbH2rMtbzOcl74
SvmtF0iCAft0PmiCwIdAwsXYVOBjmcIycUnLBXecvwhv/fbaRn4NUHToQo4KLxDP
3WmQiQ+MmgI4BYcRPulyupqFyD67H+8wca6qTk8yH0ascH8y1bl1K/tHPi17D88Q
A/+s02WA1l833bUiU9c4WBmdRttkm/ES/Qu5FS9aizlTNhl2YBz3sbswWVzqA9rJ
ivITB3kAVSms+pLb6oYLhLtULPO4iwtcbEhoe2l4z5PdwyCJmyTEXdSNanh+tyVU
SRzTpL6W1HEiQsYZqiZV8FqSy/uZd/hbIgqmf7A1mg4iU66c3NGgOoc0/6p26p/O
5smubTXyZXXv3ssJ6x0Xikg6QNlI5xVWLo4iwQ/aDVdE6JRV/mx5OYB9HfmmDBEU
OTjWtm6z+BEbVCZ2kKPnuramsOdiWEUBh8ZmdTj2j+yiC2Kl609RIjPWOYI7J7ZZ
/rjzY0eVQrvra8PUSG+CNXbR2Tvb2Tn4ucI2Ujd4jRM7CiWBamLkhe+auLQjzKc8
gzd3G//gqewYpoF+IeqmSGqdKlR59iKqKKSDUzv11vZBHuwG8g3irIrcaTXHDSFV
HPEA19UEUZCZbTbbLu7fY96VFfwy1C2DTBBFlhfPWVyO86HI88ZErrSMspVQnx73
rSurk13hMo0Ddlaz0W/nIdCkyxcNVXA2LhW4Oidydq2NGrnznzMDFdslrN5WPOnd
ZFvfmYLrzbi4YyEoVyAF4h3GOMdV1y9zTOOogY12LzZQaqx0+n/1KPwmEgcxIK8B
hHCIRx6wBPrKK/iJ8Bib9HFKQv06HBhLqePC9Uap9yXtBCQSumgRjnyhfdXHxobz
HuhqB4bDpZf9HJRxLXQCtFoZCP3wBnNdYELZdHwAKnbkjm8n93d3J90OMzPEk5l5
tjdFm8NVcjPjOzbixb4ZvJ2jqSKk9mHcIgsV0yfJDGN/PhXtZVlkPJ/IyqWdsu2/
kfX9HkQiF9EWX9djBBq71I1RLGY7MwVqW4/taAzTUzvrNZ4AbcTdkjtE8kg3e+pA
h1G0S6vA/RYj+QPKmGwCyW4d8UyzLXz2I/v5/RXvrZUI1nDYymcLeGFpyhsK22Ex
QsvD7ZqixXJVs04unPcSQ15y+GxF1X8iQlZMGHZPvWtgywML3iwlUyo3NIK0cwEG
rk5hOfAj64BeWdnPaeQq46cyXj7C5EC8DqXkGmIP6z66zHkEgqN8qqd2UJYJhYD+
T7PmfKDtLBDHmmSFDM7rW7qBUNXmZVy4vWBbQyT4I5Y2Nkwts2MMg96R5Bg7uRRZ
t8PkJMtV7bD9gfEqEr+rm1q7+n87K+qvNFEJLFekF6gaHuloiHPva4wxpAFF/5R1
d3bH7k2/KtqGAGeLQcwg3QX71iUgykridYuhTvcFk+fRMMmVVinGFuZtAx3EXIz3
PzK8erasUZqv+IRDcT16kaUDC1fj2cv2YbqmYJu1ego/ADLOi2qqyDNEHkbWUpd6
1TY90KpxKXbcFd0Xo2LZ77h+oLamjNqjpX8lQJunaBggWpZzSrnEfyP+btFTMFHL
IGQkDhb2YK+a3Rjf0f/l5oKENlEbECFNG5WB27SV83xp1kKI+NxvTuWzQIyD1hwc
WxH1UJhjdsjZ0m1aPl/UHlk9FGGJLFHo/EkKuOTii2O9yiEp9osUZSTzzqTkLmUi
2TIETq7a1G2nrDfQDaZj5PR6w7KPXa3hRwVxWaSyu+0bC37O0zR/vH6ADZCTvg0f
HDu8ePGV3Xh1EMg/fFjxcqHNnW2fzUCGJ3LLPef7LX3eRCUu/oZ7DJUcg8QWU31L
EAfQ2nca6tgjRWKgjgcyCFUANbSLB9RyuJqCfIKi1snwbpLyDAJrnLGwKtzEga0R
F33gOkYNa8j6gDT4ByBxF0F1OYQNkQla9L6pZtD2hgbNcYMOIxpcf9NfjHZEpTUH
vVW4Oqf/ox/ksIMG6pU5yoEJODJh0syuPQYLJcZBKDq4xVG2z0cmHabGeM7b3dwl
ea1Bx8rNeA/UJOpcoWwKtSwOFLovVqwSoZD6eLvLXRUWg/V+3OPNfFGxLwoHGt8i
1WVRq0Z4rSvFDDUKjqP8j0b9tArWj68nZyWOp9jYHx9oujgxVqq8XxuR4CcSGeUO
44O+y68uv0hxJps5JO3C3neY4C0g0F6S2smzWNe6OssPu4LHemjXmAePowB1P0xs
sI2m9X6YQTVGqFioGdxqNNeSUaxaVJ2Wx6ZaA6jiexNzjv8A6FsCx9KeKOeN5a0h
nEjA4JjxTwxlpCsyt0nboGnD0ZTvpRQU/OBgwLqg04G2dKtngL4ikiN6eKfEyX+K
7BDkq0wOg90j//cI8Bcs/XN3UV0nqnRsEML2oUFYYo6x1v1Eb2Ijk/lxCaPjQjh1
JznfPIXVlYfY3x/GlbxfLlY4WI948O8vrR3pL0+Ts8xfDszmgjiv9zbeOd3ai1mw
8HsnUQYxi7daGS5SfRbYlTiQEGazWDXOhAA1txclc3wm4Q7aWkoTZ9Ps9PX3/dtB
T42KgVbw8R+Uf/tPqV4dwwBStcQAFhz/xd7X3GLEgTMrC32/lzwYJ/YbIPw8s/4T
k2z7hS6U4rLoVRkrXj7OW0CjB1xwNtRdXNmeyabGXniJNfHD540fgnd6gus+7IYU
9o3akfHeRiryr1gdw9fxFvw1kSPGU+mhUTrpfpmDl21UKOR9w8bOood+OK1Fro2m
ZQ8eI1mqMoxJmTXAstcie/S/dn3zYCWmaMhHcYtfhL8TvKt/2Bh1K7jzvnuJ0ODz
OAgp9PJZBx7Xv2WCM1Cakn+QOvrib2hvJd1C39DoNWdQlm2XW2WelKNg6pfFPLRm
WxFvBtMEdy1fDYGiSNz9P2tmjoFXLp1ldMZOvuGas4I9ryONb5aVBgXStGLRL828
UTnqnrOJbkBXzKMBNMZLXBOuSyprtYnuXa0MieVvLLhLn5l3SXQ6fLrCYOtG/n+t
QFz+hJyitocw6iuDXOrOxvfFNUZBU3lF+SlAcYNWRoTOh2wqBXcXTkl0V9Dt/bt3
GyDe2fvg9jgtZtic9/ZZ8TWvuJ64R7/YFVgWx2052pjVmPn890LStryt8KEnVayk
MryPCRUDaPJSuHMam3rGwSuveHe0g3UOiAKCd9dW0bBv4CRjOLNQM72ARYCa85c+
eA8Eh0+oiZHEISVl5jkqijK89drXuiAKBOvktapRS+ndAJy+xn480PdRAVvC7w1A
mza4wvRNbNrFqPa2KBHNjEbaFR3We1yIdDj3Bj5/sxz66vw1RfLiYhQnSbV4f5KC
rvRDMsczbnK/acfZiBkaQZZCuqLE2Q4XCANw7T2ZJY/SuTmjz0lXzR/fK+JTE4Qe
G/qE3/NKp1DXOYoXYsQ/rU4HeGnuysU0MhDjSnwzVxdA7Qd3p2VrC70Cknc49zTV
wSBzJzqHRZ19vCNU5wUCtBjXVIpMIw3z04hDNutdnxlBkF5wfmUuH4/9CKJVP6TH
/nOc4OSl1psysm2YRf/HzDVEoH/dn+syoaXsCO7N0osopSXZdvc3gl3HWIJfqjaf
MZgiokjO8GqDkU+xY3TIrO1CmRkzQyElzC11prn8SaPXFufCuJrfDJEBvB1iejzL
hB/cDsf0R0xv6CEt+E9cz+EwHXhwrMW1SZv+Pc02n9337iNxEFQVDnvlxEkUAQjL
EmJHQW3eXtHIOD9Mlj9YoYkDlS+CcZZx7qSwkKN1mV2uWc/mTscA+DvwyC+HYEn4
9HRF07z8Xaahze2xTyCP5Zy7qYTX4/TjRv7s6MWcRHtaJBuuVRKBK7iEj1HU5rYr
QKGASAL0qjghez5JvF7KoIgAByFqmzxu3nU9HIW6jHzDXo69P07vfcs43B5HGZ7i
tNiJ5KMjp9aQ9rlotrE2Uh9ZObsFVgkCEtREOay3iLUr9K9/CBx9FTBOZiyWaM2v
qZHbRmx0v0fVuXAWp9/Grc98ehDC3d6+jcxC3DKWmHvc5R+afnJLDNdFpFGvnALo
dOfmQChzHTcRQRPl/33SuB1R0s0tCsjAKJwvdfXYvD7mCkkLavA/TpNu8roYY0dH
IoUGWj1jvFETrTcU1ZGxjI0AnWqZOWzBLTt5lKyQ8rsA8830NFW3kb/0Tsx+fxYx
pqP2T3YOf/vMOHkRnfrMVatBUUB6AF6dzaozXHG+PGO4HRrj0pRtmiS/fosgCeKQ
R5+jT/rjN87z39CrDGcefYqatuGMQVp5mlWuuF7PQCzx36ZGTgNfaYniBnHWqM4t
4e9fLoA/kbPCmFz7/Bx7wmJjsopq5t2ml3VFqCwntp0vqHEJVDCGnWemNWFGXsti
SXRW57gWfOzV1GdfnVIiuKHcGUEfEcZ9Aa29RZiXWiiXyqH77dJTuG7hW7WIfpzk
kasHhaWVXzD2XnHlkr/a+10Ujo6CwNcC4BOX1E+5KEwxVTZYaFMAYojxMS88hmXn
w0Z5iRHYbV1kRORCDcOXPKkEl4vlDflpHs8NH7wxdUcTOMdvBKN7A4sJWi+60r7X
uNekwNyUXnNiWmaKk5yNHP45SryXpsnsr9B+LUS/OtaWcSGSGILbzJW/m+MQS55W
/g0FFdMLOZAZAvhi2sa4qLAicXmw1gpxWTjODmG1k+3C630FjMC3ZdkmfRjIAz/V
RJ3zdI3YFvhcky5Yo+xq+oeZcto5eQ5IQOXWd3Q+lqZKaOtmcOToilwheaqkciu8
qSx9cHytVFDuMmdO/HgGp7DmeepMmPrTU2iO93J9t6QVf7ukb//9b3cqooD24QXR
xKeGrKexsDePCGcu7Xd6EWOvWdg8CaGszJJncnnDpbao3lQZxmmfidSTtSzK3xrn
LZ6WLohEBh2z0eZMd3V51mgyS/SKg25d3bUO4/hKuKC+xZ7Dhp9cTbqesxQqnyKY
8pvjVw4csUozfmtvesFOVZTMlUCML7rgHThT7jtVs3AI1nuGjEFBgCAOn1dNXanK
8aGk3rRitCZAfahnwIE9eobih0EJZC9aMtSvaxrPr8OEjG/LyQsAPfVwLERRFih0
8mvQ/yYOwAfFFjGgqi3s58TB1AHrc12GREUpj3tQbsYr+EinVdjZD6R7KlpwWl9P
7F5zr57WdoNYON9rqUpqv6VlsKgTtkat5ffUshlBezp6Y91jq+RRiF56eos/UGES
uERfAFgSPJ6tIi3fKhDFs88t5KrO2vQ91vZgLfQubI1bUsaVnMrb46XvQ6WKNAXE
4CirebfEZqkQueRSzqUA7BYmgjUHDA7CkR9bZb4QxPa0exoKk3R9hnLuacco8Rtl
rLAp5Zm3rfx8I81hVzL9g4nqwwmKbbiF7QT5MnPoMZCHznS2Wx4Fvmar07zWnPld
E4gkt927OHPZT/dO3CVt6HIiHXfaE4Nad6j4SVJsPKi+JW7EJaUI+VXRDb694ITp
Z6XakY6Kq6YrMzZZV3aBcOpaiorP+45Y6egbBki7Dfct8X8P/SkpTDJCTsxsmiUH
o/o6b3eI+YcS0tCV2VF6C2XvHyScEMaO/6E4HGE++mL6A1GhpJLyJu0v1eI9qSfD
JtvcGHuvp2vzt2h5dz0vKLsEkiPKkqr78kdGWlMZH9iXab8ZD1pn/+XwlknSHqM7
k/A5jYgVBqle9uJ+G8N7kIhHEL+iXfF9ofVW5QcK0tFLzZmRb4yCk+23sepxN3mI
fUNqHFbXgOr3FWe5CKH/g5xySs3HH/OBWthMK/hZBegAFAADGOjY/vY8PL7HquSc
vMLZ2ThaooPyTalkH4Fvm8TylIaGhd3O0meWWO9wBZErDnEC/zQELQQZEWE322D1
lF/a8CTfCEv3eZgPo4O/olMPM2mINBl0W+KscSXo5944QsN+HpvkDtR9YN9653ZH
2nD3g/vL28ohjsnESAVwXPeIgYwsAAw3WPycEdL0wPA2m+LZTgxRG1sr+zMusq18
BJ6p+5F/rTdrQ3IX4VaQUxTXvAG6hw1SsKBWalxJLxmbzBu53Y+Oy3FjBqQ1BPaF
g41BQwm2WxwUdA9Ywr/vqMb3kE1QIXi7l5UWuVxlq5GoDyTNl4FahiWsZXC91TaO
CUcgnM/Wm2OseMW1vdDLJ5IYZ0Mk0Lg03V0qG2giH3Al5qmYc8HUIDuvTtYEsh2N
yGDSLaR8oLGrvBcJRET8pyKOk+ABbrS5d8fDjPmYeA/ZcRuepQSHWyoTbwE3n8sH
sr7lmlbNa3vdEw2xhOdkI0Ln7EL/rZmlsvhAmJObw+8a8AjUZC6iFEaoWQKI5nXO
FBxn6ZeARvLPMUccwhVwWX0hijaVaUwj49s4Gm4jSgmSvLREm45InAmz8cBCYPbA
HYvSXlnX7JVAZHoHhthD2S7YweNDXeR4pDb8p8DFWLecf1quPh0/+Kcn3XOoisOB
AzqCRV6kcAzfi9DrIqRQUaTEAH7VYhl2JlQ3TdW/3OMi/57DxOmqAXQmWhxSdb8i
8cUsU1gHyYC3twJyR193ocMZeCdRT5/D9IM0H1UmKUwhRBy4dgeBzCnl9W/iq6+n
rguioiuaU3qgC3Vq/16zfkaR9IpRFFEaGdaRGW6wxAe4S0eM3c6ciRrJ0/myb8O1
BeloX8weivZSxtHrpFPUvvczqROV3kp+sNDc09ll58VqHSxmuQ2ldfWVp4X6aE3k
ioPidtaQhxp/VWU1IuKbyXJuP6HGeRzJZ2moSHFV6ho2KUFs8WeVXOCAF3W4lyta
OWPAXE6JMtSty/WwmOO319j39FXAmQXgd+zpCP7VYhUrmtawynySqpznzi1JZFMz
AV6v6C32Xn9IVBaXLMH2EaDWhgjWfXJm9Pe/dePQ/Az9fePWJE1meyDrDlA2DsNZ
RjRM0LqBuv++1HeEk0IZHN+gJoFmpzdNhF6IXbqNhhAXTxUL6FsFxdvSqjUxSY7g
xlaiSZFuurNIvJuJfbf4y0WA27VqgDx4++nCNYRr2lnDOrknpH7fiG6uG4eFjTst
7jSg5FlSGqm4LSTJB0c8/HpvNGbUKZMRZYjzsrwXB3en4yKumIKgAOHK+68sHUDA
In7lbg4re+y3mJUSqH89KneXIqPpesra94JPHC8nfMLjOuOrBsPS8CZbm9fi2qHA
EhnyDuI54ItoP+qUpkstM7eyUeLbYVqtflDUAOJT0KtmuZG34gc8+am3xsrTmihG
Px+xrXIWVzhquZZYeSeYc2bTOJ1je/kt6Mk1c2GyRNmo+kiJVkunGjxV6AKu6uYL
dJsAyfeTo8MZkacCiWo0cqxDE3wREm3v4SMeSddmm0RoUwHzy+M/ixskijtfMqab
Y9DJKe1xSUl5hOUifuQVR69RPz77QT6b2hC4UxvdrYoCE0zXOQiYe8EvgvA9+LgX
BpG/xcZZawcV2cTBQT6b50IJ/wpiVJSF8yMCMyW9Z6j7iKzU3bEMeduDJBbBRQpi
6CtFZSR/p6XAcadTvJyQApVYSisTv9jLMaHDWlFUtvxcREPvQL/wF8swj6GuL71o
lZcRtXhj/w/gP4i9wo+GuuC9K5D+C89D+9MgZTBIgXKWBOmsrbURcv2xy4oMFgZU
fMb/EwlFD/MhioFzTSS162qcnpcS7ylkZ+Sw6ryE3LZpBDWzT7kn0qdLgTEqoqL2
Lu4afWE0BGvbXzadyAgKRHtARduxKx5p22T6Cat3ry3Dwf9Q2vZZEn/zutAjwv6A
HLKEzf6NUh7pqZi5JMAFnWzAc/QgsdzJqbEqJIPuxPimEHeVBvPOUGC42UN8okwq
8yUFtwRCXWohy28P3uhXc+zDjX5azL2VXSsLM+cg6nN5cxTsSHJG2kaadmb96zAz
AGydVyB6iXSFjwE4r/ohfpEkteyee8ZovwBSdROAvppdJ9NiOcwJclwcvNXIYKTv
dfgh9Pl6CVbt9b4oi3Uq4GRdwS+EGrEfL4MOHYIrO2Ho6RW26H/0E7ugUpBLEqNI
Xk8vGn31lmqOL7Zo06zEX8gI7bUyedRP8SwhUy+rV6LHkvT+7Cpr2vkn11yHjXPT
zNISIr0AhArAL/SiIFmnCvZWlXw1qx91P6rxDWjAOZ8rfcP458JoNRHbRtjOiec2
rV2FoI2sT8LbjUnHdns1tWWl2aXcs/LOLX2fhdw5HTqrqUr3NCccTH45/gF/fTBP
PV+7axdLx74yJcaCi7XCdkZ7qfmVL1rr5h4NWkLS4CZg23lHe0zdfvcRl11hh9yG
pgwGw92sd46Cb/qpEqGIuarhK/gwZT/h4inK9pMp1xsqTDxVKtV7cr83HQETw3dY
XZ1aW5fhbmOsQdfVb5IEUiIOdoZL327UaBdsCkVb8CtSrx1XiOORKCA8NnpR1c8m
p17sZnQkmP210XNfDrRHeVDeZsOQKGgPiq1TQ8X766MDG1jaT6Xvc4oBa2yVvPHp
pV8XYNuPZmk4XY85t3BlD4EIYINe7t31WpiYgQNzu94t3DIRr8v6OfOx8NGHxcvO
gq5dklPOmAk8wknz0l0i/ArHBZ8BbX+0JBUeRhz/oWOpGfGm9VRJaxRTefizTKos
/91CmjMEUHMJKbO73nGsrI2GxmeagaPFSmNS7Kd+yJTrxRg1iF9FCEgZIJRgvheu
jltGPQNbl/ArtmJBppZFVsqhUjbNC6IwcJn7FVxB1l9War4OtLJmF5aNGTP4dXry
sSiGl7Zhhu3F1cOBz5RAHnm5ZSg/3rRdbPsvHkxiaEnCFZ2ea+nFGJjtQ8Y8yDSU
faHGese4nqV0EbXfrUDKj0IH8TL6K0L7Y/p6fsTv/+zRYNgbw7a1upUhGgWdmwaP
ZRezRmLBE8RSNjfZDWVmkDhg6yWNP8AGgRgOY+Q+SQp/6OL4hnSFnFBEmhq5zvNF
UuOKuKaq5X/XJaPi1DyxiPSyG2gKEWiMwlfzU5S2a6pAQo4oC5jwe2y64jovjK30
81bhXGz7J1ZNE90CesXpVphveTtI4rLqrZxDxlbbcput8QagCPhx5CCxd+R1YrFw
8UeHgJY6jxxVkei6K2ZC1L+KMX2LLO56B5FeBx6n45Me1C9bPsl+sEYFAitrVm4B
Rmv6GOjtVOfQ2ZX+wQGi3/y3cAcE0rrSA6jU+YNf3x7/t7qsseVh6ODfp4duC1pp
e8Eo277kKJoFfKziW4/tk5O6b1q9kKLI9SX4q6f8tuXK78sQ0epebaqP+v64uAvv
0aJ2c8ZIk5flYrAGrd4d14/ONfh5EKdvckUH7bIp/qJlLHbTvbJqYo7w4B8J8qDF
eV+qIkRPJnEr7N4LEn/NBJbKj0wm/jABqaGEHZMGhPrZUqjrMGz//E5PXl409ZCR
tCrfiLTqLf8NfOTnD1u05hcrB+1qpzBp5hghOam44kiQhdlfPqwMQjS8htOu4oT7
IA8tBbkkI5p/Hl41fKojAYUKI/RpbzSRyQJ7mXvYz8XRmUXUrXglEdDDi1ELg4cz
KGWJfcH1AH2kG0VzIrgGpkrgTbCLRSXRTnnYKIHHRp6zkNi9ntAa+1uxnWLeo9Kz
aiC2r07eNUXHXD/25PjnU4Dg5XrHU3GzeGjiWN99X4Qu0M5DQ5w46CG3vOsOi091
Lt/Jyb2keEOkXtM0Ks3UZkttfv0ztORz2S9wzyAukub7T34ZscDZ+/ywPWHW7Al2
osEk0t+vb1UjNQKEjShpMpQ9fgZEezeoFoXuH1IH+h1WzYTWfHsc1876HvhsMaLe
lTw30sUC5WFF5OTYIYPfq/7AHpjwlzCzPUV800yp4Jn3YMKD4DCnEodeyfmIm5Ie
suujEaBim89D4XdGWu/WTG+aMPhj13GEW3n5iMo9nJwzSgHCVZJ7/q8y/o4yAHz/
uOAsDqDh/EeZzCKCfba5P2DiATnSuPTBk0X/9WDDrpQhruYTM0wAfsY3zGWQBrNQ
qdhFBkRDdYtN2drRvVk1nOLBB6L8U4Ms+MMMJm+c2T7ysskZ1taWd1xO5AF0YjIo
WhOjQI+slqKSBezWZlrLTaPVqrj9tC7PWt6QnQLFcSWwmWMlckIwEWZCbXohQ8vj
9HQ8bkdY2NK5SOFmklLFEIBd/9wwwwH7uql+x3NlmLPWgRGSbCr6Gexvgh/IPwK+
FZAh8GVtFCsNPHdpJS6cu9oRhI4ZsE48N11wsWH4Q/gNBiJWwPMJOGXnIXSUgqS7
p5XZTXVN+nHaQR168DURfv97+h/i9L6gilxTwL5LjpDlRN5dGrEdsx5gKn6cHQlO
fzbdt9FySy+ry4YhOmR0z0BChJ+z0G9Zb33OZqtt3HUlqIIAk1pID+jvA+l6SR4b
j4wBE2cHviD5Qxs5BJKJYTYgQbymg28fM49CygHNY4dVfuN8RENxjZWXlOAFGV/r
42pGN9vqYVIVkK6GqaO7s6gqeCj349o9RABs9QE1zsK4u0rk0qYfi9HbSiaRQ4nv
J1yvuyxqs53KZ1L7xoZ7cGjeRG9YWMfpbff7h4qFzFEAA69QXZZy3NDXcgLeij5w
08LB1Xsh0nhNgbtUhqDCemh+fwYIHyUOrd2lihWLQopdWhJamPVYdKUYyCP7Imbi
qh+7+K5SYoVgViYBcC1+HdS+P8ca2jpeH0qbq3iYowzDV/HhLW0t+JGE6c0ZV/gq
+woD6U8aaeM12iPZ1I58zhdrNkQzvw5ULrkgIQsYsVu1xpHqmTEmBYKD6zOcplqo
MSvf6TI119WQSY7v06LUl+Hxol1tkzosM02LMjlFruycKGR/G8Iag75yAhHH6F7I
ZoJg34cngiXZkkvbBHrYXIT8pnqR9UFBt+0rI14O0MWwjo0fQPOaGosjxy0b2r20
4VK06nUPabNj866NMWM4AB6fyJ8ukF8J8Cms+xNl6xkpsMa24m2TE4/djcyleu5C
Ez2TT41AYWcJDqcN5RZn9F9i0UDcdVh/Mfpmq5l/SFoNAluN+7fMXCFvA7yG050c
NhGii1nOk5hpv07hmmymvUWHGBXaWOUg8fj9iCLtPyvkDJs8f6b2i47r19Isx2ar
CFmkCVxc3xrqu3RpaHPwICgmwak855ZDKjP7c79YqGR8Ny1TdV7Nds5khDSnN0aM
ATsukekDTABQI4L+Rj24YQ3BZBlhO1vGjlFvBdDMoUknyiuz7UV1o/RJeZHx7Mb1
ISl9Bq+GOeoU7rj3w2C2p5BvspBmsjSjUPck8LbhPmB16YKu/JiRDB7tLCQ9Eke0
yDMW7STptLwT7pKg5oqFQexDnZ88Uyu6Qv/JTWlNFPTXQ7it4nhNRHvoph1Qaxap
slG0ci8wJhdMi28BvEWc9IwJXH4/9U24IRSKPZkPakyUz0KB4DE3pi7yFiABO0mg
Irl2fiUu/wFMSL1UzeUhtvGzJmDhjCYz++bmzyFTlsBNvpGSZhVy5cw8IzgbswRq
Dy3Hf2gtQvo6fpxfYmBI68VAOriPNi/8JEeF/iUwxIZwzAw9w5BW9KHOF8lmLdkc
wBwaxBcQnZU4ztOSC7fyOWgrCBmHCfO6Mv9Nz1mIE19lT8hhtUkOB+vBoZxWKbvQ
loR4IbVA5dnAP2pgaArLcv92mrnIDOSm+rWkXCf0hxBppRnMA3IzZfA8WFemluQ2
foKvxddrF86QEVyjuJxViZs07cSJLzBDREmIThUL7ycbPtmDTIna6fnkbpPTa9uC
oqdpPujDp/krr1N9sduU8DcRIASlZg8VT3sBvQgNL1eI4pOgRztO5kcnhT1+90T1
aTjLkiSBGC/g266d8vnNEY47DWQ0XVG5vwfKTyLRs8EdtQScxSInph/xtMeg3AjY
SrBuUQrLa/y7fV6mRBp6s/zdHg/9tE1TAaxHtcQLMncDqeU5rqTAvZzOxRiWNnE1
0HGo5M9SottTCoHeUTxZjv38aqCxK3QRFEqnWHqGh+sk2dVp0dTlYVc1SZM3ADoa
pk8C4ikqCH7KesftS8Xl5F57YSlbzsc1vVDBnyejFMekX69t9zik3L/0/TThJYGV
z2qlO04t1gjPoICRICyLHtQIRHAT/QE4lxAhonnz0r6vO5ofdE89dUkl63sZSA2h
oTtcxCiSwePAQ5RA/X63aO6hK505j4Z26AQdxlORieZlhxazCeNljTgA30T90DDA
gWmDZpSxnqTBxhYE7RaWvUY2NDzhwGp78RTsoDQsex5C6rODjnXzeOEipL9bcW55
oiEC1GfpnYSQt1wDIJJzR/l2pw5TOMe1hgRFMi10XIOBW8nEm9UDJ4LikHbCtVK1
FUYW8AmQLgeOGbZc1zLJ9qA4xpYfVyzxaTg8mlt/bNs+xT30tT+kbgIpznuAV3sG
2cmlO/TbNBaTgiqJJAA7va+NporUERybXFWKnaqmA/sabL1oIjN0u1DMzHIJDrr9
c0HNjqPPvtPeEpqN9L7xjizVGfZmTq1UNyLM88qByFibzM10SrYca0idpEWx1B2G
B3AkZtO1sIrVOqs2g8w4TzvgPRzBc52SWrFdwqiIpU6XJpQyncOxUuPL14asv8bs
cR+7om3rEnSIt9Eq7p5iID37IbXaUogQQ0e0DQKwmOTxYdkkSkCBP2xetpIuZZdl
jN9CQEbgKmTXE8BHMA6InkxvCgX/msxKyN8hzd9x5sfhNPaWdS9wnjDt/xSTW6GG
LhDblqTPk74lQKkPmeqJeiCvm9z9YANRzzGCJyWIHUS+G5NFlfl7J/98NQEWpBs4
7Rp86EyjozzUmfUzfMYbBNjZvlhCmkNh+kmRLuF/Tz2jzGyiYSRD0jTsGig29V22
XkO+ddLDISQ0g+C+R/ghrMXi+j3Eo/eyLQ9lPG+vnRvuaJVPStQfTbiO81zyW5mR
mNjIIFTW3OA3W1G28+n8NBGI8A5mgvfXGg9Y9UWKZmsEKPIbu8LUbnFroK/Opf4d
fK2hKJCPEXxd0+HzsjXKs+zyKaU76TiholKUzooE3k5e/tGeZ0IA0EmXT7Ash21X
xtooWYEwvkh/PMMoXaj6L2pBcP/vb9mJKPtCrXJmJZK6I3eRPvCRMhFVo6jTZnEh
AXZBO2qgwOlNEVFcHCSjsJUG4BIuR/nho9Y5s9/RxdjxMjyaRLAG8fpvvqImt/RI
DJge73IEXTfqWLf3PWlXnEC2rsRmXSj4OBC7xXtZHcrTE8xiJufkSaW+z2BLcfvN
vNKGo9GhlBdC+x1OK/Wuz8gLZ4flPf3g0VJWODbS87bGqVC1cN47INpG6HfNrVA+
M6p9XrfmJmmpBWrQlQK+0O4Fgh1hJQ1xtrwiN54tWOzHqiHe2Rk6MdyqNZiSzJC7
iaE0fR1WfhZxaidfMzDD+k2vYMLsmFfNT8q2mro8AXQUbShI5IsZfekDFeBIV6Q1
hg64YArXUVRcQ5773lISYNdRM3rqlHJ+zyk3ZhHFrIwYVC8oW9x9EWXSOAI6Y1Zo
YlFARcUGPzZH4NXrlSPZQ6yWqjcbiM8ciHu2Z9qWNnWO4QTRKDHSTJUDkx3kGkYU
xZbkEpLQNC99MJ2N62vOYMddV5cTfGry3ZEs4pyID1gLpzWYlVYAMV5VSUi2fV3T
qNJ3ePt/8Fx1Ps/O/qesvTdVlUl0dPYdOg74TrkAymNdt///9hgBOczVnx29f7hy
yFr5KI7cJPJd0p6DYDZdd6UWEJH6u0hucycfVBa8OrqgLEZb7C+3w5nE1SXBJ2pr
DuItdF8jlvodYFy7sy2+tG8a0sjZ3DjnvoqA351iH/SBW4nnZnt5y39UgzKhu7sa
T122oHl5x5AV/bC6lBDlzizC7jHma2FUtwkkNKQB5vKbw8KjYCJzaJdhppeZEUIo
QwMO9sQCzz0K7nCDLJjMIjmT9P7IXjGZXY2yrZqC7qafUTqmoBUwNTSZUpQ+ppxi
405zH3EU2VHsrh7FWwEsuckan1xyi9LO0NkUvU/uQBGizteinZwDOEmesLH7DO+M
SOO5XAoTu0e45OVXD5ARW9xg24CEPzwtWONQ0ylIhixx3tJsJ0bPerlSWVWLDFZE
PB7OTUy66dV5Wz4UwFnuBty1pS8I8ggWikrkb2rwuDrTYo53Oa1JojNb3Jlkvk7F
dDfUQX2rz/EFTPoZqpQJUVMeaMLcLSjNETxMfhjWoZFnsYTlIyeVShiBvLZnMwgh
dodUOwvu1GgI8Jaw0WqQ+hSdAgUmeC2CT2hoj3IU2y0SZgkD4mQ+lVUXvYfnFlIP
QmSpJFQwu6Njv7E7FajkG0nfuOj6NvAA5iwr/ZNodIs+4qcVPQM56jTbTZVEqdrz
FsKfIf6Eig4R4v8sIrilFVjBJXGuhccVEATEsWlTC/UUXUXC2Zw1lVK4bMF31U41
1fHfXuVpdlHny2eV9X9ONX0GDFUdBOICn7d+KnGGr0tm4A/GovqRoH8i5+7ZGbef
SvDxrW+Em6UOuufrmh/128NkJYJ/3vv+rvIn/Wn1nvfNHe8mk/aQExLEaxgAkW1x
8egjV77FR+k0kaeYOus3TUJveL0fS7ssIY5sN/ecOUtZqwII/0aap7D3viEgn/xR
W1h975SRJMpzyBDvP79xsAl/PCF/hBTu20QaD/oAMnH2aKTuIdwvIH/W7L7yd7Ka
8DnIK6Svs4b8nNFwMjpdBWhsUQcfL4MyKQorhEKElsGHy4zdQyhysMoImiznI+vv
h17ehoC/P7YdoH0V5ZAEGQd14PoE7m6r9vj/MZQ5tu6Yd1ZwnKlOB9JfY7FQwtrT
Q45OrWeyS7rWREC8yHPnY7yICVJocDKeY3Ohd2FDuaGvppyIJwp48G559qCWM0ov
zXH8brWhH5yAplhHA5SGjmDDkN0oRLTZL1+nmcM91B0gCNzKbdj8qSsum/vcuXSR
laBitxNnLz1O8hW1ICXoR0LZJ9M8G4BU8X3P2GFNEjGs7uXtF46joPHaE0d7SirP
Q0LU6DNk9RPu3LYNMQfnNclWevqb13Zkb1SUjTWrKEBMxUBNuUIK18MCl+60dF++
9Z6v/bck9K9kd0ITFE4sVs4a6CrTLsstn9Lcjll7N5/4M2nUMWa7bRxNSJ+e/DBT
e7Vzsk6epLX2hVSfG4dz5OAEekacWUzH/6Eo7jwshErY8Dq/evsAMKx7xRZTU6fP
qPdbWIGOk0lzdpW+3u+B3OLwT1JFrVe5dXTfG64P8XdfehQ5pClN3i7VnXcl0k0p
NqwtoGY5EOrTuexS1bmzcAWk7Tjxqia7cVXNRZ1xMBVMmFTNf8eyMZIZOsMQN3hl
qcfDYJPwfl16rqAIKLpDBXqiAsdAre1c6HOUO3IuhqbrueJfJGMZ23dEsnVjkpQy
I008K9QGMumdC+4FMWJWiie5HPI2V8GsgYJMwOqTMAqiwA5TyaRVF17tMR+cWDpJ
0dB+JeCsyKbK8AMJgMOfNY5bt0O/qyyErxHNN+qfwOzwJqYSkEOrG2udzLWG1sGJ
L5QVVN9MfICRe0qy80VLfgBqckz/MFMIx6McimHcqHc=
`protect end_protected