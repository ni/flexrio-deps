`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvqr1Wt3HGpZB2xHiQ13wU4siyl5kbTMtRk5PYcPSgHq
h0kAJTr1SeKcLUrJKvxAg9t5Z0fBfH+ePxKzmQ4wrfPNPQjIiVzlWheB9QYPJhr3
k9RgVCMX+CxAeURQUYwir+UOFjxYeqcFJvrp8ThuF/tB8rvWkQroCS14QRQ27hc4
GizUlR4OKUTUSitBH5e0O1n84llC/7z+gR6PZfp7+zB3uN5EjLWtUS2uoPRizwNw
Zq5lLs9Ii00EHrrDMw5UvfGs4czN46i0vUaEg0xUKaNhRDEMlJd/C/moRHMQXi58
ciGu87TJIJD02fRiHJUgyVnqBu5lEcfsBp9cfope99z4N3i44z3F3HHsMC9OECSh
jDBNGMrN/uTJBbt5icE+yo5vJoF27/1YFYJ/YLZqs0AnhikW+RCTZMmWxgqPdXeA
k0+zyyQZcg6W3wme4+MSK6moZsT7Fy8rQa7YEcYrRrg9729e+IwQuxmGtniS8LlL
e3jxm6nsWGqAz5fdcvn5G2oUGK+49bwKZ10Ki1DvzR/y+jQbfXko8N4T1m2uHcn5
Nkw05cBknCkHc7LqHFxB4XaFcwEx+aEu29MrcT+MeliMk1T0TDE2jsKhnWAyVMRi
klHhhCqObw4HwKTbBNqSKL66soF6QNhTb1D6SIp7TjdFd1ZxdzWDNTR5To0i6v2p
sxD2C8E6VxrZ0u9S45h8iv/rLbs0e4pVtk9p+E+shXlfOWUSOlfKpyKagF0P0+k0
xd6zPziW0FFpk6KzUPeR75crT/b52RKUML93OxsAMN6lKnFuWJfJomKejwFop0QW
XHVsqAyG97bsoHIZuJEMYCcxYrLtduZQv9JZypuaBMevIszDttyv78RKjLl8w8nB
1s2ARQoXmYP37non//Elkd/jV6VIExwHGumkHO83lTezeRMzH4B7rPfcFyQkVInG
5bSvv9xoiY4Jxj9LjzywZnFkSIuyCrB2c/dxH+zX84dyBDNute32sGTMxG8sOj2V
hQVdbF+8afx83Ld+1mGV+h3hjVJmRdFD2H7wUmncYNRZXWkBPa2WycwalWGXxhk2
XxvSI9b03qgwBacThK/MEBkexdU3/WFDq3sS7Rr9tblXK6rtcWs8U4ys0m24rStl
IyE0hn5hBpGi62n9frtNeJvkMa5eHzAQ4+z0aHbM8uJ8PV3l4ye3gzYJO2cN9+pY
Ut10JwrHzm5qoBWMou0AMoJ9+NbtkakOU+tJv80r9l7ZAfQu0xAk3oIz+1Gg5a2N
r9xKxSnrHxQCIP2k4Xi/5W3HcLKHHD9UZc5ZufjRt/dvc+JdiPbjswy7Mz1/91ZM
n8GFRy4z2AIP4Gwsdbf6jrQK3mBw2AEtz35dF8akHyBRIBh01+q8zZqIYt2zeuCX
XmFO5cKfqhdlacjNCeY534RV5LEwgd5XNt8HxJtVzqDNIjRtZ3HsUTz7pLeHAsVO
r07ITOBBZDZ/YBqkDrVnkPrldUcc6NbFWkE/jBWBcwKbPpsRFml/5gBHXUMEpwX5
cQkhGzsOhH+7HIqx5ixbRkWz5GbB38QGLV4zNIHZg+538g22quJ3kuMZpMTNJ3lf
jXXQwWH8fkj/4vJgDkKxQpsgdCwOTTmVdTdQCcr6hWpFz6V1D7Vdm1S8wZ1EZUXt
hyvySa+tLbDJKQSnDJonsPMkJSsSG8hPr4sRJJH+I/wBmGdM/9yHS54F6Us17zba
rOap8AuxJ3x8jX6iR8S4GP+q8JYv4DJZ66eFkmeqgdbTbL9UqR80UMotD34VbGG6
l+UEcMTnlb+uVIBTDgOS6mChoCHuLO+1vwcVXn0xStM9v8OfR5qlkqanDxuHdMlW
jNiPfq4YzipbHbsbxatXCHj7CE+5SdqVzv2uJv5yC6DLWgZLl1Gs+wYhbBGzfwvT
2aSY26s8RtLBd91jhPR9mFfkBDkOErGSEvaYxE7RI2Mgaw5+q93qma/7aXxMgbRU
tqLuopKn2D2kcBVNZp650ll2REo8p8vVbQ/5AzGTfazQZNRDFtEQx0hIXw5gkJOw
Z1ZXFROQEowO2M/claMfuUNaxqjepqVT3WMoq4QyuCs5Cy6jQDbRWaWmK/QmsPEp
LjheaH6rYd69hV18Jhv+mDePzjgxK9a6bQkQdqQuN9d7ovdE/DG7VRe4/gEyDxNp
j6f++n4w7mIIKnFRQO8HoIIPnbhOmsOilIes6f2Tk4jdJ1mktkXcNn9LqYk9oZ5/
fiGVV4Wyx3mefooE5+5HQdJ5+erx0lfv9gihghonf59QIoLLZoDuQk4uYJIsma4Z
q2/a74rdnU2/zV1h/CngYXU/qvuHfQw87lsFS3Bc3chQzOCvl/oz2n7PmukC7CGg
IP5RcOhSMJJnh+XS7kcxZJtEZg9r55bMS4pseedZEnBeEDXeRKEgfgctATo4IP0l
hL5M6cN9fvZMJr53GK8Qjr48w2PCqHDGCdQ4PtNF4x/3AWaSQAqdUxx096YB8gEM
Aq286XNYhqubCeHgj9740/e94P80fAartnlkyxeY6mkST5VxCWzPQELSm1O/aHtC
M86u2houDToNgFDxMwzzymbAtF+5nzqrcjio0VnoAHRUHtbx1n4MIARp3kipvdyW
oEDfZAZTUxh3c7eHgDt0ZVxOe2m5f9D+1upIWhUMdSCmznM4KoU0lr/eETnw6lJA
zIuGeFVeZyAkYc9b8n2fXmsfLrcvhic55Uvk/fUxC3D7XGfhs0o98CdX+oJW2HME
eRFSeft6XAP/2qVchw2S4nEWFzHVfKuvnRKzzjy9ZPVtPu8JiSScpDKfzF3GXmfR
Kv1LLZ/8XAnX5ly0zvhmbv0uX47Z4j6/xpskEzozJcmRC1YLyVdROhETZOqKklPs
yg3Pvsg1nWyzoDBZ0aHxg/8vmSQ05fuwb19ZH4RhxrTWB9uSA5xrW6cn0wYIuxzm
GO/jaRAfE1+ScAPH6SfCqharpatxu/hqhnSiZhGspemHRes+op8WwcCOdytnYSRq
V9EW/4l/1sf96+oV7CgLZHuzWQBW16cEGkssT90NZNGLLP0RF5gcGWBRTAy/KJw+
cq7jkTzInJQnW5MM4GXzj9zBNXu2v18tB9fsX7JlocTsAiKipx1TJLjbAO71EA47
r9M9r6DoMfzJ5mzx2wD7JZEdktrwb0cEXae+ccgMK1Wj5Qlgu3d69H+mNoEgsQoc
qvUUiNpD7f1nnBIhPZgaR8+U+fuJT7hIhKHrWKUcmTIYXNTJ0POOJxN/d4ulkei2
WPkCGIsWhZec6vuCv4fqvazfe9+E14fwVUFg9t49UVqlMB1fLx93e+zwZbiBFT4A
MeTGYn+mzyHpowGbzUv9xZU6JUhvdi9XGGnDvX6ngG+sOzKdJkpVdX4uSGEUSu1V
pKSRd+rpd5AIfvgdt1jocXwkPuy632EtmE+0AZghLo+IYSbgx6JnVEnFcqyf5GXk
SXvtO4jo0lVTxgjgO8hLy4BwPsVVvrQBMAHzTxrAiLHEdF5hgqAjaHszXRMpaDOS
M1At7iq1dBhuo9kFSTzqlYl6ehH7QKv/ZC/AmsoiMhXc//vFE0U+LuOaeok5Gyt6
xCDlVU3bg3jcPSPmheybHJkjxMZ9y9x4Ymj30rAN4WfJRculS0FbpMPnF2PTxil/
AfR5J+oTBXqWxCh24Z5c4lUdU4Zz4XVcJeqWCytah8ibdXSFAYQ5mkKkJujSt5d3
QyazyXbl4CgSxIZAaVwciJHwGVP1UiLL2ZW4mbStK7TkQyeqm6mWOL3KMQw/t3x3
Ztv0NgN5LJWzOt26zmbNV5tA//0MzMI2H9HXepsguVdjXRwB+J6RJwgmqZfskIV2
+5tg4KGdf83xhbJ5afIxnM6CXm2hY8a+EtO/JrG7isOMIMIP9z6DZBWzu5fD+Ko1
BFyI0WzxTvBViM52ASz6ufffI0sobb7dEQov7FX07Jym1Ct8Dcw9iWZOXGsm7f1c
58WnCTOXNaZPSg+S2bQKdQFwRcdM0Cfn5HpnCZRmVvs6gpwHSS8fvbxSB566hUWH
36n/T7m7D38KDKgvWmEG10TOHRp+SoZGTzXi7vqEzPC16KCoELy6EnFS+8GrKJ0p
UAzv1hcW5NFgc9BJXiaE4Xxmqwvypq4E0zJ0R1MuihxaLFhQKjdcektJVBAuI56l
59XwSnSneYF+6cSeQomf/UlQGq3aEjmRjuUfnPxy8lFASb7qo243HdxAEf41x3Pb
Ca+u6ONzh0DC8+vqQ5lTIZziygMU8XWFS3cAflK7AsgGoWuMwA7MQtCcIovfNlTw
OXohu1PTLgANHTzyDH6PSACFX08Pjvt4N8pOodyy3S0u2PJf8AJgb/q5gCVzZ17S
h4iU8OCcbqSza+5ckaS4vCYUgoLczzKNZggS3saX2YWYkubw9KUuyV43kv1n8uc6
RHHrTmJNxXNGgchGhUHSKvOqAoBZhT3+gBeh5KWFOIR012dXqagAXY0rW2PBnz8k
2N0Fp1KbFZYAbONrWtiYjDXLtrmWzk2ymyW8+It65vmuN6dF6fBknf2Pp4DPlmEk
oB9raEIVxdSYhC+mcwQeWRiJJI/CdntS0kzC0z18MqFOkCJeB5XwmTH9oUOtW1Hz
qo+EpxkaToXPWJcSZeyRQbVhPGGyrVpoye1AmtR1zfH/DHkbd6eghTrpJPWb5O32
ebQKuQKO+zFCCAbpGxSSVqAO6ZuXzJrebLyiXYl1bAl8G07abbSCMp2XGS52Gw6a
HHBvlmRu/PBcnDZY8OvINf3PMldcDPh69U1BRcwx8/zFJh16Oo0ZpSYiOZKBrVOP
plt6BtQOcaBjGpMXG9JVcufuBwwVBPs4V5K8f1w70cNnNzOk/82H0U12PwjuzeK6
UIrzH7OawEcSE2cvXV7K/srAyendAWjcKqiD6DhlX4UO683ZUQ5HLmlf5nmIOMzi
X9sZRXIrxt9qz2l807ClNaOLgf5oFoDLQXW6xzujqdgryY8oMID7NQvIexll09GB
QLXQeg77u3I5+0EjMmYdx1xPhblwsyCL9YkjSHYgCREEb5QQRoqAIIUOBlOdBs/J
ZR6/HSznCyFO0HgBS3pcZLb8GbKdjEa6MnoqKWMDqXHd/v78HWeeV31oU+o8hILf
+aPpoUWJNgm0BrsmgGUpzSzvbNjD08bNr0NhJ6L70U8tFz/4bAxl3fsCIziKQOVD
DTgjKCwwh+38D269nRHQ8hdFtdWmucToJNbG5ZWp0wkHRSO9Oe4suKt/YbCdhuc5
zPVxRtd6zDX0X5uZiNzcD3Abgv+ChCMZP8XXPhnavqLdy1E9idrbVNwEHlYE5Orl
E/VOUsPbjw08mo41w5E7qDTN7b7yqadjm+E6yo37cx/o3LW2IRD1N3z8tvYzZTjj
hOrTj/UB9wk6v0dw4tlBJhKwvPJo9i/EsK8cUXcs0wEOzcp70dwD6eiy33ymKj8T
HtpBVceS0iCFf0a75hbCD0vy8mohbKE4tdJjCDIDMlMi+Z3kt7wmeUyJucfumSgU
yLO3gbv00Yb/riEMYtLijbnyI6YK3Y9kAk5PZ/cXVcsoOD0SxT8We6LvNkx9ZeIl
2bY5n4VL4tVJW/K6Bh1AyI2dZNsrVJiHh0Tn8ZzbBH9D80a32NX0RszDYSmgPx/W
4uIiBQHXbpgdr7F7N4btxEx6JwmwZAA2O8jWsssuMNmG0x+Zh9p5SIXQDcsvKOrn
toE1YOpx1sdoqCLPBG4S0Y9WDK6YKchY6oE4Iv2Y82hrPnaGr2Q9R4Qa7ZQIVEAC
P/1K8GlxueI0OfVD1DJQZekCHL225XSfboo17x/XcIcDHVHaXULtt18KbXcR/1C2
vsVKPZS4OmJVxuStsd1873inhvcUkCq6NXiPu2ak534m4ZOIO9mH95OlTpYENAXm
NVTJyEDe7vYwHQndIRuLU44iK5QbT6EH6D5EN9yyiy7hm1tSkGxB7zFDbYjcy+pd
VZxj6X6VxYYpqXgoCt7XDhzgAcGJ0H3ssaKdu/x0g258Z32nBE+c4Hhkv39BcZ9f
1UZtaiU+32+Vrx4iSQ4lI3wRM2uN93nusTMWxmOcvIucicdyw0Xn4wf3zpLGWdGR
NZ2tOGVx4pyOvYI+09Mq1X0beDIbPwWxBecd/QERr95gYxJUfBORX07FQ8O7wIJH
hNJGrXl5YN5Ijv8iBEAtVWDQw04i5MaR6qok98Xub8smHpmp9EKCRUE25wF0IHYs
RPB7wYtABab6tZrn3UMcl/j2hnEqEv0+RbM3XCZn8NQMtSFfFpmaAPspxJVIHSIK
ufSwYwYIKv+LAYB1FIRdBxVxwUH6YXeere8YH4E8ErwIfhVyfqCWGO7yP9fbEfAP
e+09fu3sehWJIZz8ZbcGLZl0DzXnXbNTAplDZ3f4UFavLJ7DwAYkFuF8CO8pJGDK
stWM/e6V2DL/Yj7ReHYZuLW7PBpdCLM00yxppBA1AEHqh+PTOxuUpDMHGqhICjU9
6LzscYCnyU5nECz1X9VUpu/DF1xHRFxcFOrA/WJcmInHk2gjYovHscgMfGYZidXE
qdjO+QTgw4Lc/Mtlf9oKFxo9/V3yk0T6GlJdOLdLrUkR13QYaBRXi4ZH0j/rwyhC
Obh8OnyifT1PXG9as6dBF0aLFhoepJTwnYOboHBmV6e8FY8Duacj24Xn2SyGUOw+
W2REi0hIUHN/ScX6HjcGnA+hN8tMjQXCXkEKscSwUeA7ogYkxKLF5i0bAOtroKZ1
EqxNxCUEuQKh+PRqxLNXHBjvd/qSjGHj6JBbiQaPnvb9ftt8qgF9+sFO6TaFK6xC
/Se6TxzRxIotN58rCTd/BB/ua0jjhBbNrqXHony7wDINSl5yBy0V5II6pRYJoM26
umY9T1ySK3M4+p0rF2vOn8Lc9NTyODC61CrDGtvD2Ld1aciVZeGeDX0M62vu8tx6
t07uzeCPUD/QQ1zVysBgu/pQkCRPZ83ZuxiU22KnoSDcrcute4Xh/1vglyg68lBW
vlkK4Jgbdnxl428xDmo9ovnMiPribwkk7lo3Iz9hPw+HhFkTzKOL6zSNdSFyMFQv
4Mg6Ild5P/GK8Jj/IOWQFlVbGAS9JsiOuTjvR+rjgvgeY9ZIj5GmCs8rT66Stg3F
3xcxwZkuvcmsDWPEB6qkbX86y7nJQXED7U+1ztPZORuXgiMRs1s+ZStneWFH3iiG
e/wRBRXYoVqpO5CDP0O5GPTCn79qoi7Dpcm9rgVpVcH5nbFaXtDE/N5QKo+MAvAo
hRcxHLEUXKUuL06Ny9Tnnl10Eq3z3nB+LjxBMGoPqljQY6mv89DE4DlayQ0B5Ghi
oa3PbmfmkFC8KJ3yjlO10I6MF5kaw28N1GGLe6iYeV04C4OkD0oFw/btGOkIrXIj
P+Y754KuNp2VPFHq99cxtN18qGt2YQbMhe4DIgY/T6VnrHUQoXhwkfCTTRXYtqDN
udgWCcnGgTfoWA/R36fLsl+PeGfRcl1o2xDN+fOd3J6rQyQJXxWSj3A6nLZu8sWQ
acCxEy5idbd6y9ssxY+jwG3DF/DzxGfoBZqbNWBneAdaIDOCOlgFzcISN86xhz+5
12+CFstHUNv2BvZnVr1sginz32SWi4LQQTG8u8UiB+5LCHtaY16RJKwiXabzchq5
PjkgpKGQhHcdjQIFsRokHsfulv1SPomw/0PUi8gP0Im2T4voGWSGow61QnJgntyY
QKU9g4B6rhYgbdEtQHgWvF4THSVMW5tL+CO0YRXiXRhlFRh6Z5mBKVNsHM0tqwWZ
+whaLp4Ygse/7Nf6EOz5Z5cV4YWvVmpwE/YvaXBrrVsLPYyDGcK5ms6j2A1V60nJ
eldOMBSPP8s7rGZPO6po1Yb2cIOQFKUdbPOLQ6ygcVH3MtksELT9DDrVbY/uZx8R
n+ugLhsq0kdWC3DI6SWievnoYWuPFyjeOhyDKwQqIshUsuf26PV5aWg9h24P7ZkO
gdD8ZV/sp+puCnblt4c1P8SOEkdoMXDVxVp8t5nRXgLABg8viEmAYlzxmMqd99hp
mj3Lw59lj62gA0p5JG23ahX2U+Gp3Zws1KeDJ9McFxm4rS4UgAUhKar6WmICC4Fg
UDYxUqqqfp3V2DKg/dmit9h7SIsig1KKtCes+bsjBiT7ZjV3eLV+/0YwwrC0S4Sf
mN/+Ecp9aRYIp0J06ZuXkZKsxTLXe/HznI15DNN8ujgzSiobEE1YSVTF0t6KgKN1
0GiujSunb76qK9tUgXmwyY4ksgy6FgMvdRcY05Hjg0crHr4xbPF14f25Ba2i2aPA
/cJG/FrH/MfG2BJqOeGjG7EULsnL18z01gOCIkxIHrOI9kFd7Oq6zZsKNNfPyYU4
KqDT47WqyW5i8KkQ+jD9ObKaPkG9+su6i8NJgMWLYp3l1aPaOW149wyJvd6nfu4k
upS9Yt1Jf1HmxF3J+9byPBcb/0oq1Rzm5i7iTFVcrBG/2S3tp4DVOBqdsokOzUdP
ArbBNy2cBXgDfH9CJSrccuUD3uyQ1X54t3c+pmO8JjFUe7/E/OZV8mV/Yg9HMpgY
wS2TCYi8Ok+ZScO59saif1vsu3x4basnAG0rmM49liMfD+M+DE4fh3MNrzYWTmin
ak31gSvEI9Y/tRlwU0hKoN49SKgOs0uLI8DUUZ6rc41XL/ZmVCS+Z1RcUx8YHF4n
zCpue7kKl6DuiN/EJvUNIEg14XBiREuRn7g7n26eOlC5b2DwWMo+fKu1vRtSCbd4
eiGFaRc+8JThIRr54UyrqbVMujG7BBolX4Rqv5YzAKBF6V8loQmcZ1HLQzprlZf4
dMVkUvqjGXo5RoIVvtHg6G0+OaPzEBomLrCkoFJbuejiGe16mK2GN21J81jLa5dS
biPh4s/8SgzEtA6430RNMNJuUQ5TI4/aNKVJcD7+8HrZ2Ffl7HlFUZjQq8IZwh/R
eKiEOByKfOKjwKVhAe5mGCDNQ4rED5NGzSbx3NazukIEqB8aoMEWMTlO/Y282vL9
NoTl85ooi2dbMNyRuCd7I/7I0ztvjRImbcdz0952BOzPK4F2lhwqEAhHnIbUs6jR
dkZ+Y82s+IrQsXwjQlxey2XPEW2P7lQuCzpgBXKLP/0AgHPf50ABWHLIb+dCGDvN
CG0wWuk3SnStdNg/7dX6dRY9MLxC3Bdxn1QtZa4Puabqcd7PTGagXCkf9hLvmrx7
r5nkraqXrxKdaq1mNr5UAB7KFbEnjq37MozCXxs1B38GCQ3BMTA/M+8+7pd9nQiA
MxA4Vm5sn6uwquCBs9ImJ4vT6FTfSjy/hfr8zt8ir0OJ7ufywWE2eOOFTeHrWHis
HjvcFe0A51jkPYTWc0NnE0pDLUP3zpsklabs55w7e1mQpuVUzvX+qnwFcigUlNAb
NSm9UWXlRCnw0HeW38KWdxH1xiQ1kKIV4uGWpS+gP7VdJOnznKAG375P40yxFVpY
9UvrldFPKPSXZrTCVt9Urmewlmfs5+SQg8tu3Q4WVyC4EfnKaq00FwiBlsfawit6
kIDiXXdOk36zrJ9BlOZ0Saw2SRVEQeY/T7B3JJi5FHjqfjDEqTVwLv7N4gRk8U4j
bxNWEB75NOiAxqhNWTX3iRp8kgcIxWtgABiPbGSRAiVGjeIfFmNiZSe7iIc31Yj1
1df41zCFzxoec2+twFDRq8IQyzOcHOiCrQfOPTFboBjDUfUp0Q6d0FlRRp6Nbd0z
cSpiRqBOVsqpSdL6ilAKUkxVl068V3EN4FzKDBVasQ15pwKOWwQmE+uztc3fmxVe
xsnm0xYO+j2uKFuaIusEPzqpNqHUj18B7WNythEYoMkDzuR0iLj15r8uZGT6iGq2
R3RsOnrBxMQpV3SiRHmN9cEY/BJdlBkCGjYOiRZkkTzLRiRwhwSNLCQgKeyN22Uh
9BbXSvFxrcmNFCt9leRK2AH1CIrBCC6I2+vnRvw7qTsCh2aCDX6b/B4/Z/MlE1C6
L7xHqPYSAtM3Cw1e0ol4OvQa0zLKzw6gyvxIjrrDvjNTbQ8TFvKlMNKZxbtm+tNS
d6HbMWUcU9s3yaQG+IKL1Mqc9+BOfC7kfxJU6of7XUWtpMYIysseSxQk8Wf2kqNr
bAhVmrj7fv6LPpkYWeciv7C1KW5Cp8XbZj/4lRlo2PJGCHSynvdjkiCpyY3sB0P5
I1mag8NJ6P5YLKPNqE8M6GvlFmNTx2CVzMn4YTB3E7c9cv4eJ1MP14Yb/J5szohj
TMoL7GsXhbvyWNpPIeoXD0X4jl/hGmr7C/2tgA2+Q9b4X6QR7R7fkbV86Euk8n8H
IfgGnpuyMLqIV88a/9eCF5zh5JpATTDY68lEhV6pfyUdJ5BYXG9QlNclDqrVMpks
BBx/XcrFoEBXvmxG8is5k1SwYX2sFxhJ78UNU0gLa11MxwfO208d2TIbXENNskA2
aYK+0Kx+1RNjaceTqDg8a0jH2pV95eYSqxpHkEKeC8mGoWdJMpPBGRfsYEKkhl3Z
4pWew1eq6/8GvHJkrE6bGwhI996ysbY2S+H4LiyXiQbsiDyradf1Z08QLjA2KRJD
TjHQvN4JvcHmOTQ5hhl+w6Mp3+wt3PeLJp++4TmZyZmzXm/NKz5MLKmf4tIHzEEs
d+wbJXv0+J1isZsKqH6/mF4mFDbP/OIRkEXSGt1iiYwIZZ7k707ojGMBMPH4Q6wF
T1vwUClh1u8J46V5nXIlYjCX3whh8SjDxugyrnmytz2/YB3vQZNZrguHqMsD53ma
56TPk4VZ/PEQgIE30HVrV2K6oKjXTyXx0Ew7rMW8Jp5p/lRYq7f7mZR+8zvqoGW8
omOewQEqy4QfphPYWjyEkIDEe2zMIscKhwRbh7lNVLF2k44dIbZ2V9+e56xzAZPx
RbokzZnA4t/QtrfwN0kYQyjf36FyjtJMSc27mA+VDPUKJbEnQ1M9rhgu+ogU90dE
CeifMOY+zT4W3LZ8jygpPFB6KT1GL5nCH17/Ecp9M3QXS+AodtVC9BccUgRixDpX
+9p/jgLOSlW2t6HE1QYgt2h0AdsjPcQEMEbH51Zp9NLI1fc/5NRJtmTPS/bbjVQx
EZUQe7Gp04LpdqU3mAzZf2xU1e1tRpP88VAh/1PuQo7CW+5+pI3rpkulgm47F6TA
eq0ee8dU5lcaFi6b2MifwXGQ/hcvwzznyJQE4qTrGDK759WDYuslhoEpNGXoi0Ns
9egY0cMAM+BkGJC62QMQq+xGX+7dpDZRXZOy67kqXNwSgXNTsgIB8h1b7Ek/NRK1
L/fHdse6WmrjMlLPAaKVBJpPlqOn1W5atWvBIDT0RZ8AybFUsOMqzqIEiC8kk0st
7FyAkPJOAnGD+IlOJbEyexqWvf9TVJlG1Trg52ZdvahxTK/9yYbqb9UbKw/TU7uj
5/B82CJ1qw6YbpreDljqNYEA0Z3u1+oo1OIAeyK9d3afPIUOJEUEe7Q9jMyIjCQp
P5skNust2EG/xccF6SxRQVHdT4losr0JbpniF3/UzjpOj7WiHPHtHd8rPozw8Hxr
4+BY+W/sT/twmDYca8Z4OgEKK1snLfv6a4ItevP7oDqIQ4Avl4BtHl0bgP/vkock
RS9bOycGtbWF3z/MW9BTlQjJKAFkH8rZbBRHdFkVXQ0Mn+3BqtLWokRbeVLw2WAm
EguL3/2w8zMfuzajCwos5h7eCVstPfSqH3t+z5KSAyzGYb+tvK2ViOofKt3aUhTG
+Fetl81480rVZL/XRb/+/DW8+PMII+zdvtsVZEtgEa2svQteMRFWm46xuqjNo6Pd
PhVUParBRYMjIObLdBiH9yrtBdPS0NRb0cEI3+TufClYGdXrsP+rJZu6idy72iYc
3okz7rwMX0UlccsqNXLGM2dCMfttIm90y7O1DNL1ydST4dVSYlCkjxHCFd17Z1My
FNqxRydzZPFINcdJY6+595VGKWZR53/jhecEua7xmMKyU50kYtaEX3CYDDd8EZus
lfmSu5Ia8lLp188X2disNDvrosh7I54B87qbBfBZ/jZCXVcq+vXtHNdUQ2BxIW1n
Ow9saqJpG3RzuXMf4hHDKRrrvCp1RJ8J8ZGNPEjR5YZLglGhCS3gckxMhqMJ+JqM
z1vl6z038b2f1TQ2LlrhiNKb8mCixWlFetNoJ/0Kh8DTGtpYyrPn1tMarCRhajLR
1a5GTzZ2wFA5ZVyYu2YGS11p3D/BwYd0jFl/XOkAoNj6o7f16nr0KuBn+Q731BwF
H+5wlvwBC0L5ChPFOMkW2yWmuGyw+FpWocd0X5fb3+I1EKsKwPd1KJ+OFadG64XO
MFcmNCiey3PlkQoaTOyAkuUIeHT1zt+faGtib3oCLXaUhcLfPxKLvqATIXUMsdvR
uqScbz0Cq0fzVjKHPZDONL2q41gvMSJ2ua7VGfJQfGRFcxRf4S72OPVtrrNNvJjz
I9LlVG/x5yal/Hys6FVc6hGC8yv0wmCMz9wFo30X2KQIcsNZzu0T/DG1bD+nMUca
DQeFnZ+ACjkq/Fe+Z7wTyHddO8xtM25vc+76+Y6m6QHWExMvDJKT/indHihzN97f
NR+h8hfTNTcBbnYAzrxjeHiqo5s+6WzUae3fWvlf6IoUHrzoBUEh0BWgiXBaYXKn
IC7rOEmAXwfbcdXG2owYny7c04u0UF5psaTgRArshgifUEsxf22S2fp/NUpmTEg2
XDkjBQmfHU1kPpkSwfccUmSQUfQZJA44Mbv3CnS0kawMPbCucP/i6IcVc2xAago+
P+G6q7R50anq6B+8HEVTFSchVKxVPQ4vrPcFWGwtLEPp315viLsvEvphgjImY3hT
a28/4Lj7UQBBjR2sTLQnIssmoOV3Wpc1ESXsGCw/BGwdaxk0SeiokCBeSQkQzdsP
0walYDj+cEqMbtMwyFNAu2V98mVnD6Bm89O0ZnZhmB7g4ZFhSBi0lqxb/gg2qIyb
QtSmN6B75aM2OTakjLYgaLswBHdygmQ4V4Er37iR0Le9MSv16BuWniDGxUUz/wPj
5bPg8Wz/CLtIXayCXRCknAXDR7/Jm76bWgPHtIFPn42Dt5fMPZigOZdyZZPE3xHA
MM1tc7rPBVK+xZSLufJbGWi670ZwmG833z+TX9iU2CDmdbq4AS1S0CWGTBxVI9Pi
IjKcqyVsF1k5VBrtVUNTK9jHM6zx/r7sWCNUwx7QmOgiPR5AkPnG3mlVnJqNImY3
jg7c4SnlVsUeHDI54mvlt3RBV9sDIOEAHqfX7y+5lGdZGqMbnIYoOX3ihBVUKHGU
zHcJWQLEMGRpI78ZHwUSDlFpB/xeNcn7Egd+GHBBOPYpmSGf/0wYKoDtN6Gs8MrT
Jkfp06sBdaVCZJosiEIXIa6SyClB9HgWsrut0Vl59aVFsf6RBLVlBsslsSoVO+dk
5C2SKDyTfW4F65fMgpAHIzQ2gIPXE5torC8gCPL9aWI9tTqo+HJ+GxAvW4yxL93E
6f9wRyfDRa7oiFOqS3e78MczInDx7gX/EOvw7LdahA9sntyLhPRrk9TdrrTRW3as
wJ/naScVV71XK96J2NQ5zMSJAZbG3U0Ar6Zqs0v6Qxm2CRWkPiR2rvLjio3sgprJ
9h3wIVsJS53csrh5GFvygS4243e9dkPt39HHcaNOCgrTg6P1cFDn9+HXpepZwgOU
YEJz1i4OcGmeiV2cPIo/Iy5vr4jbeGfxmlH/JjEvilE32LHxhoBa4GoY0dn2NBUo
7QQ3UVIkuflHb1qCwbaVcNGLlj7lRmJXvfw5P+xNLd6YXVrHYIPQFFVi4xoKR37e
OK7W2yJvP5v4PmA5DHenYy7emGwYoclh1+PkFA0hg66b09JhI8+FAe4p0n25H6r7
9NYSAeDUEsxAmsRhJqBjDGWHLJjRSPwR+oL0cZ1orW4mMIyF1bqxMyKe9S7mHE2l
pGk/MgJzr85q7Fj5uSraU6ZjCE/DsUaDcSmRoxaLvF6CbSxuoEXVnXCXFCPh57oY
ZRoG0NOKUY7qcTdgPzxWrDnyOKmnnjWN8h5K6KjAEch2tVt/nE2fyEgxiycsNuDZ
lPx5CODsNbEawMoqU+TxiLD3DtjrMdok3DncrnPAuT/doj+Y0+8ufnh2r+bn515V
/aR30MhpeYzX8oGxyZqJIwN7su0Gf6v78GY2rl2clhlYajx4avc4lFqJOG5y67/I
ihy++rKPmQ0Euwwx0QxpFZ/D7NE803FFdM0xyHgMSX/1maTMBHS27Rx1PQk0EO7f
1cp7hIV2o7PrPPtq+LA22Kd6c+kMbIOcl61DQTp7I6pra89guxTfu1KbQFQPnnM6
MU8akAHsfgQg7xkow0GecktJ/nDDfws+zQf8QFQODDME5AcnQy6We+kf/fkuAnxg
yZaqYxhmFwVxAOVM85ok+ugLjFQ6dgnPVGFZP3EUW391A5sIruQ4VUI3ekjdxTKl
W8UjkE9madG/8FsPADxc6R3JjmQq2PJFz5uoPBt0DIXqKFCidDYPJRyR/TIg8jtb
Vr4XImOe6zzm/XSPuCgcUCQWyVcWdRb0dcaR4HVb6lEM7fnEKE2ZG47k3jVzGFMD
qzv8ShNvDPuuyeqGmgc8T2s4BcztVDMJhP7sCKKvPQWjQlMOPuElm2AFXQaVgBzU
qttTGC/z38HW9Hug4CP4Os0ftEZXWrSTu0ndL4mhQ9+FJLUWlnD2gOuYxbD0v3p/
WZtySf+MJrG71kQ/wLkAB6GWiydcLEtc6YAUdizeVSpA/D7EpulduUfQ1VN/XVSf
tT3MjvEv1FbAJILSbv+sILlq1woQSGAcjo/5gl0Jh3c/fP0i+ZdS5wusl3zqGHZD
WBBEXItgu8Tixj3+XzAjvWjzAx8Ws0sPrB1HaLbEgcOmaAiMXwUyULYF7lOPpDbm
3F6Iz9ykWT47iQICI29DLLZJQ1MaH3rbIKYsoBRz8H4jpDK96wYfvE4NTyytS4di
FXLAsbxu3KSBUsL6SjHpl+bCrj8PLdQtPFIC83VqcChMKFR8gf6N6rHVEnt0ciPe
juJ1BiJJWfVclQc582FgYqkGD4v/UPGxXukXPNJYJPPaiTxzU/Wn6uLe39uLBiDO
kpL/3CM7B9Z1pnL5K2N87yvfRHoEcdiPxe5Rro53wOENEPLLJy1JHF5ZWt/WwWp+
rUwTT5dAdnOz+0Ivh2ns3d9gLj+9SKaH8lho0wdNoBOzAZ44oNTXy9GBULvCfJBt
B5Hrbdm5Be49puELaXANRXA814X+YNyjgXKF2KK2B0LVPipFDcrXgmAyCxU7PXOm
9ECOPk1Qhv/aJHFFddFTj5xN+HhHupifuBjEiYo1wlWG3felfMor6CEBAHaXJh7b
4MUmD/nvs5WmLqMSdDK4FMzZRX9Y+yNcwz2lcVfmr0QBzRl5dRAR3xcQMAPdjZgm
JGb2CdDgg0FVTN6t2GBaFjHSiGY8owfmtsIT5ga7XpfnRiEJRzp4W+fLkSeyK1ej
0qzR4Z6WwxwiN0ww9+ESbcV73F20ik3rjIHMM62iU132JSxc1LG+v6wHZ5uXAbIG
/HeSxpUMslIHfksVw9mHcA8kuS3MNVouzkFawdovDKPjW9qAB3kSrqbtu0Um5skU
/vxJbEuZM4ZoWJtulclrRIxUgpwVww+DxjBqg9dnEPc7AZv7q1UwEqj1WnsDdl5C
obNJwvtg3HiCngKEOvq2jzSblcr0MzSpytQQZjalC7cFNzBYOr6yA5q1zTp+wJYb
2jG5t5xRdnENdJG8ByB2WFNEqUprGxGnbPb9HWmkLqxdBtWgDsbxMsb+XVfhRotY
0idHXC/dwwmw9SVS0C/UltUAYhbzv6RM3vDQOt/mpkjaK6o0+Tw2ZrPEdzqpeAlk
GnI46UBahxK/TObVRURYVhe0BA5JflemnOhGX5kMNbEMBm+7JsabEGww9mK6t+5y
xs2EtoAAv0FRG+nHDiInn7t/wQNxykGU7pM6rNXXyX9KHqmofM1INGpGTnutquSZ
nOv6OvQw5r628ZdGcF2uDdxnrTQcubHaUUS52vLaUw/zMecx6kxr0Qs9/hNzCabi
toUPGB+8KF1gJKJqIHG0RTmsZ3nDA5S+3i49Nj4sS/O3Fad2+XocpMpY+UwcjVxM
zj07sC74nbIdPRMG9m8rxGsR4wGFwpE28Bg5Zw7Ax2qDuBVa47ZM6iWkQUE+kL2W
bRb5CBhDluEonMZQAvl5yCyvaxOa0xKMspR+pKwjfDcD0UbampaThqiEqBZZ5xP1
q2yjcjtorpedOmQJrVj4vuByXsb9mXpxZrriJBka/+Ysm0Y4SPxUBbfwPvFJDHp1
PAPftNT0dfJxkZ0RO301fptqhwONZmznTmbfjYp4xIuJN7OmJ2mVPEyrekWTtNt1
h+aTunsZffFW1hoBXFtEtC8z7bKc6vPLQ6iv9bLL6FBWA7iJW+MninjRrNndt+7T
l0rBDrOqebuHtnv4RMWXpkufW6bdvW+eWDLga657I7t9EeGlWeIqfzNAEjn1djQM
CCtPzFj3OXjNy5IVsUWJljTPSWQahkK20oYAcjd05sD7wJ4/KQ6+YKgxMa/94oMo
kBjR2GsvRGaSlzYotg0LjuoD7AlwbMwW2NCkSH0Erg72eLAyWFxWAqKY3QNPPBzr
XpYap/309gx4bsM8mJTgDUdmvol2Iyca6uO5t5aafXafg55Ojrr3KW+9DYK7d/zp
80dOs7FzCArhi6BJKnr3OOQvAlHX2+E5qQ4DsmIpCXgKjJf3qOKTfbD6GK5MvL0u
T9wRiHkn4RO5RrfxFTBV6avxwX/ZPfsFtFZF4dRcqT06T7FTJfXOSPvVKECbJ7fC
QWzPjni02HNLmvZ+sfarZ8jdYqoiR0j12Y/2b8LFjY/8y6Vaz0CReZi+NPHIH0L8
Cz2yIA2YEDtWirkRgLe15jNX8y3LmVRvc09BKd5078R8TfE9DsJ6xaUODt1OYMF3
oOZgd6LfTT1jpmzA9t+5p6TDQK1aH0n+PN4b/g72S6wGT5RfnaXzjdHpXaXa+4bO
OA/jTMHblpa/A/OlBf15qN8L4boyh3BehPzaORvibYoT5AgasSUl+z451iyeVk41
8WumDNf5r5UpZm4XgQ81sEBXndPlV4WNFmRPnwOYr2nKeyF3wnw0GSZEMxmB1RZb
7cRrb+ccC0n3GaGE+fb2RGGSAo+nACGt4DJlOsXb9bs2MUZAxM4pFjMsO2LCABHN
7Xv2XLyDMGzYCQ7eb+6mFspIoZYR/MDtXBUFaYvUb4AFtYaRkooT68OxNeJhC10Y
mcEVoAePFlws2bX2s4qSJsb8gLkBvdxAfNJTkCFqo142A9YSDDpu4H/2wyTD2f+j
WnFuwKJUnR90UoV5fr6GacZuTHRyR8rDk/ejL0MIVYndmk0LvpotQ6zm6cs/Rxv9
vKsOgiI/jf7k63qO2EZuFqqcG+ZNzvaHyPeslKo5wiLPsFyZQpA/d5EuvwGyZm6T
i/xvDiT4IryzwpvV00XtDHpiLmiqh/MYm7tTFYt6Lt5Q+fhrJwFmjSk9/qeyrHWv
luR9uZL7WRNdiYkc/N1uqEyQ87oWKJUXEPou2OpGVzjHXSRTJJSdL2cX8HtiM4Vc
uV1RneGYqwf30ygogTjbPyJGPB2CeWNOGJLuonTJHfiGgzQvqG0I8ga19R4kQgeh
5LG8ZJGF59ZNngFZ0pxTY6/cw+oGnheLCh9lhaxqK+2eK5K3oJW7Daup+DVkkxaQ
7GIFoWQ1bfFrURIb9/JmB4bPDHPxw5umWMTIlqovu7ljvKUi8Xv+DTcBMiposQ/y
yY30c+jVXRn7do3e0DkoSTi/Qll9YBrAyO2JgqPzClneoksKAWw3Rs3cJyA1ogIN
QHE5AZ10UiNzaAlBSQ8Q8oo2VG6ZqFQ++z4oxfmyNXvIIdHcV598RqamhZlElKQA
1zl6jRc5NTSvVXKuYHid3+h3obRrETj7BRNzd5ms91IWJ+EGNRneM1TBB+VxqPR4
r4/0YYpKAs2YNDUnv9exVv9pGRuUYhptzMafMmyi6qUCTm+CHwVmcjzqjhLp5bBg
PQzC8dA0Zy1XTUU8ohAGesYX3tS4cv8PApGv1c6hhfrfYBziPJq8PuNVtdNg8eN9
0hLve35OvwSFVzgylw8IRswnx8SYngh6UYfFata7BILh72NYwqtSFtXXop4xqiX9
D3TegG0/GMnDb7slGKWx1AYF0BD9s8dY3fp2tKosoC35wSbbnYAQo5a/wgHMBkNj
KqWzYuNQKhzbjGPc5rG4dtqF0zRQHZYDR0g+EzDgwJGyT62WhW2w8STksmZyUOCP
VrTyy6cHXVD47aQTE7iLvEX1s2LfnzcR6JnUKn09/3a7I6QcVomKfkzvw3T1+wDt
pnjbL2fxcWcgRlVFD2jhjUk/Di+//BIft9YRUxhD/Nw5d3kSR9izNTMJnYQmHtyx
wX1K1QzlmigEEMfeyR+il7UE/7RIq5lDfb+naNdcsKWgDt1TSep2fTBodJju1sAp
HFOUHzkcECX/yggIYLLReYTjAcA6Ya8QXDIDj57Kxxb4zo92eRiBeKGnZagOvlJt
uFIRB8THhV2fNFcdXA8MRBEUGzJx5G8hIlQwYiVDzjnBljFhm15KOrOkQw7EQ9fL
rvPCwsQGwaAdnufpj0HdFgKhti/PKD9gXaanEeKdUGyVex95MSY4eNWuhz4Kn1d7
Mb5JYlPsxl7lmCZGDzVAznr4PtUvean/1x/Bd24ZhKfiRZ3HpS41UAU4XTFagprt
4DhwQ1S+JdB36AaTCcn6+LZbZz0GjPEbSO0sJMJcTZtUGvoW/nWw36OIsEAmVDJk
DK66jW620hFj2wcyGEkQSEPKplohTf1wjs8NZMhTD80scPynibSmHtKpZ/335IKB
EjdxXjzDSf4EiiArtSeg0T0c7G6miq1lA2ZKkb+h70cJpHBye44TVqnQC85DcqZw
7/E/kpmGPBHr4wZcHT23eepcALtUO34TbLuxJ0S4qr2cKvRJChqQ7Ou3vq+r+us0
md20+5aILEW1EfbTQjgMOMZz10kpajStFUs5/nSnVli/okZAl3l1NvnJWFME18pC
5efigX2M7/eQbDs93sDFc1S1kq8Ogx6h5/yUBFhDowCVTBn2L8MQeZAVUvEvt6cq
xy1fXTASPleTyw+dNnR//DF5iQRFtil3GgouEiRprGCppmooL5Xdh44pPz2suCGK
e5YHdrYQMkAf1P/SPRRVSfb4KGIr1NMfjAIOUrmdeiM5RKEv5EtAUJIiFxHRfSfH
ERn4s1C9OG+cHpvxY+PqoKsoX3hOx5hIk1YKayqhAoHxcYQiqWb6mpSrF6A8CukB
Oia8Inh+6j4TkjErMugI5HpwPLgnjEZE2JXGPM/3yOQNfDT4aRAgoY9z0YpHPRlc
wcVeQhGfX6gkVzHG3SSnD6qI4luexk/3mDuSJKXbvwvFrwFAM7VypWYRl6EbXDzu
htWLb6GUBOtLEGMKeE3xRRZHH+oyUxnZ6bIqvIWAlkBtkl1An+spGGkb1A5CLBDD
xSjTqeeDWzw8sPl7Sf96IdFqdFREDlU0LJZ5ra8GujSnoSN9LQfRNEeC/AQbWl3F
MF2Nsn5YIn3SojjXsy1sM5OXKgG0EYa3OJ27Zo7FoxCEAp14PF4wx+CqdTFglkQq
xBc12NBN9IrZxggHT6ytAmvg8BrSY9xtGqaKma/o9XcIPuPxbzCBYMRJTnh4vd0/
n4qto47+U7XLqIcxRnS4DLYRVXD47Ifs504P/wasWZ8MPkuVmCBfxucr8r+nE5W0
6RK4nntRw5QRVetHObA3jJ35Hyd4qgvT5odu/0HPU7Zvxvq2QP3DfnUlknWZYTiW
0wOroYMqQkwpGKtomzd0O2O1pToYXFtvvPKlj7gkUfiOnkXMDrYa/nTEYQoNI/L8
Uud9VBGc6wRN/PGwDOSaot4lU7xrLAq2n+3uoVQU04hlOGF4t+5QvSNURIbRZ9AL
eQliWxbtKywkcSEWMrbkTrC53ck1GZy7e7cAtcRhilGwQRGb1wI9hJaiNyS2fQyo
ODBJgJTGAso7/Gk0klPAngizEqQvB3WfSxD454hMup3kxVUHEKLeaWDvc07e3OEz
j7Pnx8ncVh45/1otkoFAdJgt0u9MXdglgHse79ziQS+qeZCvFlPHkf90htfaCGO/
OiutntG6RVmGgLPniFiNAMimdxs4PgXafw7Fjbfo5fEe9Lul7pWhcwaiWHuXFhgo
TOTVwN03S1Wl7x0/8CMEUasqX0QljeZcStqpA+VJAtGtGiGI3n9JBB+LF7inP/4Y
9CzsTiYoyp10K8Bk/YwzVa0sW6LqQI5l2JNWzeP5dSP3AQl/0yl9EmW76UaEA9Ev
/v8SCHuJjAzfWcTAKU3LSaPH78k0fZDkatl+zdjNxsYa8u4J545jhE7QUU1z93kX
3TBcWMfIaSX7FFLoLuaJu3sl5l2wxi4yYKdpNFE2w1b6mKbnSwZPW2U7eaPAhPF8
L6+CrDH4qP2RtuLd4ooyKTHP1CdkWLwamAWiR1QjAYI2SlR/u3VbvA7Mt87LHGYH
FtYHUZhfrDEe2B0VXZZdhEy0m39lV9O9JPLGHqPFiNQ0CTZIkQJJN0vKvj8jfXic
h8arbTrVYSgRJlahfEuQvQtUGgAap55nQ7QD/oeJmsq2/SKue+XW7ZpEeNhNsZaX
lrxqhpEboX9+/u8wMGlXb1aYo0LGbIYlR43vaX3D2B+JtUOtdATYifV4HlyTek41
JDtbZhP2ageTr0hUgX6v0OFIc2ZthHCSpHCrn7nL1PTWbvlhmjpIOV4nhpCt8oRv
YGt1BaXx+9+MRfDfxr2y8Jeo1Jab5kIhROVVK/lVneRuxi5Rf9nxuY7aQvv4n40R
8AuTiJTvew/8v1IuxiB6XTOF6oZerngF8NnWGJTnZE8UVgPOqPcIjzhSEQfsbhZX
se0D/8IFyF7Fqyzk9Nq4PbnkEF+EuEW4J8tQsHxTF/I7Elt+hR8Rost549ls8aTP
auT4lXfpfljWsdz51FQhQnWjxdxA/0urnkuJoPUCeXBJBLRwzQo8oQOQ48/C8fU3
4xNSJM07jA2+GtJzIeLgxSPfXmq0w0mojaKSrfx7dqQI8l6t6sNl+v6ZoYG4xqZ2
M1n9na8vI/OwiYr6uf5HCV0FPkfAMWGV+jXHM6muMvzID6n5zKFFFv00oGEpviGX
bue8QfkiZM/nxGREg8mk0jsyEHDVFsXn+LV7xvx/25k9oHey+O0C6T5I2sm7heTN
UZ3NXJi9uckfEgssOvAikjUTPk8k/9gwzzcpPKz6PU22RHArC/H6XONqX4WFVJd6
YclplI5wsbnticu1f2etPsTA2EZ7DO1TGkJuczrAnVf29tWtcDw006xIvII3clTN
nFqWjE0uNrVTsDy0PpZBmwCFn5OCyVcpTMHvASbXym8L6SIHEC7Bdkr00Ey2K7Xj
R6yLQT0jCt0NyJJZSyKkS306NBbffCiUB5pK9W1TdjZIVu32lHv5gzad67kJLjLC
h69KUuUPE7mHicBrLkaPh0+OYdJaQ8Ak5RWR0XNH+3UDklSrLjM3kSUHoMEwtE5y
aXN62Dy5rvHigNahCo5iV/TP2mi5+SqPqNPNnxLQ0qCPx6pt3ZFLRqwqgOeOcAqH
u9ck+h0bNcpUegUrb4aj7jH4xQ/zku2HS2jaYfb03O0fUsUL47M9Q9aCpVCJ/4g5
WDeCrU1/mrhJH1XGtlzEnOTbd8TOzSc19tC0R2kZxOFefhntDF6OoYlQ2SpxJoMR
oZDy77+g5WNTOpYlpBX1vaM0YZTEAiM/EsFtHM6GvhTz9hnevLzGhbG4f/JDN188
I4v3rs3EvH9y8q5dJytxkYS5Z3B3ssUooBauX15BZqoRu2tqcwhLFo4rOckCJtI5
G4ZaBPw6pLxENvBf4Y5zhpNb9cXghbaDDRG8LpL9ELyQL6MoK/lBD6V00lDIEjCW
vzivJkX+MhVDi/ycwllW3mMVf8h+Lc7ri43mhh3xMWktS+aL0x1gOlA/7jZenBsR
fxpDAQ2RDi4I/y0amK1sVG1HsIJl7/QVanFII+X+Z2OGYf4FeKdHRJZu9FRTbWDx
yTIaVpwIV7/JmFftQT4+QqpLq0a1qfGJR8DcvzLMRWeh+0sOuGuRcA34JRIAEshb
y72nKLegnm6rp8F7nB8hskdOiG7TNH8JrtECL4UeGm9OoMXoeKPF+7k6TUz9GeDf
M/FOzei6d5T/ehspzRt2eJOCCPJ3DUfUw+UJDNIhNCywBE1HA6kpqsoAMo9SzpqC
2/xOtWm8nRFlsLQi77gnQdJNQEoEsVAg69G+cqBMjQXIai0xbIWpXluRCjNLDYND
0vMJ/6iCSBbHShRnz3MezDhJarkkKGfsoImjxDqKWKCw7OwRkdBScOXU5bne7HkP
G0sBAKjG5FEkS/btATvepwyi9gDXtCnP9cCMontvNaZs/hNwMPt4uvntJW/jekI/
zxwlRM1sH9P/XLMPJGDxBMi0xqE7NqxSl8JyZ0UM3pV1fss+acWZ+VqoytLcoomZ
CR6AEYFrTdjVo5NaGE12+ojgWCziis/zcgklcUfzvFrWX+2zks2GPNT9cw/n6uGa
JQvP/SjI4ujSM1PAB0tXDZ796VVpepGJuoEFl1P4ISOyPzM//qAWWfWnZUvw+91+
PbrrqAiYXCjDnKglzOISwrkYO6cPcOrKaBwksSFkLEYftdNmaBJXshfMpNe6zNFZ
NNaXBnvntBO9KuttR5B9EtL+2KP7mDSr1jVEM/YbAWpbbGQZe8lH0HTsfBRaBft3
/Hft+aT+HbZ96Jn3NCkYC5k9ciECXTmIM7eH7P/IzmAMreIfdiiKJpba/Qa208AK
+q1eqZVUnBDTig+a6XpxZl7tvvpSWx7dC5TDNObEdw1n4TelMUQyWITsaScObbrf
t0ghPbZ3nmvKNIEguOm+Cc3jeBEMzw7jQyBZFdFUEtAkeYBhXTaP0yXVWE/4VThX
pSu4Islbddp/p9pxQP/NxeMkr8CO1h5PEoGm9hC8xcseC2onvjQyOiLk1k/k7Rzb
od9F4ZEnY4oRVUeS1NmogQ1vwGGeulO2YpcwsvXA8e07oommO/d1fEJ6JQXMfMSK
Y7bJviSug2VMfN1e7nxXBJbGgqgCZZiuVGGQq0QqHlFb/7ozgwDfrc+9LKgKexuW
U4SiaazcJhnYaENO1QHLc9aunSkwbSyUDeErFZdjmPJIwQT3uinQd7vOig6TGUbM
d3mq5vhn2qIXHzsf9M/VUurELLktve4dC26X0Vjy4RGDF6V4ANpxt+zSYIVc5gHk
I7WGHO6vISSgBudy8Styl18qSWukbrDl/yueoI9IHZfYkugnZlEKoe63KMKMtQ0g
PdXmj6csJDb48Dm1bFdOO8XOBG3EvWcm4i6OxBZQtfB/21uZQUAn4GHvaQMWABas
dSki9chbSLWUJZZNM8MQxGEfnwna/hmtzNw4RiBD+Hwtp5+LpkM8Nzd5sutKBDXR
TC4aECy5cDn/H+WXOv98+vZG4jQunJYF3fWilLD5QUEoyDr+WcqKCN4yf3AyTLrK
U690pBaxHQcv+S14FbJqhxtewrH4vCvLNUinFS2s0C/h0FMQBC8ZJynEV/zATb/E
VzGjEa1aXd46Eh+LwyeUhTD4+ZTytk7nkVHZ6Ndv07eQxpzkVqYtt/8UePms3Aah
U90RP/9rPYWhIW6sYl0nBNBnZp4VmR79Yqhe0Pkv2wfSPim9q0lblWvZP+RhYJbZ
NEDSkU/Wj49GFldN3UmltmhKqwKp0QMHUvi81f/tTxKDFAnBGz2yj3daDtGtI5zd
K1TS782rog3FPA+0XsmrZee2GmMlob8i5HWS4tGfYJx5rFYQXHzVraROlWeK0l3i
V/HfNocHn+ZF46ClNk4msg3jbEsjbt/Y2SsEAn+MFws49KKleZr5OGejGa7XohFU
nhS9x/NfW6Y/3z8Ax8C/9ZF041S/H8ngdfEfMjZPStzxwHpTMOljpZh7Ekmg4g8x
AD13aEmxS1OlGxwO2iCize8EGB+y0g8IvQk3Z6zyYP1WPwgtR5CJXBNRP57W+eGr
wDyQfQQQvTv/MTfxBniYOQJv+dLj956xfq1eNxmn71Gl/eRuJCLspU3PfBPTVH3X
vLbYsG7RQAF4Wgoq20HYzh1qcM0JaZ07zDoCghQT7p08+FvaJZE57477iVXTEyB9
9ZUyGlrdjGJKWw9MGx9w/87gDVW2YKCi5Eu0/Fxv7d90qiGqrN4Qgk7F5oW5Hwfu
diY9kjY7yGOFWPICniqtY1SkqrZrOiGPVJgWSku+OkZDX98K1URo2Clqp0updNs3
BdhXkUEzu+Audk70heodrojj85TJUS31Z/Ev3VfcQ2vG4r4rkbbzdFlPBWEMhtI0
AtaPbGFkj+x+MFV6tKC23xSpoOXbWDeTuAxouNKKHlhFC6TmLcBmFmujwHlYl0ll
wMhSBcapY6wmvldS6Mt0EAkj78QqPei8Ttyk4kBfnR+cQr8gwDPxIhcN8+/3syzk
fSWdhURxtQE36+mipKWlIGy29SW27znkziajqp3G1bvZwYV4ZZwD2bcFecy55wLE
6qkWOTCY4CkFW/M9U6bxk2ojjGtTrNz7M7GwPeubvirgWDadDqel1ha+8y/kXdRj
F2QlVasRIkLHKoEiJkQXE6nGW1VGDXKfgg3PXRX9RuFXsVv+YkwCnxrfinspwG4Z
qmqT+P6dDbvlJRiwRTtzRsSGqVhJMkT8itH0XEuMpjad5L7KRLVa8cww2rgrLG3g
Ssd9BopzfJ97arcoPhOCqHp9I6mP0WdX8b4wXQnEanhcOb4opH7sAA5v8e2aR98E
iUTZaI9RnGOUd2AUMZvC37lw4seI3QwlPj79ZHcteM1R3RrFbAzsRl3ZhB0YTsjT
XG8BB1Ui9w8o+dQXEsiPfAg89GsaEVKezpdiYi5FK3cjEIu/RY4cEHiD+Y1Shg5f
8X2GHkTl65ZxkAPyPstPC04ZwV+mbTEqJaqA0pHd1WITWdQZ7IPSPvonFhb4UJpt
urXLo6TcGGYE86oh8OLabMvsiV/9fMlbldKbpVN5ppDqEdloz+6NkJSN7BOaI+xT
a9al4yfzuNzS4MHJDUgPND1VQegewfshPO8WTBwatb/XGKO+QvmJJ/RXVnfCOul9
FjCVqaHounqbF+b6zymwzzvJsAvizRwyIa2CKVI5vQGsdnMh6F48Ti4zemAWiE5f
Rh7sbFjBX8eWXUX8PvocJid7M2IJuq1tAhyIRFx1V01lOjUGdY6fp9kZys1irAvM
nEjyYs8CW6TpCyEOQrd9a0uCzunrVFIY1HD11cCanYa+iLE7s7zInjATDT4EvUjl
gj74MIaHuF5B51oAIWGJS8sovcu+bjTvyScIWO6CfMq/kIUQsW7E5bYvrnxzEncs
hCKcAdeUmNkNNUKzMrhi9hBYWGXXiE5vmjLZx5U78GTfxSH6xk8Ed769fGdtyqNA
i7ilCcSt8lKDtqtYgSUZiYBiuWJ84UjTbxmQ1odLjU8ud7Rguac+CRGGgySlNLOj
NY5D8GYew6UX0+R5aw8c/EWcJfckn9Bbndre6iqFyQTscK7AlSCvvdoP1aaLnd4g
pQAsZLvXP6oQl8PLIwfoPy1ok+p77ifcpDL4darC4u+43cKSZKLgpX6UO1Epjk3+
siksqf3/PFnW0ZFGvH8s0+03kexZyK3S9QGVAVnQzdU4aNR9A8zkDutrhtItD0yc
YrGLfNIHAtrjlu6vCQPbPWDYp6HWbdQQs98aRE7hSI8TdBRhynhs0jQq2STs2roU
LyC6ajf1NpDgXKt/5boU2CvMipvVNkaFq/Gzg/sCG29gQTCWc5iOXCxBE1FaCA39
x5ftqXh8hX/YkF/Z7p9gdz5SL4i5jxY3YbbBAw6TOIjzsylv4IWR2LPhqZQqSAW8
tstJrCtzg39unGGWL9We+IE2tIuoAfP5083+cK+dXfwFZ1z6s/3A6iFI/qW783Kv
RkQXyOjmqkHXN4MgYhT45LID8IXADChkNVkain7AV8U3yVWSbFcOq27WoEG5RXgM
IEXrooBLoTgBiu2n70rWLY5+RFMdqgIRxgqAih7kLPMg3J9zO4T55KmT+SP9X9Pg
L8ERHOSImAbuH/3DTyQHUDwOyEDA1Uk298fWIxTOc3d0pQovt7Z1mi85K443oW5U
8D3Ly25OhKEWGlhoKaR6Rin0Nj3Fzsbw7p+5owaAThHQUbuuoUUbWUY9uYt9dG1z
b78sK6O2OcUYAIFM7hvyRYMHZM4B0NT/854iqe2H0sYBaJBDjUj83E8gja1XHp2o
lWrzQqwh1XUkTWWlyeTZ9YO8Xqx0sFF/z3VL4SAocG/9FF4FZ/bwAmAJrXwLOJD6
//Ph0l64aODhhzcIykJqODaYDtQ9mNVj1gbC8rGFmKpxaQT0KR/4ZlNaj1o+15F+
+UhUC47Io3IUOaD5JcUyX2ef+jm8MdeBRteI/ZAdF6yo2ktOCFqa+XTxtj8FDLdC
tA0o45AvIc40iUMQPKBSAdfc8876K/r6eIQonqLVOo2OvZzJFvqb0IOdoBSZ2MFZ
WR1pEJVsA2SCeaKLa3WEz8o5hq0gLQaF9xp1FICJWJEAUIEsjegHogNlRUUoELG6
kbGW+Tfmj50felHiayl1VyYDpHqHL2J8JTJL0m0xFnaasHCPjW86vf/2M8+mdkZw
pF61jFu32srl2AJZaBal4aH6TYxTev692kMckmNHGX7x56T1x6+lRVvudUHBiega
GGCQo2AU32vgzL3Yg8HhW+j24Uv5XMgaiMrxXjKVUIljGTR7YXrRF9rEgPL/xycF
th987w9vsFVk2E/26rLnwvFpOELBsY2/X8BZlCwmsYx319aLhKPV8kXzMUKV/u/m
D5rAQe0hRZnCI4zY74Yq8V75U/kYrBunlyzc6b8UqmYeORtqJRmVb+Kkbr1r0RiK
SPTVvu7oX+ZAGby+QUDzkYNf1MhnWkzCcY7Q0z3wOGXN/4GaUIxXOaa7EQgB17yd
iHRQz/KjOaM0Awx3dRhc1XQF/LPP3BjaPh4uR7sNCC4h/c04rC5LlJdTqKAc/G0G
ba9YRvVuVB88kQIf5I/98Q98VfQ+KYAJYM8GVfSDFc9+6E9z9CL/uZDlJjmUrmO0
q8l2FklgY0VNYeaZAONcZnUrmjm+1rnH5mYJOpdS+KlV36wNlWykOy6s62YVzvqP
XkSDJW2AEiupS835HUAktXapshPoQKr6wSUomUGWQBNlM1bkNjIoO2MzaPSixSrc
r0HCd8IhikF9K80jbmmr340i+frVWaT5Vz3Wb8vVdLdQq1oVuUqpo+KcuxUzJnFq
/DUUoUdWkDObRKej7vhlFo4nViVZfJpitfLvgiqwYZL5x16eoSTdHZ2bDM39OXKf
W13XZ9jjiyEPpsYVdoxpmG/pQWs46PbOgwEU30AO3253xl4shPoGbRWUhexUX2aq
fchWYiWxh2df3ax8iorrZoaQHjul6WxlmXEp4syLAywZto8YnvusW2RaVJacqBH5
k1HfpGi+1MjqNjBeJXIU78LPQQI4gy0lDTUpQJtdT3oBQhUA1VTXbvYHxMzC2xdN
mo01xOfX9hmNn73fzV9GfVvLRwxfas/z0h+go1CIwQss76LlOS6Wxby3dkty6kBj
OMVy1lHKxr3wjbpyZqo4fNiAGQ+8xLdBZg1O4wE9+unwObMsI7RsOLVxYGbj2Lxn
Xq4mxpm2+BHQejk3/I81l9shT+Ro59vftO/Gcc5/subCtXZvudVIbh6MF5o+4UKf
nCtB60CfY19C8RbQGiG5V+6fmemmvJmkVY7shjC1TTn2V3BBYqoad2zOW95lmFJy
tKEvzdFkgjVGf5+S1IFepJf8UZzHIstXMqmZ20ZDeHhm6hl631LktPq2liO9snGK
Wr+GMGfl0nL6ZmH4Wj3E4gAipME5KUpiaSkOtvmL6YJZcO5n6Q+aEshZ1ici0/T5
O6SVBAnY1e6eV3aZ+/kpxJBHsKMxK1w1GrYVoqkY19ahr7AY+4Omp0seZFGha7UW
6k7iXx3X16bC+zSkC7ynKQOifbMy7+f2Dwmk1Q7J72ACAhIFmdDRsfsP4hDvUQGg
HqvoOxu37TRUidiKhPLvaY5IdBB6JjXJu75r8ZKGMAti3VHjYz+tW//GddcUMwMR
EQAMh0GECCNlt7KkvNABxbz8hmmsNIRehgLwbPR31JOAAqJfcSPW9PxmQoLhyu9a
6D5OuCmSkgx6nTLtDgDhzTWUrlAm91LvVHGOOKsUobwviRrU5dR6REwCTTF8K+E4
lLPjEjoYC/3QuQKNzKE/mRvrVOtkedY0OeRWHfJqgYrMF9MC5TLHpTzyBqV9l//g
rsHaisbpfbdUK/el5v+X2JxGNroC3NhODWRISNPYJ1qO8JNrukuqwg0z4vuwxaPP
wfLFvyRhbk1jM3BkPM6GLCi2wqlFTTkGZ3oeYJe8PoUC2c3u5PClHxr5IxZAa2gY
JM3VB9pRCheWbARR7X5qcFU0GJPXlfPmuHvoDBE50f76mKdVxzQCOjbws4jpL1+2
ywjDLdSVCmmurKRYTMhsQNNm6ej2vY/pap8wrLqN0N0R0Zr/ET00VSrD5Rbnb3Zm
VpO9T42Ymz3TUbgQFk6ndyA6hh1SSmCsF03urp8WM/FA7cb+I4tq1cKgt3G6c2Z8
/K9M+nJFbzvcHpqvnf5QheWDKe55XrVFJ252AmlBvcQsFSuDXI/6UxvP4HJPYpIV
ZaWD5jDwu32XiSgYA8jV1Z+plOwVZCbRG1eCJ+r6r8gCcXz8nk5gNEuj1dQLB1V/
SG+yvnjnFDCAOq9BFH1nVWw/z7Lu8MeQWgWO0MkSHRQfAJ9baVrLDY4EYffoKo33
NhNh01m9+oPVVQcRiJGnGWiryYhC1KXV0L83+L52a4d5k+4Iy9kuNDdVd6hTLu/I
c51j2+wlvwf6e4QscrWXicJsuYqtOKw5D0dGBsLGaT48+PrY249Tn0KgGzILdOjK
syy56BIAB6wzHLSiJgGyaHk8aGeBrQHu9iao2qnH3hPqSWMQ4FW3cIevhbcW1mXg
YXKZhJiu8YMunMq7Q3JYMQZFjsiDR7i4Vug7Pz2dahHE/6DDLSMnIzDxtFrgdrk4
6xHUWEztJwHjmQeMSkBczh/iobgIZvBkfJH6ua+vSxi8sgCPE+rJB8NazY9EpRbK
tXDGpgkxQb00DB8GtuGLf1iGNZj0wiMAvLQuSFRMWjp8ETuF77TxUvqk9RiEod4r
jLP0ElY+5s2K36lZgnFA+48H00pWXHjXR3XSvGr33QH5I+dnr/GIK2BkBVy8z6nv
RQ+wpC8UPXOIOgC8bwWOA9dl1zRIY9Mh19H8fPUDQkig3QfLZIkef/cIqLomWA9Q
GpxQJmUT2QaJNWyfSNQkzOVk4BES57ENzWdrw3kOsIcMyC5aTkZgsAody9LPF6R4
HugWzHrzFCEidoBey4/S+xLHLPzRq7gjbiYpReyL4h5At2uTkUPMBb2kRFeNL+v8
gywwauUbwKmMtWPykAVE7NJdQ9hiGLoelRrU8YSDcMB3onK27hm234f7H8NGAqHw
7IhXrNERp4JpIDzC5V89ZGtEkTQsEvZiyl/8+Xnc84j1F3H6HIHKett4AbIbN3Hp
KiN1c6AJg2A0oHeeLl92omN/n09iQrHe90rB+VQhOTjgY1gvtOcBIS9ZU5nPiEce
Pr44DXXTYbMAS9Y/RFC7TUqRmYzBC/MkGAqS8ihP6zHEWNCojMSLDDJ7C/bqdedG
oBN5zv9JJYGXaFCcgj5nYAK3Ox1lzA1G0QyUWepq3jOF9UBy4/s9ZVhteEgldAvB
gCmh3DfJd/p9Xi3UIbSr2wP+8zTl+NEgY5xl3ZPtQ2LIZFT8mW7mDI/RWV8LGf1k
OK+kzXB8R84o+LB9rK56WDVGKg7yY81VjpfBLwgRHMbTvtLsHEMiCpc/Q8cMCuai
Ay0YzdQa2ZpbwczOQCE6hnlb6ni3/hF7KT1fNzHHcAKZ9O2M8NJQpr2ZB9ajH/hp
m8TTjxwtBxqW3SyXuOQKnoCa7AO64SJ1lATHVLDDKsFFo2P4Ki0V57pjjesCFehi
P7ae4dGkzVCOrWl2N4rsBy0sn/40yrCt/e6kNbXJbQGMC7aEM3SjFiCEu4HkHG//
Jla+8o9e+yEf133llPU1R8GcanW7FpNqW2f/2XXQZH7f5kh5ynfpKRXcPk59f+fp
/MbyncUNLHVBTRf7+pZ5cljbw6BznYi6LXPwZpUYgYqcEz3DUSME+F/LVPqKXtFP
f7u544WjJbn9+ieKAxMMx5hUDIt8MK/qaBTf46kLoskITjwvVYdL7yNn9HhNWOPv
V8Q8O7k80dwx5yZpmk7XD+i2l+s49eZ5+RSTSfbeBkdj4xR5DOmto8unF/PQiNhU
7giKlfgA46BoZ4D5YWCEkyZosgtpNtIxcrxoOEjgExrYXrvnlGcnxRGY+3PTS9F8
q1WrK26/A+fLKgI34x4p938icbpn5CxsNCix5J7O6hZjlAPo6IiegVJjKy0xQSPX
leurdCLqkw3H5N0dzSXbgh73WabDIjthuPVHE3zai4tpP7QmKylhj1LYagkqKYEr
V42EA6ijh0eku9RMf3O3CvZT4m6XGusVH1wiDfz5VOk5v/jcfBeQl8zif31HOHs+
ey11992wx0rG8YghAfFsbQb2xYMhxvkc3UQH99mg9IR65ODUPMW0yQMpvXmP/CRr
cOwf19uJN4A0fYV6c6Hp99TcaMAKXIJZ0t+GpxgFvhWP+CSprxvENcBXgVuw6xi+
e2rsLyDmuEY9YFn+sVTGUxZhoFn5qmNBRyrk213O25yGX33dsbomuI3LULeH2OTB
Td28cGpvTlXR0UlqGgbenXbovTUi6Y9BISmJ7Pqqe2BaFrxz6smvw+epIc7G8mA9
Mo1hHnvVfq3jO2kBpp6L4fRD3FtOktUtqGdqhoMjiMWFjYryP5dKLOt9sDCgMGqE
XJ6R1VeO329xcFm/R/JkQBMPPVwOcaD2s1WfK7kH4LdX3lm0A0d/cK096G0c1nnM
GExDxx1vcjLm9s47c9kKXEQKma7IZD8pyvxn4AkW0nS+qat6yf+cTem2DyJP753v
mVlTaqTXgNIPxN47WImtjvpiCgEhCpo1RpHYTMJCBIUAeiTqlrQrAVZ6CV4aKK0Q
AaKPvStAg8Crf2V20BpH3IxroxmAl5FfF0BYj457RJjSNbeaFeDzssz3RCyf2OBk
N1TexeISQrnVzec+YszFhkzYv5fb3YACxkhKgSs8nhHSUdKLLmZ7vdvYaFwaky00
FXrblUIEgwll1Bui22BAL/naK++md/sgV57muG13qo40ejD1PHeZjXgTK6Q0GgTG
EOLStq31wSrUqdUzxESGsejXzeEvP9TintnWYBETMa8nSlfkXCsZ/gAPB+aX7Pxu
FuPw5PVFf4qcV1gK53yBlwF1CsNkfrINPHbsMkd0nwOnztTBiyq8/PWkhmwDCpIO
GWThlOVUdkn8iL4f1XoLIjtSTjFOAs0l0a/39fEOuEDltgGsBVydQazTtLr1vHCv
aF4amwkbKHOSwlBiVOhvuRtYg7tPqGLQ6O0vdt68mvIfqRw1z4yR1A1WlSM7788H
9PtR2wWNvvrk1gEgAT3FqOgnU6JT4DuSuGVM49JUYAktldZyiNsxV73jOWUtvOeu
RkasZs7MbQHXIcQ9cDL9iePO2v5N0bexsxbu0R0cmOH7jeNBCeI6qa9OWumE23uH
mFnrpRIbZs5JgGssEVqaUT2Suh8BhBGo95JSi+DtxqAN4914DcgJBW1nThGb3e8V
O++ymfBVmjq+EQK6AmrGEEC++yCTXrGXKj6zulm3oow9vhIH9kQ0PPpeJ0uK3bNb
TmNyTCR9liqm1O9mmbAlrK6P52PPrLnWP4g5i+Y7tlm7VJssePLX5SWqI8UbH/4S
RZ4twzCr60cnb5vIoFvlTMDjmAiZ/CgQfKxyybKxmZWARiOPeH9MJx+JWRCGewwH
S0P12XU5td0rkV7gAltJ2dBTv5V+uflimRWP9yYqZUEqMPi3W0VSHauq9qHrBGl1
AqWuPgLOkqcvb9NyfEY+gG8aPDH+IluWLhtempL1S9MLlOs68Povrp8adPU6CadM
CPRbCzNfiYqX3Y7u6jQTRc3tJV+xTH8mkusyPQeEyaZ53l62exdqNz8LN/0E5XtP
5Bq3swqhrdc3LwtQ39rS3oPGHMhDFH75ls8/csEwjib2iuN9PGAecQTv65TOFEAk
4RIRpPy4xQDitilyAFLaRka/S7CpGzh8k3KQShv3YXCtDQCxRKw1Cfc2ZbJFZqNE
OL3MqtGjelqovWIHjdTk6tmOgvhuj0P7Pax1NYupX/geoCu8tnLsTUa/tJDSVfl5
EQ5FL8VIZR5lPsH/RXmGyvNEdPw+WUb5F3blg8ipxg42X+OIXOqnxpbttIVSs2ET
subSFtO0wPR+D2Ppf0GFmCk27IYrb1J02xEfXr8W1a6M+GYywfv8pYbBGIYsYhEH
QoDNu9Zh2PU+cdYOP7Shh9jyiCGTUhyAo3kiRzr+B3VysZsklvta98l2+6oGVZlL
U8uus9hXJ5TPyrm67/K8LOaULBoPFREKLXe+i+tm7gzG1yRe+Qv9CXk4aRulFFP9
P4RZZ/mUVOcDUVNBYYo8s3vNdDeVrgVDFu0TJP/ppq9uJ413IE9lhxVMUC9m/sV8
7xu9czTPD4ZLsh5JQR6vaj3s/KEGhwvHeH9wG7Y+V7dBZPUuseJ24DzLbISHc79l
DIwggR9E/zuuPRdL4KL5POEHOqCY2q+2bdsAOrvXFBN/AL6Jx/gwG8HFc61ttyxq
UpKlKJNFhyqzNmuq2xOdONJyGJL+X79Eku1PT/LjHhunVwGkvFBuj/27WUh4vTT9
ZiaPW+087JdxPPXE+GR5g9fhreZ8SnZ7nKocZMuD5apsxvs8UPwZ7o2Q1EtrWXKh
XEm0hMDdpqTkKxhlkf61EFnJbr5cECT3kdymqv4CIaWR5sCbpp5ubiRhXUzJ1pSW
MVXVwpInSBoxlYOXQNFgYs+5K6oVwklvAvS2EVj36Z6ewGM5MKDwMLeS4m2IEoGR
ICbUWvgALtWDzrknkDxciNgY0IV+yUDwztWF9bEYNKzSKkHjzKkHGKOx4kwZOsTY
OctmHG6f8LsFmKouCJblE9+DEbR9Yo3BE+G3t5Egk40KGLAW28QfBsJcSmiDs8Gn
mRc31QPdKwQdmL5TbHC8yfkVKCmpzRyE2I5+U20cn4cSxhU+6iy6aFgqvRifD+SX
YVIVqXfhvpOFNpiKnnny6/SHNMmxjelCDe9R1vPk3Sl7gxnrCDoaV6CqNzFhUVEu
mR3yx0xW/42PIZnJw5aepJkSo/FuxbqZ2ZCluW8W/tt6jNBG0gmb7zM1zL0r4izP
JGrQiG05jEqkjhuQ01y1XxGlBlb+NpV7p0bbHklwjw/tNa+trV8MJQmaf8ullyIZ
1/+NURPXpBvG4RBJHbLzAWF30gINhEFnceL1hA5xrGaqCi4MecZCxR2N1+YMwzUf
Rn3+ZvSwmhiHPwI/lmisOhTkCZx/QR6YZpXld/w741V7tTnGq5+0SxvQXzqqbQXB
APe2ZLxKQ2aVy9CMK7WQhonUvMMAU2Xi22ALehdTibE3FolrkBfsNsPMC/AY26q8
Rt1yWCDxgsuA2NP1th0Yavq7njTWwzQgWPaK4OLgq9nxnqSdBSgS7F1ijIPEqJbR
L+TB40nEZs3NoQHd8D4zTJImm3jp5YrguNRHDlvWaOXvtyBclgB4PhqmHm9+HvDx
OUl8EhNHOmKnjHCZQztb2DXwxQMBYUQ2oldklOjsg8OMBsmUuo1CZ37/M4dqWUQM
4HPemR7wiB/8PsOjUBd3/n2VtQMNSWLHakJ23u1P6R7z5pKZzXkh58mKuoAwmu1S
zPT/ussazBksevFfGMsLEp/DpVfi54emFPwJYlNVTEN3Zq1iz2kCWdhcS6hX/5GT
xjSN1yNMQ2LGX858fizjMyfdMR6log7+VS8f+/tfDmA+QKy8PYjLMKKalR3GAZ4/
Xpt5eeGfE2Fvk5zje0OMiHw4inW+B1ZV6UYP4jGxiiVnOiA2TGGD6AO7andaf5zS
U/2RwpoqRyW8VhVDhq13TOy8FWz7G4lV+kupYIoKRv/89wS/FecyhY8JGAuKyPTr
QuJpeP32yNi6cbGBDV8jT9wz6DNywUjKlniiZnRCGEckluuS+jbfDDyHB9R/l2fc
HK7eN7SdOiWtAE87Qo83G/JELZFQRg064y/PKimHNcLSFGpLLw3Z2SB2AiV7Le8Y
itlBqAYDyzeeye0qrENBSEX+loiUH2MeJsbh9hIxO+270Cx+0wZEpIhYh2zTPbi0
xqbyQlk1bywJaqroPEEYXWvGJDmMJHdvvOSpFZgct8WcTsEdoPhC+pjtUcIljrOY
opPKVGRXJtvE0bWEF9h/dRvUh/l/4y4//zbZDCZNfgGFrvN/EoEWbvlMlwzj9+T0
yhTBFat5krWEEd21yAGT8fd59hWwbBFH7Yr0Sd4uCQQuT6SiKDc47xHLnObgWjJ0
Jtrv5uGnaqLqyiei4YYUmHuM9tkJwtzWJtVLrQet7K+ZhCfEiaMc1t2i+hU6oXZT
8CBEwsRaQMrMDGXGf71aHhOlnHp1sFT20n0v4D0DJkUAPBtWvREmLZezZYvxuMDn
hY60dpLiwtd478VQ1yEEPzQLKqOmCofdLBr+DGr0qczxceW2Mt0M4flSagriwkpU
60xAkxjqnwrU5UuCednSHawtXB0bBqeEl2DOkW4iPEb6NzEOutsvyWKE52+J+eDc
kgmuqXOvzdzbl9EOOBwWku/OyLgHc/IeJcj5yL0HZm8XDFVPXs1rFmGMOAFhE4Yg
c6PK5YPAaLCUFQBtltnhaAAA5r4kgi00kyJOpeJvM4O6g39VErogjwr1Qm2awe9H
/c06S8TEeZ0oTqt5c7rmj++25XIGlonfb0bE9b/J6ivmssPdJWkran0fyX/4FvWL
+uHXfTrel1zfmmQpFZz0fEb3mZehVbPYrSd506YZAlojvwbSdOa0KwY2OekEP4th
09ZbeKfD8ukmaQNcoSLurayLql0SzjQNALS0A4KtuEZm51fdwax2c6ZNls2Hb9TA
p+V7oVPB+zoJbM1pYp0DFJiyLC1Ep6GwqFqRm423vg3c6FAksHBIYIfKFLGoKext
d8XxHf3rLyANeu45N8QsA/xfWq/PUq0nzgfRa+3qO29PRHa1wlCQ9Y64xH+pP5iN
LKZdiWqJ28q/k+dR93/xmY6+TO5JByLWH5wUw7ndubTIMfj4RNxpC+CJmjJhZjiE
0wL4DS4Y4Gll1PrDLeVGodmevUdFltDDtGYx7JrKOCd0cRYOKKjQ1+cC4WfVmMFL
ugG2ZWcU5Cmnmz/8EOXolgkZ6/Ovv/oF7Z+ZIdMKV7/8ipB2srpAq96akRtus2Rj
z60VPi7MhhVFj0SS2fOtFPxg8BqeT8HIsowKcd0fpCl8XVPwOXKa6871YSiSuL+S
TSxIVKdsqaQplj3WaapTyeCrWX/dOjY4CD7Z8xs5zSfwiNw0kK9LvKvCv2O3WX53
CN2eluiw5fT5rAnCZ+62ZQPGaqpqUejLc+wOjViGrr9c/RrUBMiWUNZtCpTl2kt8
uoxzj89uIHg4vZqOOHSujDz0mjvJgwCaYaSPuYWk2PO/nu9e37wYfOkVuHccPTp8
fURLrRh4LytReOqy4KMGNbO/11CZglOXDEX1oLyqCdUxVk6n/EEaK5TFi8BlJIc0
EvO1vTJA8NlMnWZBhpfJwSdxlDrCJq2T7DNM581vO5sHCzTYwljK9WktVPWbdv2q
7ys3ktDRR1nPhz38K6ynlOAIMW7gY8xXMu0h0BVvGA8jW4OWzWMaGAxa7Bijj6rV
J1V5PvD/BBNSidfgFJm1F/Fxt9JsFf9uIOynDyqtNsqmMnFW2bNFPWqaeJtiZjbN
rc1u9j8va67eMxJj5FZ7m99aPeig52oakZ2Po4T8DCb8B2LQ2zArg+tUva0LPW6S
WfYKF4HNeYuntVwSgzsIlZ9L+jlseMC3ruv6f+JM2/OVZYaBAe4PGPCfOnX+K+Gi
ZbTbtfJCptYrJ/hAZudNaUy5X9I+2bcY0x+pk60jTcSxaXPcLyfgqTFPOACqI4a3
L496MFB7h3cRlGIg3ne/92LumJgOVYREfz5Y66EX+fPCM8Dm64UfFKsZHVV23mFo
OGT9cOrSWolqZRRV6I+g2TJwmbpiCICft4tBaSzwOvHb1q+yc1tLKK6nBDebYN+k
EgAfGhCmZOozGbMhMA32vJfu6a4msnfZukucUWEjiuiTAjyygFb2Am6XQ+x8b8Ll
04sRYN4B4yCioyKNEiuq8Omn6lZwA6a3GytZWCoUiP8BQ3/ymwOJaCJC8wmrcSnO
k4qIca6uyjjV9eHbAITCpkyHiWCh+N4JZJHbBPmBvuiA5l34v0vbp1e5Gy9sFvml
7FWzsuigP7Ipow175jLZyXlpuFFcX1kT/StbZVT2STSR2nXWEFDmVRTcceIw3DDq
nknC28GnWYkqdnZsiM1QHjYFS9htsh+d4ts1Px4naBtjFiOXvnt9MuEC5zadcsON
+ksCuxZYzFsyquLOETEtD1yZOrG6FebHZhO8pfmtvxiVJmPidyghXH2amMLSGciC
u3L4BED+BrRepXfiK4YbVZElrfpVqiEuJYbZ6Ly8zprLkFAGKByMDKB9WmIIH5eB
X3jTHGAoiJNGyPwJblgmIxSjv89vX3YzpJHf3ohq+zWETHcJeETdhqYXc6dkiW7V
VstjJZRVrUcM9Y3szxWVQbm8DkMtCRMJr6Pew44w8ZvJgZZzfsKC290aA7mmbGAd
ie3V/jB58adD2VBf8+P8o+HL8rxqZ4cX5iZFAiEyHKP2oST0RTs55P5IqD5IKmtK
+dOn46O9gXdkiWsa7eEJHoTc5kfhz4wF9+bvAxbqhbhqwsUzKVPaitAp2bGYuwuR
wggQzi5S6C/Q0YIwERAgOAB3rWYFSwsudzkYQc91Ct2IiLkw0eLD4wn3sSaz93HN
95CbnJmJbFCVPrIBUuJzvff3izHmroQVAzXiPkXy4rpUBDZTZ91yUEyq8nom+KfZ
fkWyocinrrLspwN4o+ExHaWlIuz2DJPffotiN+r5a32tdiHsLgcro7Gxj23bZrD3
4h4wNBHbeo1U1EiLRl3VaxnYpJZIW0FEi3H0YXZYsNtSvzUFxL6PMKe+u722Vadg
KHFJLtUJFR2++C2oXBxZRlXBeJPmLT3DbLtW7bsEtLDRd5rOZgfz7oDjCcHiB2LO
qJ5DQJZwDD43706KmxpuU+HjeI+kuycPfbJBqdZesJdV9ULohqxu/kNKfIeqQIC/
yvF6DXkDQyk3BWkdsDgY5+0J0WGhSw8UlKwoaZRsxAPTgM0Ag6fJHEZ+UFxGwMV4
5k4HhcQcOyQ7LC45jqU30ITtoT+IHQOM0tVxZrg++5aBHsD/iajkYy9Eetew+TN4
bFpf/67f1ssGUMIs8PGvVe+8qcXMZMR5mMdnQvjit0lR4dWf0mHaDYqoqSI0xN9l
c0PIcAcou8m0YrE8qVYx62Se6G5IocFAQ0lsIsBbA4TXiQWe21vpYWpQpgtboX1M
PFJqqu5blAWsu2WSTiSZFonI8ghu0ZwPqgEIhf3KEev7ARERDZr7SldTlQvs1NUI
IrdPV3jiAoZEuxMavhp1qJ9NIeaQu/MUpKbBp19K7D0Vp7PsA9zez3vogshUQG6J
/FXyoJvibekEHqUxp2mdZaEHGjMwhgh2mBRf1GlYWqC1CahF5cT0vIkrKHIDiJpn
L36HaYYKdiUncAHGqSd0brRMEdCGWqEXGdDuE3mspCA+uGfAwBFNEb59IjM+sJxr
km/aRv8GR9Gy6d1D673RIKl9IakYgyBiyu2QlUL11inMRmjtBn6+VyxANJWsTmkH
yHOO7XmigEjPvhn6K/W7j1k577hA6dNfNu1iQYkh9Km+4uSuyZTDrhmOG6S3sgJr
Q72/8DRE03h2/sIgAhX6b5QtUUJhWypXA234uIfs8olLLQ+7R8iGjOccp5s3IVO9
TwwAXl2vPFCG00EJUxECGqqam/f3aE5EHnqEMtEQwdLZYkZIMzR2A6vLVnkAfVqt
7ENTP1Ty09j7ajfnzrgMlqd3wvObSlpDQa5k7m3f8VNoN6XufDN7BlB9Pmv8ESS6
xmsAgyXrN+C/RSq1ZDNuGjdHAFF8bfTTKqKEcXZwwtykoja3Fl5UzQ8ehjLlsu7n
EapditqOuX15EZffO1iza+IhlNUTiWXA/x8o+HVNnXMijfIEfABcqN/zYiFEWi3h
trh9xTu/xsSI/z6iWtGqfs+zRBv9hMCrCu3FaQ+I1XMy0ej7dU3jgbAvzoVEU6uz
9Y+u4Au6nTQOaeVA+3ucDetwBN0aEyVILe7nVyU+zfIHCeTznhe5AmrnrHK1szxV
XJbhnk4jNltYS+IJalNvYsy9UDjqqf8YkbUx+jU09ByVSuGOUJO2YjofiEprRZp0
RjW6poST4HCAulMeqrlt/dCVjuW2jCmoBpIr8mBZdVeQz56LwuH89ftiydiNYcVD
z2RrqpxMkz+7HBVGiIJHc47Tn9Tuw3HzJlAwsLHAkzoN23Kr9/NiwaEuedgwLGoq
dZmcEWIZ9yMVIIYbtmOlksULDxd9WFpESgXy3cPf/qxT7oIrcBcuHiAYG9rqB9F9
7jdZCapibUDlNtzod4RtoZrNkK0iOdrA4YO9nfJ+ToRTIjv3/fqI7ONWGdmKOC1u
8IG5QJv6lKap73ZEzO6SJtAmDjnurWiq5ikkWSqcxXxngEjJ+O0k+NkPgzTYgz+p
r/kQIqwzjfZ4vJG0wF90svScGKiXt50KPLJ5F7M1IOXz+WAnE/PItSD8KgyhRj7o
elZp1NLMqzG060ZUKviu33pF6uHnj6aYmDxB5vvToFqIGP21IOVBL/AEFHxvIC2E
C9jBevT5NbpAmrzFz1om+4469su9KsZdksFGe/keBRZa9ZJAPwBEte2lQHwA5mF6
1uL0hEe1ggO/u0+M3DYT/qkoYYyWHdggWBdr1Xf9dLH0rPzGHCO39Q2iwup/TkXI
MfYzA8CvUfoZa4KokD/X1kr59GAvXFpp3e4TpqdNNgeXq2+2SQHl2ADh6DEimnL3
G0wRxDmuhzRIirAlZ4IS51RPRV8/oNDf/qC85IEm8CO2fPa0Xm9zx+lcaItCYrpW
W8mR04RRIk0N9M70pTE+UGD8OGtqlnppGzjjt+pilIG/EdjQo003FoOVcG8U5Lb9
IElGylBNqmSbTJpiYoDBvTE+v0PtKyybBAo0kEhMLElGQZP/S9000kTks1Z8boUN
7zBWCIC1voqjOYCV4DqiE6sbCV+stU6g/xpgV3ADBcjRNSypzbD3AzD5fI/cCWnr
5k2I+iyb/11cOczbnKAx4pzRxs11rpk2o2If1CuGSIefqCirDWOkKeVZBumH8OUB
jd7FyLToMsfYFA75RL13iYK40tqqvy4JZAKHoZ+SNlrsnUDVPhSGwPABeITmhB+e
kerR1g3SYAllrjhpwKc4dzjqjfAbPP6lJHotZtk9bnKaQPqVOuFE/SwoxJS0zvPd
NRRD8KMfIBhDpSrqOgUcAizIGVKRZJtMSa+NMxlL7T9j1vrJC5E2KX/xZxMaohHN
Ms8zg0djaBdh3vApFZYj/kgEQlpB76pU/0MrBQpbKHzqbFq4wHQIhOUWrWmbVC8U
1kk+2w08o//YDP6gTcc6S7XPL605O6WQwYa/wyXVmuyMgTfOC4SuTKbkpkzcxlrB
CIFi9W3ljRnvJp2V5ZvdAnUf+xBF/ZRh26dnyd80eTSo12sFDFPP2XJXhPo+3/oS
7qo7d/KOI5ISiQBHZauwohWDuQa9+TrlL2rzxK4ECP7NBbP+baVuv5F09wbKumFd
oEuoXxMA+3pD4JqYrlFBS6K7MwGxZ4DRBrmzMM+5H5o73gG2A9/oK4WgE4HxKGzF
y/xwoNLIYOjbeO6YkQT0+of4aPBLRzYlN4bg+IMx78PBeRfhQDAMOB2O+inYh94e
W6c8bKMeVVYnUkQ5H/MU3HLt0NNDf8yajFww7Xl53UoTUoi1a3oMXRyBhLdOCZfJ
/gD0W7npm0M15h0SgU9H9hpRnJXRbD0L6PEvudZ4p4JVax8docIZWpfSCuJHmkIV
AvZg4fsbapLYkY0zGPW4LyMrY4xO0YEDjpW7/DN9VD2iHMyTHmkrI7CVr4DokYpV
/i0u16AqsjrLNB3/9G6fhDn1v3MYZgOAuREA9EeCZzZxc9ERh2mLQhgob4JWZwag
Kx/t2NbNQlP3j7QdMjRUiAZaSClvUuIa9+G5ZgvHJ1/Aox6pSosRmc3EW3jQeOry
0qqm5N+8xrzP3tzqBE5P9I/W4cjJg73H4dtLfEiQsMRGM4pkSfOVYvexYnM11RlI
yVIshx5Ft9o+K2lLLguIWFjHmqyv1B2jn/BCgnJ51DpauEP1WQPFbx8r8I9UP6RK
BjtVzKEkHAfFpcMncoIenRL+30+JAXDVxVoxP/m+tqP/743YxfuycmvdUoi7qjRL
kAKhz8OFMUvQ7XcIiKUoI4RItN4t5/vNcmIT1HrX78h4Hj/bguexXVLDSa4rPXai
B1C1gkR9rROpbovyOb7o/tWllMLsK/4GIUFMmZJkNcKb/O+lFU+u7p0GaKJWwlyw
/kPyyotlWwcjZ2HSSknfucPoU1OuBx4xhbHIkDgG42B7MK79dN5RaDGvH4HyS5op
AvRsC+H5WNo/Pj+Tx44nabkpqvc9GP5b/bLirbzhVOHZia17DjDNReMFLUedCJWf
Lrg/Tyoxy+cnOcxqaDA0cZLu/pDY5ETkYvjuRjH/yZByvjqafONmaD+uMclY7AWd
DI4yQtMf0/xgGUfsVegdxmjqqjw8b205VIifGogvS6MS/jpYhz9jmuzzb9zwHts/
sWsWgdCSCRyvjUaQqjhdGmu09df3Cip//RnvkFusOdfmOmCCW9tONDbrOBy1D08U
ot0obbx8u/C8OCLAOOaucV16kthKHX+LaMR0LQ8gWY4RfWZk92j4tIzzCoX+HttQ
kmyk9VLE00tTyaqx9losU1tLPIE0oo8k8zFqKOz+sDU3ED4VaD9gQfqO1jR1i5rq
1uU71opelx7L7NJGkQMDPZkUYdha65sW0LuvSVSjMYTaGpG+cunYXiLuc0ydF5bl
6mw5bUGqOyaoHeLLEH3UUUenqf6y9Me0BFqb5rVDHbWCXAbAJTBanhIHXSB0kpHd
xIhs7VXDcHEpwiHUtZALKBfV6mefBN6dUAJIDjcAFrljC/XEmNX04xX83q6QvZZv
T0/2HkXi3s4Fe/nUkgBu5S3lw7P6vGFjQWosXRGiKBOh9icyfNCu+2thLybYhW32
BCTTxKbW+B21wTsg/4MWSbR0jdA4Ar6bz8ZhJfLbgSMekBVoElbHLJOsrfNkqerU
JDNq/g9tQuz5S2TE3VgSW5TyWrTA17hjXRNUOWae77y3SykT/SYovQA+wlO22B4f
a1P4clMBzCVWmFI4wTjuoy0fgqxDyIdKMu+VIBk2i6Tm+FaaPLUq8AHU8MuTJkfk
UracKyQtZA9EeKhHvPRSbeUrXN9oSg1v85U+e6vZfBTH+ROdDKmoJkXFZUieCII/
DCF5/iijU4B9jzbBfEsN0iQuuz8IlgBw08jVNkCcszX8DvZYWfie5n2UTiv0vVoW
cYfNjrXjI6AExHp86BHloeRhmR/48G0f7dSgNv7DXbHFmdJaS/G+nrDzCj/o25nw
Pq/WQksN9//ekt4pH/AgFjGj+kdYg/tVkWXb1h94ZsJW3pHS+rlRbHpqOEyzkt8R
WU9oFP+P4Pe05d5N3VzJDZzlYLxAkcRnsHZl5RcZGU0ZtnSMJ1j5WXOBfT4kUddc
7J9zi3tO6rymLDfv4cHLQiJS/5UR3aDKF9b318x33S7PfmkFREH7nOh0IuJrehea
NSCirol6gWXOHt5Mit+jIfZtGepz6rVsk/wLjtlhKtrzV2Lmq5Ix2YBCUs8uShgl
yj9CuFN8gzoKeSIWLnDe3VB60qUqnT/mnk8crJB3PPmbWDtjuSljs5kAcjbqVb/k
2ZZ5WPE28Q77wNbrxkMXfZoQMvAngIJSNNK3xHGl7kgsLIfIVpzAgoqvThbNB2O0
RR2icgkSapRLPzJ+RHF0w1utaltQhFTOF5J3sBAnTtju3RDiuBnEKRn2PeAUq35h
UHuftN2EcWGAO2PIHAUvWFHs1lfBU1/T3l4HlaNOaiFLf/e/Wi4Dg4WsRWIpEw2M
NVfMoAw/Wn+go/k65akvuS1FQc5TysuM4GqJERnq7d60jLsWD8qR3nSev4bJgx3H
/5DbxFUS2yIIEkyIz1VTNLPG0OR1zr7c2E4+/DxCtl9TqunUArJ86i3xr8/sSMl/
mVZSlULcOhwt1QHjz04o/JjOD94/1p8FM2+XZCrJHKNbwtkieojx6cYyn1d4ay/O
l7vgsnZacyk4lhLKr/K5763HstxqDRG2WTMEdzMHkIFxmu5QaSSxBaqqr+1LC6iw
IYzMzISoLVVxGSGPsTyNFiLzPmiZQLmJZh0BJP5zLBBsWs4HUPN8Dq8riekaBLVK
/x4BhQm0g7KeEH6PJwhoJVrwx+ut9zM70QsHGf43bgcXq1fHPsYBhMXyoQyf9f6u
A3ExIFq7L5sIDHvlUOALNCMw/xFXh9HK0+bja94HApFWF1tiQfzyqBu6e2xV8RRk
Oqi04kyC+H61QX0FUPz9HdsIoerlpqtfhI/cgqTiPvrI1/I58BJnOUorS2lT/bU1
BRVxv1H81FObgYBXMUzdM5u6SoLcQNwrFw3q/VWDz1Q3Be6kttz9l/dfVXx8Fftv
7VUTQw4/A1qDBYRg/tJDVZ0GS328onpFY56NZXrB5WqvHBuSj/m4dqyOSQuImWwF
aHiz+/F6y28rpR//5QDXuYylhvhD56YqpmXt64ZfttHw11uA2RukX/6FG84M71fU
wMqHVGj+H9LJwiqGMRBW7SYj7G+E4MCySPNc+kLnOA4wN6UqbrZl7kbhTd0mgZkr
vvHh+GleALr8kam5In2bTxSNVki7xlEQA/c0m20Zh9Qg+3Xg6W9tYBAe6zNAsubL
71RmrDrWpoEFh2u2mdpa4KFTGQEvMAmHG75BEavory0qqDQt6VJRPfQk7I9ikHP7
S40gSRkbsuBPI5+PVbouF8bG4XNAv3Z9lbKEWdX/UgzLd798Z4jLAWDJ00l/o05v
dBIWvsBTMEiAdLWElx9JnrtbyUczwgRA2dmP+gyf0nAhlJqGap4NUBrkMdCVwky2
T2LNRWUq177FD2/GGNfCQ11FfU4f7MUi7UfCVEjkuxi/Kr5dEms9roy3IagzioDx
rPQkky4rRFOSvBweKXUgpRemW0+MefvkSWh8g3+hh+WPtDKeBnN59wUnufGn+VXX
8aKgdg8rqa5rrPyLGhfDIcHpnFaj/XGngu9PtO1zPv14uMi2u4KAlMsEg05PAKeC
LV0ai/r2qcF4kZUfFF7VqJDWs5OKLf5H+uhFF8gq/Ojgl/7FczbU+jioceGPgcLx
QRCRaRQfCo6PARMoPZmezF4oGn1IyToEqc8xERjMe6bzkl2GFmaWKQc+Zr4qxues
7SdLYr7plN0Hzzcl2XKx1Uhy7iDE2CmT1DRkingFc1rHJ7jsfA6fKJSqUHI8RICF
xJOTTxdctu4pHxMKDTOsbUWoUZiLoZmkCKroFCiY3PzQ6hlkPkwqDyku3SvtGiMr
rgOYzdcYby3Tq1hiayO/U7cX7f9SIDiJGQLgy/36p/wyE+7v1zkzEzY/OZ0zxpLT
/gSkm9pK9bjSAn6ydhDwx4cBTYnOpoCS2+lwC64eDUd/nHRUUD77hBJqStaPJX5K
yCc8WRH+Lvkb9XY4sq8okooa2aJZnswpxV4aId4HqQkS5H/ER6kRSuWcRLB674ce
WZCXIWJgi08Uu4tn49qrB7dSnu2tf5459U5YS4Av5+RAVA2z8E3O3IMEdH8YD3jz
JxqqoaNE63ywSD4xkj0hnme/yq5sJsZ1TtyS5IrHqXxWLdul1INvG4jhOdFQUKkf
JIeECkce7OFNK3ZDIA3D4iaqDGHRwyV7rcS66ES5NKKKoMas0D9PEz2KajCaACSi
GtI25X+gdz6JGFrdyeEEUlhiHblR4Yfv/WmxoXYS43U44NutIUKPbGo8RD3iSNHw
BCaApHdvxZ5djYEZklwxwBxcbNutx8EZq/JK+vBmZbIUZ5g91I+apQ4g7Q+O4w4x
jJ3OSWgr+mrRr77wTynjbbyqRIgUupjkQFmzlZE9e7DAPHQ2AyKdEe/1nja4Nuew
ZpU5dBfWGjKgfbIN69eyqSWRLZwWkSB5PoRrWxQ4qXDzxXf0+SeNdXCBIhrXIy/D
pUHa527fueGMBJvP21BLAs3HjaO7Fhab5Uy305XW2wyHXBel5XaKiTpAwmETYTop
BdMHxS0zbXpZe/ypxuzZqmsIpPMzJbrYZrlYc/FSQmH5hImGnVSvaenuD6XsIKqe
3gV1i6RaVPz2pkhZN/QSqs/Q+ia5gbbZVx7hL6YqVknvimBx446IVqyywYvpVIHS
tDJUSysw7YuUcttBm9umiLxh5OZCqjnj31fAp1eqPfC0nCswDqILS5LZKLyzPxvf
IsA10DqLZ7NeaIUeSGp4wUgF5EtKirwL8AdIisuY71VPsthqdA5wHIsD8lKNn4mB
Z4lRm+V+C8PVRZOgRbxH6W6rqE9ifd9qM5252AUgSfWct3WDyFew2cyp90PYuTnA
zlMGVl5iiFJWzalyZXGQ883mSkRMMkJ7Em/Im5YW8w2lTpsstpNSS5vcgJ+S8EQ0
GGontgOcBFMlUgLKPlCIKBzXx/Ri1lPmm3G9zG79omh+1TJhYq/Wo/32lu5AXaiH
/AiwcvUUJlkbmi60ZXia/ljAHeIn6EZgx8qL80y9nHt5JfWakB2RQi2WGrmbHKUj
3XFg3Rrx3dPwUTyKeKIlVFZvcyLojK0rxHGp+yZPhITn/IvD4ZC/yhIB7P463RlU
dD4zUZVpZmRVHd9HnVAtoyNmfFM4bk0lv2f0xuCSfgsjTXMemxJqu7df6p9dgRx2
wz//ZCiAdP2uuG4hIstMbjabDU9FpdQERduRlT6mIcxXSIr8bqHRh4URDBUWlupN
jT7sfTTQiNpWvMCOjUam2zblpnwo4rbBIwjaq/mJxnivzpU+xe7ONVZtRHyEkAOo
GJBTnhiH/IZE2PLSmnjpnYvdgmDQk2xWNZPl8F36OMF+r4o3NtSIUh/ZUBzcG5Om
zxP3OTnkwjxPj82Lk3SrvD3jBNbcRvYJpk/XaD9LS0F551uXSrp+q/Ofh2MYNKgu
fcAHd5drM1+NEhEqDoSS12+8Ze5TM7gjuIJN86Z4i/cFOEnauJBOr59Qj3w9iNbc
CWbQ2qxjidyapkN/VLxgWQnAhUd25aWcJukDS4V2i3r3dp5+uFOIpK76AnWqzC6u
vUGwd6/YxVjX2x0Tl+8cjq8NYV62L7rRitZNXThJ9W7D0pSV3PXDxta9ncKIZohN
zaGE2VYnMCiGBpGzzhxB/6MZ65nZfkS7WYxfAyIfNDP6OgBb7K99GkkEuJ0vup2F
eSWfFqLBbtc1/uGlqYxquHcjqFaktZABxnvyoLQnIH//kXZGNbcwnPxmWd0kEnP2
aiEa1U7EZoPj37WwAiK1mwAndIjzDnce5bkPIICepcn47oNgz7x5fIv7bBbd9V7E
2KaUueSg9eBdNZM/R27DkyVQ5G8ILnbFSFjFLAtGakoMWgSa6Z4zAd4x3vkJTm0C
hrEz54eUy7rqmVfcrpKr2e643Wb1WODVkTraBno5Tb2F09jZeq9Ohw2Jxk5RYLSf
pT4m6PKwwCkuB032uE6QB9EK+06+T9StuCdNuL2XpwFgsWw95ZWaibwJCwIH1m9E
WdBUGB5rOrT5JBxu3gKZisLvxjOshVHK+R1KiAL7kANO4l3oNXIfE1jSR9HDwJhO
o2QapnArxDCLKBf0+WhqR3mYbMFYRHDU4W/w4t3XiTNbSWtT8/r0vTkbFl5/0M2k
UX+/wjNXfuAlnBsnDZqoJrVQobsXtukBBxE+6NTN/9b8bmZJI5XSgngnAGtddKuO
8JpyVaQejaZh4iMBmBS75+YW9H9CXvypjYDgThAm3/K8f1aHThy/2RGugqU4TBMa
TwhZiA0/mIYO05In3p5zLd9k9o/zb9QKLQWNL2p/tFzEUT4okPOqywahZk/rmce6
eC61M5PHGP6yRwvdb8wLjxDO+HCmCtRfbhPA+Va/IiHPDKhHp0ITslvMVyHLEW4A
teHiRoy32APvtPsXA2EqBp+Y6/mPgqnMK/sstys/od3XLO+0jhOGTqxRmqqiTNby
R/iIFOLs7aXVSobjowiyJS5FqfrT9woTV91fAuDbQY1QIIPpniFuS0RrIbkaz6MV
FHjcS+7YqQkGBACnTPTCQgqC2msZ3fTSnu0rPrrj8juIb9tSbtmD/bpBA85a3rQT
6+9iWPuTKtyeL6YoqF9erOVZpvccwf/ApUsRKLEtd2ylOfJRT7/cNJHYyaVgzLC1
BDFRyCrwxEXpnqQIhLB8idC4T28gcC9cwxo5AhDpynLITz4+8RE8hBmA5plgraX2
/PjHkbKJX+M6QA1J38o/CliPpJ7CK5xkJsJoZxRP6HvLJt1c5wKbB7UiyqPMWdl6
ORuRcOsVxTIiaBy3YsDoZphc7Ockes05vAWtDFct02QprKUWh6MjHcXcOvsbB/W1
ib2Ikz7cwEZgLuURdLjUjAVuwfws1+7fMCSFgPNzO9TTe9Q8jfAGDDW/8xpvy37S
QQl17qIvFcaJnKA04LLmSlHHUulC7l6lZz3pAIARqAIG7iYdQ46j0nUtbpviCHL+
6TQxSiyjX0j+nUaVfElNC5+MwSprFv0fiRuxe0oJ5mI4UH8PuQFCpFxLicTuqL6A
KFF/2h5CMPMCdkdGkAMQtK6JfqUTC+p9dTlshD0wd0CrYiJ8eUKcJKpjdcnczgbx
O02aLFrdjnlToKe7EV90rY7cgZVqGGvhBxj+3t+3AZpoxtV7Hphh+hzkLyfzPaj+
mx99sYvUlDwqr0jRdDzner3OVSOXXWu3p+1TEz/HlrAbtPU+ozmD9+fpIli5zewW
XaEkJG7o+/SOSa4Af0JQxLvbY7KprwuOjP+s3Zwd0QP/nnvt8WROoJpNoUaKnnSt
08AdM0XPly01VAFUQGy32RcOp9bYRouAL5Ov2apdVCKAnW44a5gnvcQMTHL74hop
n1J6jBkqAE4BNRH5C0xV9iqcB/vWopvRI9OCTZlv1hwWtoV6QeWgi7S/aHBilGt/
Js46eN41+Gu/yhVZuzR76HS7daIYCRjMc8ljf0AikG6F+NEhEt09HcIO2PLtP4uP
lhA+zt8x+T+OSvopKjYXKXu81bdUoCqn0yp9GGQk7udFIx0o/UOiu06btDgPzC54
N4q8FsKJP7hAdU9T6WHCbzJOmeS8RN6lNegb83zPjBiucmYHt7OaVpfc/h88Jx1d
+0fG3SFEtqa8b+c5OntUsw5kxOjF32VHNm58BDDk6mrSVpfSAhAGEGcjFdpV2wTp
ASIbptTJ78MGfpmNh/yoduQwaw0dMPajRdO4STJ4QSxh5dfxfGyVGWSRLaIjK9bF
EJXIo5jnaMhsOMApd/KuwGRs3gbVyaReWd9MjrJ4N0IoKoQyYx7aTRdRVgQ+qB5k
MC/sXeZzzApP01BKDo9JUzamNVZEkiBtWlAISltodRtG3dRR2QAdRm/MFVYPz0Uj
tB/49UrqS6SjqdxxI1ivb8/quit7uUeUWQ3iXtJjBBEsU1DbKM8X3UMs47zrAQ8f
8G4cBTFu/y/2EN4yl5KqbAkxZv2EfBfOMiXN8XM0sqRwDlJwP6V5y/uoSfvR46DU
X5hoE0Z1mXAmj/bD3RVacrQt0YdDtQ8aPGLdXTgT5h8BAh25Rs4EtRboR0lOirHv
qWi9/ixCrO5oWSPGMkrA1PDTJIaILBVCX0VSvyDZM5+kUVEtNkwaucghaspUTD2W
ejY5oO4h3ekaeAYngBDPk+rD7IZ9KT+SrGwiIFQe4yWCPXg4Y/MccIFi3W086KtH
61wdTvfa908BpsjX6pXrT0unCKWvRW+hzJGt3OgsvRtutS+/hedsSsWc/mWI5ult
JQjqS+Q3ZDxWLfq/TSbo5mTrYbAfSN8klTW76CwD//CAsH7Ge30pjFHMsx1fxIcL
wZKr+YfvW5wDwT3dUg7sc/MrhFcsR4Uw+4mxMwH9E8ZRuPj0J0dCPQjnXLHSkS0W
v7u6gamQsTS4lAzkfp7VLq4tbcHcze2/gg5p/18bBGZ31SeZ14AlxkW0gwq+du7C
qJihKEeGToSFEDHRSOHFEmWGPMiKD7lw/m3pgAwZL5kZKJQvvA0XoQrXzw7YuqxQ
8GKqw3H3cQiN9dab2kh6PFo3DySkFRGbwSyevSO8CSapsu/LLpgJ6AtfEjsQs3G4
rGM0i/0HWGo7IG4qGbfwEigeCS/CxHWYwnM1c4B0l7I9N1boTEL+0mIXOANghFbr
XqD18x4iEDRZK2K5yahFExDY/zdoiFl4jDX4N1io1xU3OaZDYSu9d9UefK3cDSPD
wBUs+3ZGIuLN8hD/h3OmrWwzOwipfE1XHkgK1Z0toeCEeu4InUWkeFqsd7XhyrBf
7nBuSG+/QclnnkmzCu1xAw8egRd1YEKfN6cnz687AiMA5BNf6clRqW/rXFb52xOd
iqPngtM0K/sj547bYF3nEN5EziKTHFRAy3/kzmffzmcXJ4h+b5et/KAKWgV3C/kx
+dipD6zN0vfSjN0hz7xagy9RECrj6tGZRTXsyD1TBDoRAjMl9LpE4HT0omSdsoWp
Q4rzI1WdpgBmiC3slcSrFmg5nGIrx8r1+oCTsKFQxmvrvwTSQsYnDzrqboWB44PN
aWu2k4sMJgDAHNa6PQQHBLrrDSevvv3GhwUlOUORtiYLpINj8QBKLD6aMZ0H0slB
5VtTV/txG1xt3ExtQzxpOl4ww4TPaGZS/hFDEtu+Tw9EBWSL8bC0798RpxY9rWhD
gaYQOX3UlwXHSUTvebTDxAGhCySR7BczSDJGLDTihODNbjuK62OFjpIeaBec/Had
C5LTcGMQOfjKZM2b4Cb5crqCQQGMMIyyQTGBHlDOkKo3Qt9hRFkYT/zWnGasCJ5I
gFL5bplKAHmkFBHohBuBJbarMIxKtGRS4AR8ZIeEZu/z7RwjHNkfIt9YuJoAfdc+
xhQH/JDWTZfgcosmkPAepl5DynEGu9xrbDNraTvK5vE0zmm2ItMdCr0zy9Gzj8AI
j+N1dGSUur39t/ZmS2IPe2sWV/w9+CXKve0l9m3T2x98o5AbJX+7usYdm552hap6
D9AR9Gkw0KBH/Y3TvvHXq3m306nlp9LuJuL7FO27d5GGoq/cUhKw3kZSUB9V2FU2
gERZG0Os+Zsk/EGBaL4WllM8eW7t8bGt4jze99x0h3wbWmd9gKzwl57hNHeVkbwx
JCDVKorDeP4HwoYcWcKkUKJTSE+vdF9Ol+hIlFB/3HWxeDuX74LECCdlWAy+qstj
4I/edno/tFKYVzxQ/PEIsIpYTVTsEZbiFKzs3G696tF7Mtgpo0c1YdSE98v2zgSf
fg7frYQrwhu+Jju1z7A7ggTytsYZY2CqOln4JS5/3eRFN3paV1Nmz2arH6G0JMk8
O2bsKuJnUCixapBZcS9YZgQAtDYqFxaRo6FhdMTAn/mGo2VhJPqQINAyxgyyc0kW
HWxTGIBVNyyHAQaC1eQlSvpW8TCfUST83BJIGKFH0pbu0st/vreCe0mDV0SKnz95
1/JFO/X0ZrbZ/j+bHjqIIt8NU6ug1DKzwEOu0i+6xiGtjUI6KveincwbhlwN0XDV
JQB4Ze/U0BQ7MnIb0sRt3Oz4NKwGapzx+PMlZJCOMZNGL0d2ZJMFBwSSoVm6gsRy
NYjU7Pq9anla06qGc8GqQreeqGB/NdxH18hqY7tAHk63iCEyIzlcZYYcRqqrA3nX
q38rwWZqe1x4USIrXwjGr4Faxxc/uQh03cvvG/MYVS2jVscbHtGA8cxHu9nLuf5i
A0tvlAo94k+e8YgaAEH/tE2K/ImdzTfwWWBJitKsNz0pDDc6RN9Ws2srnNF2vIl8
DTm1WnEYM/tPVMvVpdNRbg11eKyLV07LpUcjx6gBW5xuuLfF7slvVL1dYx8yp0CU
bKkOAdDCGqxotApiNQVNl11y0Bjtu1ztPGOM2hVW7+I8C29Ng75TrEgHjnUij/aF
VwzrSr9lpG1kLrb7LXfSoY77n/i6gcEy5t+JXXmpW3ATRxwg3gKJCB8y9ELWcyCH
9MaVD3tKKuK7W5azpRT1rvGZw2Odchqk81xugkV7v9uzuYFXqhw/7VTTZS/CGJ4r
PSpiektulg8KAbVw1Khi5DR0zQPNswh5lGmtiWoYl7ng+0twTja0/16FrFH+JkFm
Jc9aXR8LO6UiU/Ii6q4v4D9ztj0ZRegPRYxtaN6Y7o5528TQTIPfzsVevvaYrCok
m45K9ChnoFokieZMCnx3/57Tut93ide+svyso3hCvwPH3cCO65IeYrZEZU6Ee5N2
/jd31ZpwSiZXkw4HsXTgBb+IVfcXPxlsjZ0zdW5fOnT0B+sq0QAstPpKyzxlu3Y7
MkYhxSCDpkv3Pn2T+sC357CFO15yNJjyV5Fkua4fosdF2gA1Ri9o9cVOKC6GpGFN
ehG/UhJAWyYLmpj2abeFWLWAevP26NGr1QKxidA1unDD2aTRt5rAnNW35S3klNoi
mT6731qj/EfTuRik/PlWY8JxDrngDs5rCYCBIia+moHyY5yQWOkhxOUs5qcvCRbP
dsKwT89pILScWDtJV1YWcl4EXtWv0+4poCTuXVXsfUbTcBmWXw9qyDy/jLTn6ijP
1Cm7CLrdMHtqarLR1KzmVpZzMINlI7tDC/nQ13PfNwohKG9XtYPgcMM5LkMqKlx8
bsZeVpJaFf1hbXhK0qbynLZ/bHumRmM46WxMiIt1/WkgPnWaqlQ+Zyg8EGYi/YB7
zDDhOrUBJXslsI7FLlfWWQ6Fs7cIO8r23aDsYocfsXd4AqR8A2L4M2Vx5HnF7dxQ
c4m4+LJ6DCKgO0dCBJAPcnnGe3uSdkZqWqZzdA64X3AbVGrZ2vJ64LkIIYUL6G+u
beN3MkjlBu9pOkighJRtbHaceI/EXW4h1bs/bm4N6GQINwh9K8q6T4QrXup6l2pt
bS6/F3QyRxjc+H/62e61FC6fny4oWRFTSxzR3rIfdJl+eD56wi7RyoIfQTzUV/z0
o2WUlRbZIv1Wxs6rw+s35VphnTv73xkb+BsyKeBoz6ecjA+tYsCEmyyS40B5Y55/
Z+X392xCZYkK4pizCXNzE7CATOJgE9cCT+5qQ8h7tGsLjGCBemiNrC2cpjFfjecd
nz1t6/xY8/nFU3erNtq7sgzG5ofRz/SOjyiFBARVjKwtCmzKioC/DSdU6Uru99iB
oTlBybwuQLbZprgib2YujRYuaCoGD+s0x454Llz1BIhDf4EEKvQJY3rYxhBaiF5L
MQN5wU7lsmZQKrcqcm2J4SRBhOWcnaclD8JnNB05W30hh3zmUYn0LPOEvDooc0pa
MQ+867Jp3ikHafHDkJTjHhw5H61WZ+0LYUc/1DSby5UOrqeo6ZkbgjZSlu6sSXca
mRvhHxdwpCglfcWGc2TzjKhcoT2NqEReoxDqY/lLPrlvxLG/OQ75oG8qbIvp2NNm
Uogv9vhV7BD9F+oC2dFp4mgna/Dr/+6ud36nJRk7aueL+72U10fVWp0VHezutL1N
K76LhQ9ULQ9STsskbZnID/0+GInseh5BsFkDAGQZxjF/sJOVgnlq0QOIFZkik5Lo
XJFMRqQEIiGQMhqN5o7jzpoSMohusZZ/3kNAtjdhwdMLujWTId3Ws5U90WZKhgDB
ZAYf84gMQQDigqlaW5xnMzjU58YmFnOz6S+LeLUcnO4C0XmKChNZfWrMxhXTT3gI
iiU8T2HF7gsrokCjZmqaZhq4z5fAwotQZFIJ8WToy63Kh3sGiBHwmBWn990jfnhr
WgUmjJlGAjnB8vcPRRW0myYq7R02fBzOjLAroq02Yj9niV/VkvEyE3loIMtHLAxE
D3wW1TTanZcRYwCLOhMD+wpwLUobmX7QxG9iTr3WazWpt2I32+1cwP8pUjsBcuub
8nWNrVHw4WYIWthmBmBAUDvza//nOutJrDivpitStk99nCNPyddeBybGQ9pybf1x
RrJM8dn5HjL8Ik1vw0Hk3yEE6TL+5Z6ugW424HWhzUY/i7/R6KGFCBDxu6gtxMvy
IXostvdjuNAcv5CwJ8EOC0XD7qMxM/tFk60S9yV/Ksuw1zvmmpRpgFulelOF7fiy
EVaAY7Og1yvyXRZO6IGgisVwQvr6hNcgcbwd/0jNZnx18K/7NAy1wqPOG4reowGn
tB5dttp+i58CyneLnO9/6lVg9c8Y2hrdDr/Fl0OI92YoBNeNBLYKhfXZXB1SyuVJ
OiMRkD/vsyH8g1JFMxy+DeSd0zu3NvWBpA0KPamvSRBlOYsRYBowFXXoMZsA+uVx
P7mg3bAgcglQBLVIF53mYiyR2Y2p/wkOaPdp1vp78cGpX83mSDt+9odWjQK9F04R
28rbsOwSwGyom7bpwMnKmEsNGdZLTL5wFgtLNHg6hYxJrWQKyo7RaSN1Wbn43ZWk
1azTlf+7FN0FvLmBJHU0jJhTuk6NZ57Qo8y1XePOH86ZVQzXG1R4wIokhFNRfnmZ
rrAmp4FJtRW4hbrA+IYRHWGNiLH8GQj07+hBw1MhrUAUsJKO5ixGPg/8SUfQA9KQ
BMKeV2j8tbUxx8gT9uv0ZgneIur3iRP3pB0sGh59Xh6SH4d/Z44+VmZRlRtfHBIP
kx5ZrjkbXPzu4aCG/7uDuzZLNJsaXHx/oJS3xLoAu+NjZnKrAqkZsJ/UdkAOQhi6
wCxKNNSN7C9DIU6umA7/yQCDg7kRjEYfVulIaHuTnQR26uedkVObIsUuwr16COye
rwrauX/d9VBHD4mj+1gQySOk73qxPG/5FswmJTZoLDkVFzYHRkYKOs305wO7Goub
dJEiUDpVXKnmt5EcaHnxYpEC/uhDpeBz3MHJWZyvPiS/UuLLhu4Y4e6ySY8J15ic
MWnAytdy8CDrw/W5Hlgkhya+ozL6pdPpn3hsGKTGfru7iGZSiWKF9G6oD+ghppkw
huvia6Zo6hXRnSJ+zcpEVl3do21erSkzFTJtg80JSEaXiBnflkhgY3l0tXuGS8uW
d+EcFWf0O017ta+Irg3shYgpcK4ujfmFu52hZcFua7Yxsdl3Se68KAd9a1+TaCaN
juJtmp+3s+ZexacS13mKvYaFqz1VRzm0Jv8cT8RE09YGUpqTQp/03QzTh9vWNjWK
E+i+BrsbnIFeGaZ/Fq2BBMjJ8rpvROBKOJ56v1aD3y0I1ouwg38xmNU6Lqui/r8i
7eR9kyInSAii7QiQaUa+bO/pfEAiROanqQ8fI5PiT5HmJXtZC9X/w/8Jqn8EpwE+
f+HGFL5zRNGSNYC/zHXrl9KuVV1Q9tj47wYrbSVs0/iZCiwlRWNE8YLfA66uUHl0
PcNS+ewUzpZBGUPpkL0Tlt2knWHa5SnYEWkbOZCBPv+1uUWTqBNlMtqeXukC2usN
GB87fx+kY4gJ6Mqx24yOJ54xEzr0t5Mveaik7ALYO+ZzG5VWxbf0aardGtCW0JTX
5JYWRm2+Q/+2aWxQq18iO+PbnMMgKnPPREawIsHY8Ah7QTHPfidUrMk+uD1GMaez
fuD64v4uBvKbvdJASv9B3AawpGkKAbp+01Bve/amDObsx6tJWrGXgsm9ulcT16kr
E9RcVdUPu88jlmu4M09C6HIlAsMISaz/3ocLU+kQiLlHUkIHKu8BY4gjYMJ24RbE
NKtjE2P7a5PNYjC5A/83uFTangRXt6MMJQVbvDxGM25hA3SzWmA62Fu3HFJTIoEb
fIoQVfn3Cn3QfXRl08n7HbEKtGFUTLMBmuDU0ryg+5kKedETHr/rej7lnKrEE4ZW
g1XLkGI+ygijNIiuIOwQ/sdVVCejo77RF9UNxfmL4kwzDpkYSNc9WFjEYcEMtCzs
bFNwkJMbRs2SJ9vPl75PENJ7oEhWts9ZXacq4PgFhmxZokf2vBb8nsk6PosQEj2E
vtyVh/qYc59u/sLfQQy4A7MQ3F09e4CTbtuOpbmNfJssS4WX6jzX5diiZ5ijR3Fq
URVZ7/YkKsYyfhUAYbzHla2ptjmJfIABV9NXuKTtyu8K5g0YF+hz9pE26ZqfU+2e
uxDycduQeynBI801AF9eosq3hCM5sq21saWKrt/tkEVHccU/f/TVjp4W7uh7Kt5m
uucN/Wp2ex+ju89ICR8OFR32Ju4mfocDNHYtz+C9jxu9MsLTNM7f+2zUAuct26KT
DI9F4G9IurwwF9GKuSPOJW/LzwwyIs9TMX464tlOFxoEdZsTFDtGCaCt2gR14P/Y
HykMQnUZ7BRzHK273Y9E4DXWJK7t3sawP11yk5d/BRvBfp91x7qSbYz9R5jbEPKO
Gz84ZF89yh6nQhBKtocOMnvhsQZcgzdG4aGdypYQ2EqxTdo4+NN2eeFp3NV8K4ki
HdIQT65ZiFxVT1rovjkMrPWyNEz0D0+JS+metem5EDXQXd1cT44WlhY8a87QbaIi
upgaQUF9OdwSV2TwQ6MiKz0RldyO4g8tgqvWKweGWfGZnKWf1MscJUuG7nMTOD76
w1K3fso9x7lEoSnNOCX6PK979/xiJXAKH9PGBC+pDt5/p2sfpdgmsrOJaNDUM+ci
Ktep5tM+4BGTXo8Z7D/ib6wOqt3uEc0Gc7kaMi46CzZkf2Jys6ThMG506rmTlEoP
UGMyK6vKl1fnKOZQ5q24LXnalP5QGOjLaMH70kR4X3LoYf+cLZd98bztbfz7K4EX
TEcseto5HylLbaBJMl7Pvo6hkoJEz/pyaog2dPXZdF976+pGtFX2isK830riyo+0
86ZmgumcEKnVX0r7cnGm4RtMcTvzwokLTsdOcv3GIyXSz9tKKaDOfKiL9/oncqYa
MiaM7lYoOKubISQE7hO0mNThlAN4Nxpqhzs7r+Iq66bB2Fv3it3bSFemSHVQNVYY
2Cygo5ZZ/mZ3QE3IXcNp0AUshkvnuH2y6Wy270zRidhuhELHQMVwNBnQ23h1zxt/
SqaAvqjWbJkPDbvs6wxpHkRYdbY3fRFOajEszaMzIZ65p77a+dPR5y8xN6hWZX3z
XxkBI0lfFKCyfOnPFibrBCx9r6b8wPzOIGlCWe+Ua05lDT6sCyRPKB7VnSKpy0Rj
REQD1VsZSvmwt54HN1z1ryn6a9KEkYEZpCAT4Fb2fg7PUsnlWUWw9SgduGccOsH3
g+qX7SCJcgGJLN+LmifII2pbCjCkbCtGD/cGkv9xdtT/YtvnIv9aBJXCB6rJzsA8
h347JQDw6bX4DAfK0kqhMgsG31mJXwHGv++rV/zFg13d3GTzimKzzt2PWoWm53wO
hqEsX/ihrPwWxd1Muj4l8rwIaFGm2Tw26wHN+DEhRPehRZsjimeQ9xJcPL3nSDX9
gVeF0ZkdGaDMkE07MgVF7XkItnzwY142le5teZO4pxPQhO38mOBzgd6VmbvJWK6D
MWqa0KgTPoZPZ3QivvuMGis03XrLiSDSBpLl+aUuCAzhqhHFqrs5V+CnAZZN/cmx
Fb82YfRenwl3i2oVJLfViJHgi1YW8Qwn3ZGMG07T+0kHvkgbhUcsijp+wHRgOII3
WQrHCVA90ay0RsWMueq6YBNhBa+TlI6/75L144qkuVjTUCJYpkWJR4VJ0c4qRGV2
F5rSvsiWXPoEexjTKGvaigEOZRIi0tSGCodo86IH8oBS353XhySJmaypEUp+L+/+
2U4sItaa2h1a1u08yOJTXwpUMLimDA9LxV4wpTdAHv72tpRW8AziylKTRs/qVJCy
9E38MkI0MH2BB0CvxVVS+n7xoVi2ERAv0ovKxd6kK+HyR6fi1d3LgrG0qoZFGQ1r
fP9byQBTdyBzDORU/ecnxTrY+GMys+HSz38Q+MLYHXv7611CerGJF8uv3yHPAT7h
TMLyRD9pzX+tJ5yKsoi289k3h+m0dkBlQPS2WOPOsbRdQYAQHUnBc1p6jIQvcnFE
TgC/IuIlldpmhf1EgcgdVwhD5RZDDlPUkuI9Yn1QmCT+k7KAT1UWhbCDF75peGqr
0B46sX4jhyFT/lfY7Ym/e3oGHOj+oQA6CSJyIJd3mm26WHjZtTpuCoMuVx84069D
cLZnUaZH+QoW6rfJFT1YqVHwlbduHSqujYq9yHVr1AmimRldVoNuDo2fPDkCI/GS
ejpZM7/wGi+unbTQtJHGOWy3fQT/HzhKAy6lxrjXb3zjBFqNRygFCyoojjxxnDjI
TdFRWVfBSi6nOVxC+unSW+Q1IzX3ftbzsQ7l+plZKpJu6xuTHrdZVxtYKKBf+ego
xl/o7HdGzBqeJgryqjKoSdGKj7Es/4e+j8chGcJd0b/6R2mta3kYrWw6IGUr5wlF
A05imQyFMWTYLWt9jsbA8BkO/GiDBlpDm0B7GvyVd2+K/p7zP8M/akzQ+bTotfhb
fgwrAlLKXHka7ERMNMl8R0U+e2coI8IBXyG2ElOyeO3ftqCfVWjVy7zv9R9iH4Kx
QaDdoeeo8dwxopNR2Zx0Nup12Q46HaUmPwIknSQbRiFlEx4D7Btdt/BoGasTiQqG
pvIQznPceboxuxBw+OGP5Q26w81ifQa8JNs5i8cmefpRBtNqbyTZ1H4pf1FpOgT2
jrZSKOwKof6wLKFE16xP/QAOtxU4rSbsd/zMEftUheosVcURvIrvtRRvij1KPX7z
/xu+J7oGwLbMOPa1/XRrB+aqD4Ptxncq3meT+jO4kwFh4aQR3qqHgKpBnOrq7Eul
rOddQwAchydvZEsSimzaK9HzzbVcjreP7dv9DlQurNw3pNDWiRQFo4Mf+zWyWhv7
JllDDpOyo8fK/2qffh3LLBr0jqOVgIoJs4OfC9pqP+5Gsdibb5h/5hsSUnavPxfK
SBwM2mbVfXGZ6KvD7YxCI2oCysnhbyir6x7v+OQ1yBzVh0Y3T3xgmymq6RW8KUCK
PQ4tl3/BXLJtd3rwPoMPHZoo0P2rMKNmXF2Bz4RpOrCD/w6MtGlTw/SCBd9eEsmc
yHVj0Vj1xHYlrDnKr43jjgEL0KlfEg8Ai0OpnnwcfYPZadPVStozy77TgfVdhhCC
74jOvua1gdWLNf7E7m8eSZ2GQyIfn22ntQYqZOJzLJePzMaYRx1cBLxd/8+l7w4b
xCoEMNtwb9e83T+lhehWB1iST8F1h1Y/WbIfgX30I4Q9avZ+3C+aD5tekb86F1dT
sfjnMRVdPL8bJo5ymwe8mchlQES+/BxNvb3C/BlF4g6eYnAj5BgYMjVANUPmwKRM
gL7ZKaQB5DMd8eBWRrM8ojofO5eXCAx6tO01i5OCcNP5PKyAruTvbo0UOT98sITT
whJ4PJzDGr9pL+kWaBffE2al0qPxi0eOj2VxVVDSzd+hx2m/lf06UbdpiyRQcFYQ
+UyjNA7YdfBYkd0MgRKktI3uQSiQsq+m4F15FRGYO85GG7T1xN5WUGgd7upwPzys
MtThRpTS0aLhmjaU6fJHs1d/iReuBXdJsp79PFlN2QwJ2bmQ/89U/DpajXH9O6EU
7nN6d6Nn1TAjpAohMb13H57T4J5XDRMjg3bIO/AaJxIEUav7WPQt5bgWOZbidW9F
OAzJv643uQ9mDAObnUqBcbpSS++STeJ2OmrPWSJ26V8r5+g7tXMQcc6wVk+vHN6j
0uSXG0qbPKe04A/lPRo5zHn5WGMv0OZfbYnY8fiReEE/GAJsFVhOMAgZzrYqFdaa
9m0+DidQ9bE8qtm6u88ixy+TKQ8U6EXGtxwOa5sb8zHuiIf9f8PHW7ezG76IQrVd
GyaLPtCFHeV6+aIY2S49E31l9Vf/TVe89pXhPM9lq8nYajtaCSsgGgB+NlbAD00e
qTdhA9JZHkTiUQuo4WQ6zEkEBtkinGxyN7OcHQNnKp2cs1cMnWUChpUO2Ihknuou
jaqBIJRDTzZQ/dGmtZm9sj0rfp39ODZNm/a94D4PIGF/agGm3BoCCd07k2Y9xcML
BqHg45E4PeQZ+TaWnw4aXOi0ZKo3WYqDKRX1xlrCzAA4djYwCdWTG/H8CBK7wF61
wKJ3Bg9qszwjJyevTUowUrLHZ9WrUmcUKlu9zeMNgA3DTyTGCauiBIZR8jQKiFs4
klThPzNVu28Ttyu4qyVDuokKcjjbKpJP04VyMaqgVL2DAWahvjBqR+2q8+U9Hl9b
N9B3HLfQJ9EIyQgtQVSRvGTYghFZMLM+cGx3oNRMSwFNyb/5hmzAG3nDAeznrP9N
awHMJODiQ+fUu7vmklp2sJFrd+jOe9l+8qnaHDgrrHq/g5Z/8hQz2PWhM3tcRfFQ
Kdl1LzVj+3eCipw/jTaIWKVGqobWpctozvpicDdhLegvMBdzFW5VPhK40p3gCrnX
lhU0/c50csQ0HXXpCJST8sqpwx+j3ewjkmCwA0s/tGeq/W7k9K2yVNo0wLnLs+g+
QWh8n3u9e+9m7tKWDH56dglD6M11aKMEkTdimFkEyOGq48cbkdV/ugZU4lnSEbiW
9lRgG/YvLGro/4LW3CZR4v8kYWuVvGRA9f68uCoTZlPImqopxz8cHsfkk6RgqWdq
iSnGs5PVwLJVlk3adlXgBdQJxHhPQAuv119suvItheYvaxFdGNQioJspHbqmycK8
bl3LMspX9qjdjtQewcgS477mkpAcENYABCvEF8cMyK3DKq9PY0AZrpqdPkdI/nkO
FdSx3IytAppAEtzLUGkJLzNpZmT0wYSId0OUAvfV3rdFPI2A9DCLrBcg5MqJNK5P
2NwhPH9jruC9z9RYiP9Kt2t3gGWE/GCjg9FAyY53O/V8c7yMicysZgfwUV7zsq/H
JQqp7srEGR5H5j8Q3q9IugH49GIt+O4eSx4b5a2Xhy1S74vrGhB6dRwZJEpH7yNS
mgrCUc5XiyNWYm2fmCWwuGhFLt/tUZyDHi25p+qyPbCoX+rqKJnmyG8b1vZGudLd
QHAuqQ423NOqz1EE3OXPZThlOk8Ya9nqwhxak0GS30kIDRmqNcwEjK/YzJmziNpe
12hl9awySLlyf35Yl2t2BR8MXEAJyxS+Mh2rEhwjeSKKfPg3NQzWN6tYuv8THXkP
f3n1bZ2jTy8sJAOtO1tydXZ4Am9eDJmKps3MNfay2x8BIILgY/vHZrAHhrUS4pFV
FJUixMGIQxD3edSEgsPFThHcXSwPqE2wDw5jnZDm6tCkTKyI4TcP0w7wDinfsve2
Ga2CHRAIuhsa/b56H+9kupoKudn0/+qpGwmuB0+8wkfrasLfWLCPd4U4wzsNxoJg
VED2J8+7LmrNF2Ba2ZRJc1YDPaX5aysrIennQqtyM8dfY7oA9ejd6AlJm6Xry3/L
+pd26s8K3jSlIu4rQgCnl9QZb75VgQeS1fMBHJfJUvgbHwfGGSXjF/l55jYmKdmZ
KawpHrnCkV0tcb0BaaPGanNQ0wPZmaMUUxtLxxtOJZpP0rQ66SDQnnuRWmZfTgge
nx9CHQG4dVCFvPsr4uTvZp6PP+2az/laiCue7tUeWE1teDgBy1kaFwJJ5CGjkb7y
D1FhDFA83B6yXVu/0INy+O7Cuo0nQy6or8TrgBpx00As0KYdkWSz7j4E1idOeYdz
xZbE3vSQpnPZX0SxdhZrbHbkcvnErqPT8veDdXY+QNExDEKHFmNYmEoOUXxJ3RLH
/CFUrNjGxf2fr4T1kIBFv8cJGPlvTm/1iHwfd70e2sS1HfyWM8ygaJQb1rjQs5+y
w8y4q30tslMLLtsvn4iEU8tLbTX06jFhvplLnkCHMuM3FIG0TUnINBPrqtvs89h4
EUQZfRUiOO+Lg+3DIqECOAQtdy96A2lV7JL5uhI0ZScbDjzhDBUBZiDcGbonO/aN
Bc/tFASn9wI/SwJGp/ttN9ogWf5O1L6IjkvyNli1ukCETBaoBj+H+maNMSS4Wz70
XPybAoDETbrQbD1C1MT08VT2GVzBK37L+xLNaelOVppO88hJ05BRJQjLKz9opsaE
UewEIAFBm0axnK3MKaXYhI/JaFWPflrJKI4bHsY4DsZdCOADqK0WvTwRPwCH/O76
EcE+zyPjPclV6ZcBrXP6QWIRq3t6IFNjB47b1i79r5N5jdlFnWb572bKX9fQOGuT
wQ31W2I+nqFJ9yepOT9uNB+Wb9kEPX1wDdP5zICIGU9TPZ5PQyvQw6OYqsqNUqnK
HTrFwNFwHPHD2nio+JtEP3Tf0ST7k+Ji9uVfYNlWWKVD5FrZebS/QOHrmvC0yIVw
C8juMcxMdRO03MgqOQqrGNwpRPZHkjb0A/WxAj46L+3ejS/HTEV1zf4WDxUVcp/Z
4r6jpg86HVc3YoGdWH2qXm7+3Pb+nr1CEE0r/9FkGWQogwTt3Y9UD669TB8lIWz5
3fr7HW8jGkDOevLv++DJ8dIMcccGaQ2+UKNvKnInug2Ekj5Sn9qO0yWa16IOd46h
J7gGjcmh6bSwzB474DPeg/Nz6V4kbBkazMvIWHMC+EvwMq2KsvujjusTvPBID2Vf
Jmdi+W1amZoPBYXXSLiAB2p5h5oMDseo5AZ8BF5XvW8teD4zhPEWMBWfRFfXslAP
vX2kWpMxjntcD4iwSHeEt/dyjM76uBMTs9g6aGnC7o+OvvRiHx6X16ptclP3yTEC
JWPLB9SPLWR3BNZqEn0rBoDz6SHcriFMv1rzkmk3m00KWxnNM/oLAL2JVfL25UPv
8HTngdqP1pJyNs20q9aVFS31sal1u0DiJf4cAN1PC99U5TQsZhe1VcPWS5x2wAge
Vb8W+MD3WiGr7LI12BIP8aQEhKwHktvSyvacHCoiEn+tH3kXKKDGvpNHcRai9e9S
TaPeUuRdtIe3EzaKvlT5IBK8SlqHvXagrfkQf0sDSqqSrsf1RdXXb1AaemNmHoOC
+c4pD0JjOl3agq9EpvAYHJhTAlQPS8a6HogaGYg+1O+RRQGM8pdzKf69rpGPGFE3
/CtKjh8QQKmgw74Bbd0WpB8dHPulypL0PO3cVL1+3VaAO/zO2CIfdhtf5i6H7ozd
lZsmo+zg1OQG6uqHkWonY2D307WMY1AY9RQcecaKGfXodm0SQ3kCOLRWt1x+wxbs
4RQmmcYOob7ly0v0c397mGK2DN/xI6uqrmwF3Neg0Lrc9x9TxcYS6om2xTugqzu5
7WWiaLJkurmE+m1bLzH4ygMVVUrl51vyUzNDIsjFoC2g1hr4CCsyhXquSGCKG8DM
Ba+fK+b4Z8lnAx1KOUUqorNt7mkSbfMYJnyBlkoexb07na8smeIXPcgkdsB2fUFb
TKUBkv9fd76HK34pNzkDk5Lo9UpFyDQBR5AS3YVeM9uz2zKJlWmENvmjwJX39m/g
FhP5nZqGWfvQCQ3k6UlEOmtWkf8svGnHoDSg2WT/WuMIi4X88WkJ24HBmaqLmpQ2
b5Tqx9yD9NCzzWzixkk1OD7icmDUE/rqB2dG+rWyF5Hf5Gmo+2Irqy90VpY12xiK
um37m0hwN+WEWoJkPdmt6h13OFDkx+Wge1FTNC5zNgniOgLcU1MOkr8a1nV9SfEr
Gy2jkV5fjay+iKgJZbgSKV7HqMwOqwW6cPY9jZU3MAufO3A7R2322f8JWRXt6Vzi
hdnckOkXa8kP2iWXbUgQ5XHx99CFAWT9a1wHMjmSvf8k/K9tb10XDbXZ3hmuRiOh
dwXe0bYE3sYW2OPbLnN/wK9hjoP2xIqwOcbcRLMnqsVi3WTAWRsordMTONP+40//
Jlt82EzwDZJ9LH3SFj+jxzCcEz22JJe1YqCtFIcwmlAsvXwprs8mK8MSYBK7evOu
hGEVKcN/t7ZQWYXWyjC8L5vO+85DiEHgoR0607q8seslJutEARVoKr0cmfeUzEjB
W8o2DlEIJ1+hlA8a2Qs0rL+4dSnWJcjt06jrn2jwhe6A4a5pDGWpkCzuJC5atwTJ
N4AhHFqxi9YYxeAbwpw1xCtWQioUpcxx4d5C6RNBI2HOkbB18FDP1yqe//uxarzN
8nG0Mz94CUE0z0tR5WPxCGlNHTaN2IA5wg9bgekalFFKPyhPRe/C6J5YbP+qzrad
41M3kj9ZoVF187wJATTdEsalR707OaYisASK+3T9ScUQEoQt1yhxhwZfK2UQ9zG7
DUYxWfQvQVFnBSNR8QO9N0WYYR0SNH3OMxRJQpj17BhDiBvRALeldm17MiKAqCwC
Vr/16UwDXm0MfJOJsnjYaZmBMibOsIPHJIdHj2dN33IgkUV+8984MWDMawBjCk5b
8d6yMUbNSqNTECOAtrME0FRRQLQA7/qS1aDZNdzAIugxc19XvQALOD9kYYhISeHD
+0N+YbOyQdqsWQO3f8sletdsEGWnmki5LQdmKUXNc+2zlzbTW3oHeLUlo08LZIP1
9yOFdaB1kYQLtk7tryhphTLbR5dvIwG+htZJTaVvCZaxSpXiZ9MHfgLLFBROX1ec
LWgxL2Kg77hKEzezdrgh7nrWA4RCuh0GIMKdczOvs8gJdmPsPa7BBlTOvsUcYXRf
J3eck+/ztxNClNKcv2pRDN0lqkCNeR1twytql0yv1jIQLvtJmEnqjxPaUXsurZzZ
V0UYg2GqU5HbENNNII6+Dsl6zcqBPPpKpInHzEj/gLb3NiHh7TqFp3LQqyMvsk9c
yFD1TsidNkv33Rw8apTiRQpNBk6Em4vgRc2DTWCCyWEvy2eb0iodcQUmJd3NTv3C
DsbG+cHuK8LXFxbVEsXzz21X9XfVaqH9SMsqOxCVeSTPTwZDCa3foUT8ueitfJxD
1GVNWL1luFQo68spjL0oMYIot8l9Q3Qg+9V8/Uw6tJtth6Nxr8aqt6SmrCkzroZF
zQvjvmFDKWi11IPCo92PclN34Ini4pv1dgAWwMENxJhkaSKy7Gnj7x6/YEtrinFW
O0mV2VZ04s/gzCGWNtyE5uEm+/cdZOWZqRmQ8VJfXz9ohLyEzMU7JuOOVdo0rGml
HAJoPVlP0U6Lsbpwg2IkJYVVGbE9mQ/QCgvIdounNwEXVt31aeo9bXK0Gi5YLspa
Tcrale/g0enpKgzso8AxVWdc46waZPiOhXWNp7VoN0juNxevpG2GVOMRfYmXc3FT
IXEdvhz9QW7g+HHEmVoii8Hx6A/5CUuoLUZ5DPBxtLp7ybmeLx+hCUzxeauHSDZG
sY1TYrz9s6+y4f5P2qvffjOqYKbwmyKMkyw93uAQ5bDKxUYOJAYxNrzLA+xUji/7
/YBeWvpZOjun73dqwPIYFK3xceWFHi4NfA/stptGfa1rVx5U33MNmWjr8cN83GlA
6Csb4lhoMnWRGt6s47gjZXVOw+2tWHASK4wM7GkLhkJympBNcE0G9FLVTWKkf2/3
9BDjxN8iglxj/Nh3x7TKgC6WuhW3/ftwGjZAym6rn4SL6hJ75JCmt+4OOiiwTIDF
m9dvXW1z0UI0Im2HZ8164szltmqBw+Yh1ghHyjdvVRysZjEd2AGYl3FXeqC60Erh
kdFtQM9YKLNbCui4+cbgVSf4dqXvTFNOWuRYWRJYFabiKyFQAYKfbGNS4/JWmKGL
OI2ecDO6nkqeoJwdd4wT25spD7Hthqfk6PZ7xUk/SBucTW3oPY1pktkj+O3rVs0S
HmXbroVVYNgBbPHn7EeZD7fGuH4+4pEozA4Y8/lUeUtZKEtyh+jWSRYG7AyWAnKF
zgQRqY56vsSlsaBkjIjoqDT7PCuaZDV2IfZKNQE2rucOMRo6jPZun9/odUQaAKhW
2Fbfy9cfdE7E4vGXf9Zc66Wk/hFleQlv1C/DRSYmJjTpPZOxKtyuEpncxXd8+VT8
qPdxFAUKYdjjcc0Tk51uPZiDwt+MCYI/6F9nt9/ggBDY8gRnP4UKnX1CM9J60+4V
dRePWDB9YWXQ5j1yZfl8RW2bb4jt1FzN7EZhraidkY+JTFe4+AJ7EOLjecA8oPk9
Tm6LU0hhat9+3cAZqZP3VPEqC3L8vdfFYPOhqv9rpHBKt6bilg1eat0MbO32TPYL
DuitYbcoYTgyeBVmFm5BYQYKoRQq2cSvSCpAySHL7NvN792UWJybZPwiVqTgF7+e
jwYhZd9B6QpIZ3pBfXYfi8RG3p1/bLuGxjKHlWh8SHAaG7zeo5q7AU6zoi/sZR7I
dWSS1OSwu00sjl7l8HK7roigDHRJwhGDB+X1DczOE4KEd/pWEmaBjQWNCVhc97Pj
g90AsNXGzWn6WnDyQX9IIzKbplLIDldOvAIk/GG4gYiNW5YNuQFJaDC4RHxQoHo6
sZ3S2TwGJeIGEUWtZYXqi2DfFGMKlEFst8qutZnpqGZSLgOY7YcOkMHbN5NZSsJd
Nx9lVeht/EMDFl1ed0kQbrEA+TD7knGczOu+3l8GXorZ9tPX8ter012cL/ViWBde
0eSIvmF2Zk6fwVNsJpFimjWN66ZXnWWumuKhNnNVA9LiFVrFXWUJzq1N6Fp7jJ+Z
Y7isv6icaBJf2qJRqoAvIfXE26973QFDU2siJSrcDgEq+DTWpmv5EQXBLFIOlxoB
PY6D7W6F+dPtqmiBQJQRVLYDzlOFP27k9bPts9WwxJk7BQ9Z8r10HoSbJq8hnmzB
pkmxiD40hBveeC9mcmyEfS5s21TPPI4nAYWnKzLWQ2bYeHQyJBRBQypc/nKxN0bG
Z+bXogoo3Gl4tvoYiv9AmJkIm0Wb3TVIkdoEuyL8Fctmgo7bbYyt4nQbTp6CGhCV
JLKQNhzoEFLuibr/HdSZJV6p7VPJTAMk385vwksGm0cF7Uyew8uZXmLPNBOXS5r2
63nMJUBboLIklkMPYhDqA+Go1OOZkZ9y80ejK8yYrorpIjz6AYV7A7lkz9aoWRLv
tYZ8qrjMiU5yRAcvaHi3GjR7UNdH1E6LPMCLx61I0l3do5jXv1ujO6p2oNlhjHPW
pg2qJlGZR0Xdj51CfytPoYceUISWDP1djB/HCKHOtP7SKDoH0Hd6PJwdhE8GYccT
iGt58A9zsSSVoNB9Vhp7UWYs/Jup2Chdp46651QD2c2RKzWtdrmFOVxkmyiFx8zj
urdynALAKYk/BnZnM70PaPeAOTlzz4o9T2tGvwYp1iplAkAzSjAZpVKfF+KFjd73
Ynk+3SFrnQ/mN36VFGX7uhLN+AhNAm9FgtOvPGP0q06denT68T7RmQvTfelAT8aw
UG5K6ffzZsgmisFfZo8U8jaIP6cHdDXAL2lz68u/esA0wPk1ceMnggUbI7p06knZ
2NGt76dG6Jkd+5tApy5AWYVVjJJqaKyKS/aB/czAW4hF11FbO2vrGGQUAKf0lCZZ
j/56518fB54aYIdw1a/OWO9Zrt8oSc7x3H2YkV1+2k32yszfRK3JvJ6fNuZQSlRb
hV6ZKYtA0M/gQYxs3FGbi6pnyd0esANho1QZRG/F57tGFP7+q5anUTg2AZIwIEf1
fZclM0QPgL9IzDmj6kXrFAXyJkHGo1B1M0BEPtSrX249EVkvauXDxGjgvbcEgd16
w7mab+F7+7JV4/hN5DX202ufjMVixa3XZrvLtzqcSa1VX4F4x/N0CKeifacGpeSF
QiZI9ra0mAUae6u8WoDL1iCQlSqg64T166ezAFxe2K/7oGbmxFe2SCApwpd1p0kR
5No4ksx/Qkm4fPAzgEwlysJ1Rl2uGYtvnqF7RlFxdqpdcCiMpXXQHKAUl5XOg6CI
L3SJDhpIsm5RomZb0rQNHGvJhT4oUNcfQBF/9xF81N2ytVYDkY1790E556XG90D9
Gxx2qs2n1U1/jT/1hCJwi1R7aYvRWuFLESESxYyAhgA17MODWpoqY+cL+VPf1Gii
A+E03naKceL6KAjblsQXFLWnyHqPRvWp8e9iXo7SD1beBh60FqJWMc/3TsdlhptV
2p+Gm+3NYsYNBXhkAGxCVGJ3MQhHKeFNHd2NW+3jX4VX0CPcU+ZTrJQ226xR7Vay
Jaew0kE29pZYKR2+xPlUkvGzU2RhvgJPo2in3Yvie08bJj0Zzikb9xeGS79bgzr4
hi4p3icoCW7CqFfgCzEpnSgD5zWZ/CIUquL2Qh0r5iMn3vyJ33z0et81fqwo16Hi
Y90AXRModSC53oGhwRR/Qq2Oau2QWIb25q00Nu6ETOUbqiNxjrwBuqvZuHuILFHI
M9pGl35tv8nYdbqVos+NTwpZwDnJzKD7SrjiQm7F90JayGfRsiIuBezBUPBqWdcC
J/nQwwTK5uduC/Ca3G5Rs2FGZM2aFQWM31G/xJhALfMkFyMS2K7oDMVpkT9irZj7
PNyEtGayKaQKWOCHDmTSPPTwowDJiXmb/UM+vp+uPmM7shtzbSmLq/QguaHt/xxu
j830272XHynxhubaoxMYuy334rpBVX+cRiL4sz4B6MwzqO/VVGMRTcf55hBbvgS5
zPZ/jfFAsXXURaOOKW5ps5JPNY5fNQruLJ3OsZd4ddvj6HkImrN8/BNsddwFnDTk
+84GIwhrAAgCvmgy/vEDL8sSifUXgImt32SxgavveuzgFZXa4CMLAnbqXDEmRzi4
80hoCEdHMyOwncFP1V/JpcDtqSf8p/0CT4jbJev9hqYoXKQLqhSNfO0TUnFatSVW
yytszZiQhyQROQaKxPhsRYgkJIMuoAoMAzBn6B35uGRdbIvAjKcNdm23mWZRYcef
/2boIWNuxd5GawT6ZR5JTgmBTJYZs4SwsS6jfxcJ3hA2bV04vEwiS4V0vdcNIXbI
05DvFPHmiOKwDcYlBeDk4XsBGMQXgkHMsyofsTDn7SdDt6asZxyZFbLbUZFPxF3Z
WH/3a8ypL8qGYToo3qTxp7/bgXvGhgyyt5iP11J87DZjYZcSsrE8xWxpHFZhiqIN
SyRlQXGGaTQ2YF0UP+1bhbpz5ZWUrohL0KFXJiXv2X8Dqbt36HAIAQKcq74ErjJU
luF3bnnrYStpm1wwqAhDAl4iUvT4GenCd7v14Xrt07hXXSgvBzw/K+TWiH/IxtxL
1ABi2T6l46LsSGNcG3p4K5DrgzAw7z6t6ca9b7/uJ7hVAQja47jSGgoWzcQvrHcg
yR2G7QKfu401+RS2BNiI13ykGFUJ/oWMSyIqCsyKL3dYto4CJeayzSlbUewWXKkt
HYjCXhoMcUEhWBIXTcwVCKJTOTrypdbs3SU2bP0FN+jn4+p+vfjfDIe2daOZhXTj
XpcqP0WbcVRx9hUJ9EqgqFIa1tFSxyyve3I2HMgyBywG2uKZsl8LxhbLhoJJatOS
YoTL5m6n1je6lwi8c1y5VfTckjzJ1JXVJdYmJiCV53TBatrWz2DEtxdSfFuWwU9m
RzVw5K6Qgu7AY0M+1meukm/WUuRvF9umLfyPWzBrbloLDHlZ6/jdV5mkVUFTnVXE
UJL3CKZjJUXH5S00x3v0+7PEgpS089MMCKi3Dln/ABYKVmlhUDgsRgqNQkWDIDmF
UT1IR70a5Y1qNX60P3yYsG+cXRCUtwmS25p2pi3ULUxpyAIUrdaAlgH6CBX6STUm
ISQM8VMyR8WvzIgxxv/7yhq4gjEm1z7Qe93G8c8ynXTBHx1nanrJ68tjy47l7OcU
Jap7SocZlkZdV93MmDqX/H8nULo7jew4iNWk8p/ex6gbeG/+SoYSrrD8RCUJ4T4d
ETiZ7XtQ86sonyVlE4yMRyQGL45rjUx6TKAwhUBQxi+RA3qL5NSj1IDC/RX6nUNu
zLExZFS5swsqh51q+jGtpz4dzNweyw/gQIeBlNm4x4/7k9RiHftkbBmNc0y9DEZp
OhqZPJ6fygszTbG7sfk7zVBtsJQH9leC5jCQt8XlvXb1vop22EB5Dm4AUS5laP3M
rcgRGsvfSjQy7JYjQNeOf2ua0ZVRm0/PvGK2Z0pllDaijwMKofMaqNpSRU93rNdO
M+V9t4HBW78uzH7q+yzVrbnt0JVCnjUcnRe6jE/aV68HWjp1KihsBhkrl5DqPn1N
eyabegs5L4xEe+SOOwDXsVl2Ss9vu3iEhheWObgRY1o6rU4HZRtNIVwhLRFGgvt0
rmzs2G82hPyizmMH2X/bUj415yy1q0zep8AmQbQDHneO18mWtFpVrlDcC3MoCEcf
+bLHiOVx7M9D/QhY8Gy34u1RSv7re+uu+2GN7KGA0mcEp/E72HnltEZeUzHNbIQy
lPk6sw8PCcif5fzFMxxq71P+RhCQqNCDgLzuhMNLVTfOSu9UlRzFvoraNqLZrqv/
P/Vy7JfZ4a1iWnNtNKicgcEGfNI1wkKbpD/yhHUgHe+QD3VRQ5MSHX7y1BWwVu33
bNniz9A3rtyUUqxhDl5zbZ/QOKboq4MwIvO2unVkzGZO5zCSXetcVX95Cj22sT3/
nc2RunRGQyrUDudbyXis1xTUgPYFOJabNe3OtGVqWjhHwwtCBWL8PmPfVzAf36dz
836Jd9jB3NWfKhivHyHFeHaaZIa8AY8eb5KIaaaUjteQeqZj0a/Zt/8ffI24yqM1
bSI6POn0XbcU00tz4dqFVdHpa3g62Vh1n2AR+nixvoxe7E7cf3k8MzSTEVTBa49j
VkiUMtFlV8cp1Ew+ED2/11Znwk4LzGMdW9yIa1X9eDahpeI7B04PMZxigys/0/ZW
x5K+SWzxpi9GJF4/+s9XLMOQcuep920jPmvzeLSLBTN5fcL/YOKzKGUqVT3SPirj
r30Oi+67KH0CROWFXBvENeRLGTRQMS6+S6ePPvT17JWJW2HzOcR59gV21ls/Nq61
QXlktkyDhyasLOlFfUUSG64+X0yq6/+v/imqDVHZvC808CcYJjfOEYALooZJ01kA
KX+6z+fSRHKTlo0iVv3Ty/iYJ+V6wU0PHMnTk75vi9t87k00EBIu91814R6On+AA
fL1S13I3JODN0XhJGEGioUKUH2LZIpBr1+z3/c/Y6olX1kW5PxlEWQJMmAzUmv1H
yGEcGmgXk/82p7Ow4fIWmJNPkuyX8XK4lP/LKOqfjwy29ded3M61Ny1iXGuDjY+8
uUBJm/taf3RRi1FIO9S/ueLnm6NsoW3LEud8pQhCmTOuiGxRyLr+C6P3qkMg2I6V
PNBdRAw0M3t9ZstvjwXOIeGfKOQY0VARO0Yg7UgqbLCVOkwaOjuUoah/TEjX3pGv
1BEUUfjfzM7eo2XvoCCnKkuxz6We+i1rXZ3NPlKmweus0aYJBIF5wIICKBZsyT+A
Pv+0d3VKsqBYhb5AHHBwUBMnXFUyQq3SSe6PQsL6paSRWntT3mHyxh/8UdZ0Tk+H
KZPpeJkRIUgO8Mf04I2+yJ5a4k4z9teFVSn1sreTtBlqguwzdBosym++SU0ogEtv
sSO8jUDAWxJ8scc4DGfWbyaMNBSQzkNWO7WMo9oHdgHnZrgPNj/smyMpSIOL81C4
JdsSQu566dJGtfpv8Ud0XgOu3Dz9s6U1AyU83g/C1rK/A/13dzQWqHJi0lrvWrIU
PqCutcJzGKeVVBdLD7LQGzhad9TOGZqOphQnrHfg4CWCoL6EXkTWQ3iPQYty892E
E4twyNMtsn0LfJkqTOw4Ydag8/h7J9XLTlF259Al+OIJdtOh+TS9wG/olCfePFAZ
q619YMXJffWZLWtXW78WLF78FL40W9B7Hk6djGaJC2OQMVmCXRlLLcrWrDBFTfq0
ZD6UQ/iGmENq8qAPDbaE6T6e+qOmuvWFNeSFwxo4PWykgmycGacVgtaN1QJnhRi1
2tUBzi37XNkx5jOLIEiO9r9qM3JGxYFSwXsG7SHgUGQ9l3rdWV3HHpvdeSqxOCbD
fhmOtQsm53uUjub14WRQoegKgItqeD/Fc1mX+j74qRaJXm4O3ATRfCBvJG8rt2lm
0uoek0EcjEXX3dJ2H9Z1UaVZWgSsOS7dlRd0wODhYf1soN342rWcd8D5cxWTKoF/
HQutJrXO1S0Sc+qLLPukaPUU4GAyRXaW+S6XM7i9WZw7usrdTySatYYQQNmSaELY
E5Ib7Iclr1XwRNavYPUtxike7ayu67KZbc76H+vwJ0KcpnzgLzs25U++geLK8yfo
yKE3H/ocPKL1gOk3/7+R3fbqInAEHDmK3kXWhXnNb1t06R0zLC0e9QSeaF1BnQh7
EOmP8GhNilHcq4MfBPydAjNvIrZBsnE2nercFV7AsZTc2kz4VcRaq59qeaT/0Xf/
z+yGVRtTIhLZgNy046+aTJEXAD2O9BSD6JDG/+VflMaxbyr2SlaooCu+N0HuhHIu
LBTEXrsBuRmXqelPeWpd7TMnmul9X7rZTqImrnJkUOyBboYL+gqTXTvzuZztZ4qc
BUxBJcddr690q7b2T/WgJVffPw1dpmhsZFDdfBRQPdXRrPxMnRgvPAv0liNe1Y0O
PEUOvMq057tttsccjJTxwzeh2s2vlciZNtijt3gHFLZYDJ+0dqM9M/Lx3TZYaIgB
V4ELPN37GavBS7AD+KpSTWg9usUqzTmMBw6o5jkI5tIqy8slB1lvbE0ZP46S6lRs
zZTos18+BmQMvoRRwshLAtUB7sdrUzrTgTfeJmhLvyO8D4LSFc7rZbXuvtK/PO0H
Z25aM2sgdaj874p5XVYh/tTbKtuxFPFx97UsW3A8yNg8QATV2pgI2hBZbIDTOlMY
hlZ5SIP15AXE1kYSnfufD88YHj/G2js+BSX5ZjB2wbRxQyoCUO956opvyU5GYXJp
3aRe2YK4F8mCmPebsYSoWH9GHLokng9ipRYyZnHl8XGXjyguhgv5RtWWLPQMFzaf
nd+0UOO85eUdQXAwbf1c5gY/pmnFsr6C2Cgmd5ADsdOkjuXdeWQnn1u3EdGAh/FL
aB00Iwfj6yx4k5zpQY0d7q+xJO4jTQNhClytP8J7F4yq8wYqgHzGJ/bQNYTHlQH1
cPMFoZTfnRCA0JWSwv31lHdw5CMCO1LbOp1ioovkKK+L1bAwRDlrczO76YpQCXW/
tF5XlI8GRk7ErGmCSW0ST+RbYish2Y7sv6s4ajOAEYUN4Co+jYCYwL0+hf9lIw50
og7gmrG5TtvUifXsQLOr+zYxr0Pi8RJ6UFST65+IzBt3aAVjgOYFM2JgtZf+OHJI
Lm5ch9xTFAv761d8iM6SyZOvxEI94y4NQ+T7VySQYMZnmKKKKBwzBDKeiw9lvoOp
1PSQe7F35C5sOKu2+/Up7hqUxZpMCZVWqMMGFkmoEY2MsyfoVQwW8rLQDC0YDIyz
v2olWnVD/Wx18vlP3Phhfzo6eoxFaZ2s/qofBUmk+uLyzFSFlrx+3+jsSqTFkpTX
o1S8cI/Ssg7BGxVJQZ2z2fU+2NxfOlDPqz25k3NMFapEaVFWr4YHckHSJRjNr0UI
8xs9cC4VqlezievJMIcDXQdiA73nnNsi20yQG6zVxQf/oBwLkJ8v18WFdV5tXONK
Poaw2ik8p2FpJXX2uPO+NW/YkuqhnC7XAv69v5c/gSHnEaBg4yeHkp6U14tvBR7x
dxyiYxGlCQzKjTtiOXp5gzF3Q8U2cpriRaRBMRWPti03LE7hWa1aWivZvGTUEn70
CRy3rLehj6wEMB6qHF+7fy/WOvVD5F0SUgJ7/MEZCl5iCairphJueDMuIIT04rHy
a2nRaSPAT/onZEfSjs5BGHdHJP8MDsYBxmBsapnWMwx8ebOH57kb9bjCOfxd44rm
cixL/w3dOcSU60JvEei/tfpPzXXezR14ZWTFxCf/x0OyOBR1Wg77tIUFewkWAzQc
auKJZ/QOvjSC3UijFivs3a5K5Uyv4/h8QU9sH90tt6vd4ZTdQSFPM6UHDU9+IFiK
Bv6glq3zgt+Jap3+e0YB17pfTHp+LJEGzYrVqURLbn1mHYYFG3rWZB7YL297SFcm
lZmex1W9W78t1HOuCepywHkXDqj1ZXWyy1lb4v99jd3jPMnT3hPn0sxGv7f3tJAb
PW/kbciqFjscJt481wcyg7LPMHIOuGEjYDaV3QCjBsEd2EHnQoGzhdgq3DvXqGfy
pSE4XYWBceou9/UEemLsz0ovtQdXwmw+VlHrwfp6gCyp4RaxqyL+LjDf1Tc1Ky+W
gJrBAxRciqA1wSK5cAuub8sSIbVnxa2vFHL6DRf9WbHMO3XOmzNJQWa2eV4vov+R
/iaUC7+RqkWzpgxUIixyWzfOEbpV1+gr1nAensSpISd5j9wPkXSX/VaqiBNJjU+D
gKNChmYxKHp4X/RkyH+yXyM1MRSz3bWuRaZN6mZha1orpSOjqaaNjH3a26u8GY/J
xVdUoNJz1ik/KdM1dSyjkjoMQIo+fP4/tszJaJJNTtIzDe4zcM5ixqtgosMvA6p+
CxnBl72H1BDaT4sPy/b0I8NyKF3zyoG9WLS5AmgH+F1HirHygV6v6q4g+fJQwIy+
Tdbq1OJHBiYk2PWwX+B6jTs9vLIK2sW5mB9JV9ab8px1TlJgc6mN8vCVTQpYRgk6
izMhZAf1ah86+AnqggZ2HwQAF2fgHG9/tKG5saFdXeMNVz2aKYcXKEEu3Ttmx036
m/er4NZphxNTwlI0O/WVD8A+MjQppR45sOgLrwsaHEqNDO4Vwp52ji83j9nJF4Km
MYu140REV2BETCMptq391hHNDziMufArnC8wyOE0DrNduci84PGwhiorkFEiajiE
bRZaVGwbPwvNpN80yaKF1WUrKAZl0YZcFseJrhvZ4lMfErzvY9/MGG2vKFvdjZxS
EdkK+NyaVU5XgkVxP9PR25j8It+KhzVE8x933C+oW3Zg8oegVY2aNo4oZg8fYTnb
ffaynKeV2acfVBGu9I0uDQ5G+QsU6kM52inpfULbsh0WHwCMjhuNpNwF+8Ggp39r
I4XGKNY8LjEN3KcP9/yB44DUXd+dy/1Np+466jbP1Xvq3/a55hkXFkSzPWarHPeZ
tPiHdIJlCXkkoA4jwERsClnKXtUpRKKQZ1FzXYhHtvzEGfm6zbi4x4OdJHZn+1T9
PTDtm9ZbUDu6GrsMRDC+C2Y6/dKTRsvv/8EfddFkZhXxabCLPj4edxOShH0kEXL0
q4DL+Xyv2NqB52DDfCcGH/xlcqo6LT3EnXVq2EAFOTVMic34RTY3fCZqNlSNDznF
E3oE1pei9TkW2cCgSYk8lWUsqakRnGVZzyLlrqwVu1ot1Nn9E618WGQTkRv6MUsQ
dyXhJ9OzxHSRoBjRzVKOJ4A2/8PTdWhasaFnYcTKBuHXoSkIEwwu8NM9Vd70iaMn
kEz5b9outTpM2nYJsHMcT3OVM1DF+ALBtk5r0nCVob8xJpOs2pFzFG6Cd6S4EmtH
lnJSk1j/ZJYGvvzI8v5CPIX5PFa/qChKWK5B57xX9Oak52jL1hmsh0NdlJJEhKIZ
69fiITNGqZBBzgzezLYy8WVMrfmUm4c8YhaD6R0IzmZcmB4RQyfcdXd36INZ9GTR
`protect end_protected