`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlnrEYb4p1f4MxzHqe2QQTvATcMRV/u1Mw0wljRqXMKi
y1tdfa7fXdDEGY/qqdPZdPTtT3/69feQs0k+PNSCn1EHjK/NM1UqKRO9ieu4QjJd
Of4FTISq2bi8N5GMdHMQYSaUBHDF8IGzYZvTkuf7lqRrf1bOYpmlJyRDNLJbBx0Z
qMNsGUbPoqUhP1XpE5L32r/yNtUTxyezKHmsm1nyqORKivpsuFK1lLKdKwVu7bYp
NxxEZBdgMndCnt8DNcUSRdZi2xsqV/pOvAD0Xg8RUKo+l7poCFpOwnAl37WBY4jJ
IiKS6E9MbxVQK3KyZfkAt1rZIANtZGPER1T0gg7X0uhAkPb8GXKiNr5AJIkp4d7x
jVUxYdlioacJdbEnNQp1Hn9Ggm4nbWch7wUplRLNXr+iMRVaJ2AqmW8BHllaMpRJ
YyU9LtdBMGEWCSuZ9FL6YqC2x9BNIVHilwNBA6Rwwn/myTwcpPyZRNMvYQsxrrdv
U7+jl/jIn63ouaU6nJ0jxVeoK5mOx3aqsfHY1Hc6RKimb/+VkOxmo4XYH7MEoIMh
QvHGqUgFca1Fl8yzSNNb5RSos1wQdyloO1oE3QhH2gTKMQCTv8lcWSEIoDFKQQaY
+rRuUWnDWcBPp+YS/RYUnTaoK90xg+M1QSt96eUO6Y0hdlAqUl73gnNfNHmuCAy2
Agctrb6A6bIXymMR51EEx2BPeDcfwXvR+b64xFbDr/Ah3Ra5Ui6d8uYLtzh4jneO
cHco82N8Egk66m610Jc3gqg0gv7Q/MC4EKC8HSTMUItV2m5D4OC5j8lf3ro9Jun2
wTlj90WDetO4/ub0BQXqQSeHTshwlc2fyus4/jDRePueSOgTJXtdzDYM+Yc3303x
ufC8Mp+/u2CNN/2JzRnaabPGz0qYGlVrXwgx59xwEWtmEtL27XmKN3a/+vKZ1l6O
dqp78GL/GqHCzzLdU9saEpeey6dxrc0GW/jsJIQ12Ej2MiqkCHo6dKz0jDq+mFRQ
NISf3eryqp8+dhzQXOnca6EAOtcFUWs6JnAedgvjeGZTRk3npbZDNvkbSi5vzw7w
QqiL5BVxup5MeXCgNHxgxvJL00rLUikZw/FiLhJ5+f1ybXl8Kntnp5Hzy5N5D6n3
cD1AmZSJIL+Pjb5X8ROqFKCS/lsw7qXpV7Ye+Y0Sy4mn7VoKWKsZWuvhcUmIvo3Q
1N5lBBkxluPy7hI3JyrCRWG1u0wBMzMQJttXmpRKw6ZI5ff8Rbop8W6oSLMqfz0z
ZRf5TY2i9MZKOpXxXBV+ELSNsnEX4BMtqpUl2q+dP0M53HQcUJLKH/NyhFvszn42
/bpNgGd1SEORMJC9+5ktrs+XC0scEabffBaifgB9/n7iebk8kYO4271RB8pyP1dX
DHYwv9ckpljv0JohDA946tixHtfXaYYypNr0+goqHrOxkQ1tnQ49dFtsCYDueKja
LSzXJkO/xA31q0/vyPXEAwa3zYZrIpaoWkY6HwbSyo3flqHZt28/RJn3jjJwm688
l+gTxx6/uMi76Uq7t4QasHfUTAOtmd3wFRkwmewVC0iqe09aph08QdyeQ4ADc3T/
3iB+eZzxFcOzlt3jyDOEXBm8iNZI6uvkRLDmJoA4BZFO0RJZRRbrLAelUVVdCFA5
z2XlWbBD3pKP6I9xczlwAH/BD5JzgEJz9t75V6+3pm/gwMNwQAvOgBw6uXZcb/iq
iQAAUsyzw+9pJnvfA+qbhFEEa7yCCWMWk3qgftJJJ3lhWlUL0SRnsIpH5/51cWXt
LvN/QOfPPLUXzg/VRrhgCmcjoZ3tQon7u+wkEwHDMTQyDre3E7lOcaLMPqi4YTwR
6M1BPQkczQOVEcffT48erTFkKqrhjoc6F8/bJ2z/qUpJJqWYxHg6m9mqoxlP7U5+
6aB30SkOplIpV1WtzsQQvt89VEikunUUgMkneJT1LO0qcOT9+GdiVMe1gGLA6Ln4
B5//vFeVOxeMsscDYgivO/WdVYzPpdRNnMf+hpgfq6uhqPbVU7B0hEDpCuxLtwwT
5SI573UMAoTQjV57BkGE7FiS2+jMMDvrAI+ivyUKrnEOHMn8Htqf1PMZ+fv5KOgU
sB27RFnj0Pj5ZPukg07daZlZ2ODIMugnMpkRs+slzNPcNuvQQKsejSoP5pUs13X2
CsAXw0yF3q65b+gaa5LOLPzoNoanBaF77y4cpqnWrH2KYaOvnGkNr8GxxZ7CNugm
gag9+M7KMqJDlDC26FC3+QFiSkVujdhhhGTrTnNOBDsfKFFaxfC4PjXKstLeL+cO
5qAL9xVON4B92eQYTMcw5zK8yQLFUGjNOmQFgvMUpLY4w71+Ie8S/8iT7+uORaAE
lT8mS5n6gBiHtpkNbngtt52u433EIdJ/IOaDecgmKppEKt2dgt5W6Z4LTj8+bKjW
JSgOCNAXaX5qfZwqdLsdCRMO67r6TSJrlIcRprwHdHjRuj0dd2O0DFJrRye0GS/a
SDRxbbc5suD2923o8B32HB+dFQ5UASIlLnnWFrmVuMfKRlF2+ClbbZyZakr9S8qJ
+88gcB6yMS9tTaLWR7NtSGC6YLiXQJFxXDJNo9ZY4wMaQoaA7S6eridL/bZ4ke80
dym26h0wiowytnLzoyiprmmMP/wC8iouWU3nrPoJPFVexIcjVmj0KIWo6xtNmdCj
Da/BmHqCyPnwGVBlobiGuPr/rq/iM1YStniHHKGkhm0uLVD/RrUryyYmE5FKRXbo
gJ56SbTn/jGph4mh7puB7HDtD7OU2BrxnzY3UQ23pk32DIEK86/1YjJ8aui4VmNt
WLda/a+7CBZlz3IKcHTUuB6z/zFuL28k1x1b9vDXtXcYim79ktZZuGxqmKmZxz4+
ZcgMHsBuLe87ra+X4Dc5kZWWCKkK9nC6uvVZ/p5J+nt+PZrz2MGvINbROL1LHYcz
SIyw9Y51fl86BHA7fjhTWGGw+iIhYKtHNsTBynIwFxOUsXI+eJ1i2vcvHzUMfkOo
f1w6vvFRTZvpuzFoqGANGaNcwmFAGl9g13qAKG6QiI/BWPCWjOLLkJoOXeOaxI6K
Gw1uK82lhR2HWjGZSq7B07eRM5vDpxtWHHYlAnly4QQW0Lp+9Nov9OLoQwqc5em5
FfpBfRhfRJzOiajzRJkhwC3Pw+8WPUucMqYgfeJ+uIMNjKfKsFC1G9LZhOP81OJR
4ug3CTOgzrBRHwv9kN5gQtviKM/w0i/JtZ0Wvn7Dv1peu5q6dqaHvZq544v7hZsu
jf07/nqGAvrpyp6tgoQ9eSEUN4AR7g3rnEFQzn0oqO0mTneMmOxv3LFmYemeZOc3
epP6GQZBgjPsXILFjwHetlqea3RXpOgvWws0fgq2Nlzb5dkeIdx6MWna65QCCj1r
FaR1dgA+h0p+KGhEi3WoUhtSjiw1lCbTPKeauav2FiDgp+gboMNzV7wEbxapw9u/
Oity5ShM+irVXFgOq6yOz8r3/fDflUP1k7I04h+ZL3OFecy3VF6ROu5B+CDwWGCR
+SEbe7cBGnYZATImIH0QdO7kVAl9J2SFn4Bg4BShUozgSZ3suzZwKsDMC/hmQK+K
GR1Qr6m39H2Z8cVyBeKKit8X/3LVMnHb/HBKphHGRi6irB2TOXQVgfLnBdJ86+Su
HHB4N1T0jxhYPl7vbNdHa28KzKRNJpgTy3jlmi5MWO+QAbN6zZl/lyInXC6viyte
vUtNAzltLV1n3/PQPQ56+dCy+3c98SDsCxNLM1+5mAGDyITX5bb2zvKKn70+E3xL
TCwtvPhiZT3YXsEUsPtxMHV+FKlbpl3tnqZYnogQCI8AnC2eLbBz50Wr8DSmjODX
/sAwUcoEVTkGStPiMXn7t80x5HFoCWCoYz82i0yWyQUHBms5l4XgwCFH7GgQsJG9
5J+ekmVGm3sdQ9R+/KfSGZZOUx9eZMYBTHUf5fwjw+XmHwkQQHkb0xDjwGAbazue
JXVOtQcJsyfgNYfYrWNXa95NWDgvkPa6SOuwFl7/d6miam+mqwlmVOb+HNzzMvou
iMPdAd/6EyQ7PgPJrRmN5hYQHPry6Z1WZdxG5GztzlP3Qpi+MD/UgH9ME6gF1E58
3Lejq1UvrfYp1Duuqx+vWkNL8HaOe9n4WSN7+oWDP+z7OR7+buJcbse+pMQ7vju7
GPcVynP7ppNzouAu0maUhSE9H+9mHtGvN8v8Nh+NvkYSU0NQ+9TZikCifOL0wGO0
a4pSM+ZgFFXOHxMNtygCS3oqPtaFM634sPTWbAhp6MDmOfr4l1zXE6net+3ldRsh
7tsX5ONgVRG7llZEPxqAxPhw/VrI0UJn2ipvwXZuXFKYtLKvf9CFuPKJGJhu3o8w
Ux9NcNgZ5a90H6l3CFoRw0rgREigtwtb/O5katvfW5kM0ySAVYlEY+QPXmJnn1Uu
X64nR/Ct+40NMy3lasFpo8EdsDI4j+2J3fLSrKRHWsNxPf2MvuaojWZvwIAIDM9j
tGQjSnPDu0wks6ctrQxVN+FSimcmzjF/u5I+gUXvy+k5FrJ3KstJVf9bqTyXoJFJ
4LOam0Tp3qVWz6meg7stQeiF/6wrh+Ia2leyU+i0gMNc2gfCvmNfzosoeLlBfyga
RBT6iStk/liAiEMQP75mEmoRb0nfj0kFI+VgN9XPkh7U1tCWlj2Lrt/6birqAvWL
bQa4J+a8Hg0dEObNb4w7LLFHDQ7m4EslXBRhD1fhKagvcfulY0cjautXu+I+0zj7
/K7/K5Y3sMrJbAh1O4eSdHQew15M1YFhg+iiAm4r/dKjeh0zudjLbJ07vtUMLi2k
SkAhoqK7jJDXq7YBBQFFF5MSogyxy4MJB5DPOkn7iFFWdLYLFKB0yVvYQT7iaY3I
eLxpaaQwpZHCoM4mVVPlFSYi1MDDefpZxIOn4nCWzTnBDKO1Yob18wHjSC16/ysr
QtojvXJhcnCkfycMsIW0HT/vw3qz0LmrxpkDWk7rprXUrOYPjBFeZ+qaMGCaaMmD
09zl6ZIuvykpqIHYpioPXRQXYm/k9R/JQzHFROE38Kw6Y198KRRAk/3jFS8nhIK4
fXxOivQO9f00ejkRThbxu41dNvzxkyGg5kS6GXERTVYQ9IA5fMnbuhyNvlAWNJrS
rY7tr7e9srsTBkpn/FW2AfppMCVipPbIKkvMRYOo26VBazF5VugAfC7uu1scw8B2
NH2kwN8ojzhe0UK2Qg7zCVuIyhKPe0t4hIWwzwK/yzzHd2oh+awfydJmwuv7CXab
+v/JbRzIkcWG3L8xIvNWLW4QGudKriUH/wLP+8pVvlF9MZ3zgJrRcdH0XmgaKhs1
wH6u0q6CGZ6WLz5c3GD2ZdHXifhVYxM94px/tVAnMwKRZL+/I0SjRACeK+6I29Qs
elQUaaTLK+biBlp7zVrM78OvYMVUrPyZDQH3tqq9H5mmP1OoKsM84/299vU+8/ST
NME8bMkQvhpFc3k0aEVDdqfDF4ZjbKJMRK80ONjC4fzVs8xJSIDTCEDVW4gTTHCf
7rPdsVKW82H5omlMqG5gY0bwLjT0HEkNsKabwammOnjsfarh54/5lV2eEQZI8Syh
cpKXjTeIFSmjxmqLt1X0DNNtm6nPcN/Uy18cYfVKeeBkHemJv6E4SlgSzsOb9P61
SQKAtg9SZQ+WaWq/hFWjFobyt03RwK74EfUMyqCx/i7e48llbCDbeGs9s8dsbGox
iQnBnB9gtBDqCqrnouRnbjZQnTmOkQfeUILxedoK/f8G4jiJzgIsUEAYdqiPJOy+
V3QNtOrPwHL+Z4/pLNlqhEWoZmeHKcyugxGa3Z66UmeMUA1s9E/gBKS/FN5H46h9
93cmEIr9NgKewy0jvkpWxFwnxSDv0pzgAupQnoki6A8KLFTW1ztJKImI4+FA5YKH
qYgQHQtOpXfHIKVtwSLCRryBox4qL0x+RgBl9vF5DQFAl1Ca3+RHNqE395pmU3Gv
8mmBjOD8wq0NJ//mWMhnjBYJ5ndCABaPuMbICEI9/MEY/xGEr1Vviab2xKx+ZosA
Yrnc3XJi4D6kfOjU70U1pAucX/oxBm/lqfYmaeNTutQKJYUijL235GDPcDew9/i9
IfAPu74yOVBii5H6UeqNr77vFH0Rmf5Qt7p1nBSQDgpZgOH4/otIE9ODNeOYTNt6
KubLnvcNjDiyx7vxj8DC0MLIWFp6n9vrcs7zaoFY57f5gcma36jwgMMh+U2LO2ZH
TbfCyo/fOVL5ticSKQ+sgq99c2iVJNGnUOawXjQx4vYGnUPQp+zVMMFpfDaCjA5F
VU/qohUfeaA8xi/zLizoSQx0a2vQU5DMWRTTL5wiYRVWrb/U6zp0BVKmW3YMMQAJ
D5n1KZrWEwtVVIwijelVyE6mVg9SENoFs8dVoC5xvYXdPI/EXgPw6hWfW653OA2R
+naj2RF4i/MV13TrQVsxMLE49tFnhbC+yWJlk6zoUJ/KZnrq32AYZhZzLydRzMmU
LcwPBm7qBF6kE3jhvIFaXKdrtQO+ClXzarRyMZvCVJ1dWvImVEsULKkxUPARRJK4
VDXvjfWxLpDwkDDc2I3b4s70TJ5yjaMIX5j4eR+WBbwv0LjkWNcZem0++YEsxN3u
uG9hgLznKH2+IDFRPvXHT3sXbAAWdpdZ36qfatgJd/MIXgHc+p7CimOkX3zPc4zt
SCmZ34rpuGoWpoROHcI7WIXK3MfEPUQebdpyMP0752E/87W5/Rv74FNlycjd9c/g
wjCkluJjhgLdhJODMwzfH/102faPVYN3MavsIxC4hDU0ZphhcpujZrilnHz5UCnz
DYvsb+wzBgLr2Yh9FCRfBKXgURYXCUm1R94McraI3+ZiAG+a/ZcWQtmogS8SBKkt
x+nXs8HlSO8DcF/tfVxYXQ2SdYZVwx7k/qoi1sw93epagCuDvxZvt5z+089SLWmL
1jbMGDcfwcn4bbcCzrkFCT31onc3ApCF5qBDXIDQL2k7TWEkwMst/yW8yb17kPSB
U41P4XQvntkaFkJ+P20vOq/fHyxpkcZqTddN0+OB0HSwJNGT/ulYrPLigznKZgWi
AAXbvxwnu1N3DSoOLh02NHH1reF6YdD+OaHF7C6p62AMgybwDCQdWUbc/kZ5twjA
gMMUU6tTamb60bL6MLFqW2CZdkbqbQv3KSQon1dyAkVxuwBEaxrC/kAE2CPb4Gx9
FfiVuFXQxere7QHq8s4V7hNklDSyKgLmyEg7K0iq5mzCamO+K7HGRjYjFKwAlBh6
dEybrsDXwK7jI9LQ+E0gVmZxvl7+jEtYjhACWOelF3WXB8yvKH4+wnlV9/NaQBiR
QUMQbB3xKRm0Kw2GLYJDsZo3g/tL3VJLb3x8yvcV1hjetrqOkQMsoKnOi+WQMCFy
24nJ37ll5OH5o2tOiYIJmZixBbrsxSuPP89Id79UtqWs/YrRH4SirNLMjJnOf3wQ
IhOC6LoKDTsJ2Tw+ZNA6lSS05tntWkU/jUelWr7BlAYS3YrEw8swcj909EFUEMzt
cv/94VcYmSj2mb6CRUTNHX0VSJloR6lEMbzjLtbUvqxSyLXrgRJKF+h6WYCHu7le
fKSw1d+A47hkd8y3mbqUxEkc7Yf6U20rM68SW3xwSwgtzqo3fpkbYC+yTC/pPPRh
4ygerQb63QqbAKQu9lDwFJfWdvmn6YqRSGZ35ccQKLsdzn3NL2aBs4gT90WE9gnv
xVaTsK/hGs16Vswbou1G4qGRw0j6BB7HMAhIGWXojt3DakCwzZYUDawA6/UMPjP/
VbkdiBGYH1MhLT8ByMI9D9dwcS08plEd5xNbu+xf7b6LAy9c4/KHYYVOm0IRRH9u
Y9jvM7TIdYjHAi1+rjRvxsi+paPO50T903E85vxJqF96PdlhRgPCPrHZvx7RCNp3
jax/4t/99GXjlopgQcbmyuCOHhhZw3lupDyACaec3infl6cB/8ZMd9WhvUzeVDuG
kmgy1TOfD+9BVzVqSJmyuZF3VsZzbgXWgAgQqd/vONpjIu+CRazuMgPUc5IT535I
WmAQpE8Mznlg3Mnql3z2B9zCtF7xtlPyxv6K6AzeLp/QX9pbXsevluwQO3pOM0q8
oL8HOE2nFep8M268tVR8JFh/l4+fHZSCLWiMxaH2Ls4KpK4nNjv4rC6e/WhYyeYL
sq/LQZLXDYhzhe6FlbjUc3GPK7muDrGMlywYVbw0RBV4vvxV4BAAuhRJYa9yWm7W
PKTDfI+Z3BpX4gohL+ruIoPzGCpn7DxECfIln47rFFv4VBTNB3TwpHlBSKn/knyn
i/F8fbN5He8rMVSMyyTq/Zc9fEb+MRSRuxipxMUom+BfCAzb5zJXMVajEUoFXiWT
ijilnUwN0dsbQXt15o7AynrmDsPxPwgYorEX48ebF21It9W5jZmgrkkF0R6c/EAR
iiXfQprJZc9ET06JZ6rGiJeUECgAqS7NtP+n1KatZSDipCfXNBBvY5i8mVwfh0aZ
5tRLwwIGZV9ExZp+gBYF/4o3opVVUvaaOmg0u0N+cbj2E2suZXzcx3vscK1Pt3Av
SVTISIVBjMRO/ZaYxbk2gYs+m0OBPxNP5+/igNDMD8rXgzjDLNKuwPQFQf/fJ+dZ
2NHq8/X/2gyPE6yvuAhPrbhHO5aEMWMUi49sy+jLdwBEmZ77IB89qBEMRh8nvXGZ
kdNdFnUotkPqqcwxsKBUvUcnOX+gOxQhbKr7V8YNAE5Y3QURzVTA2EO//B3SzR2k
lrUZhBs/4wxr4ARMohTeEwQBz0Pqiy8pf+/y51kSuY2SyYKuAaKbCzZCjywvFFop
oWcnbnR+EpLNjgQz/eJr2kviuZB7l78XgthEMrHcEoITHl6H/s6L7wPy6LvtIIF2
kqMglUKtCt50TVc1WJYchTQSk2PuAwI28HXCREV44wpKCl73lXTHPCqHYm6JMFTV
ctOXH5alvl2adEzk1O8SuzJHMj/8n+mfiERrWVwdpfNK6j4/dq/2M2m1s3c1i6XJ
J4NdL899oKA5BRma6acn+oTH0xWZVYAe8sLBkYGhfLysFmKqOEzmBPmAKVRT2idu
4LHq0imSraf314I/Qi07fMaZY1dmmHQrDWYBR9aT2zBjDjGgXtMySS2oGCPNgKGz
h1VHfdMwLupAZSZ5NuF1QSmRqRrlt2lQBf/WtAbutysHlXjRX3wqWOXJbQ8Kqk1R
FIyF1ijC1YzGdeE6fDrPHK6n5X1HyEJQI05j/Ba+yeXaKt9oKhwgHfJ8OYXzVr/e
CLnrB1Cn64hqEJsaLX762viAqP4o7mlGyPcvbMmNEL5Y9BT2g2G7AvGGt8y3m3uL
i8I8zJ07KBQ1E0nHi7qKfGqvyDM6dN/1CclDwmEyTxjP2CTcurEiT0DH8l+seYQQ
XX+ZDRy69W5/d5lmBAWQkyxgG6uM7EWpUAP6IGK4yZKEwE8tYWtsl/ymfEWXPh0/
veqa6D2rjeOrRq2f2affIu2TCb+86+K8GPJwu2hNEmDWzo2TwWki8ly7Ky42Mp+I
uU/zdVrWAAXAyL9HmHwgAWYqI+szHD8WsH/JYcgrBIEE+Wdtmcc1N+2qSKL7iMFJ
qb8CvifNaBw3KDHnsLjDs/ZTHpwfNH9oJJWQsuABUhGrMPLyrQkzc4rLZjTtzHv8
jR5xdEWP2r5Ss1EQny15kwYb2ulmtbXWgyRNlGGvudW4lOrXaWHExvnAWu9JI8ek
1hndQ5kxBKm3SNPvL4oHqz0f/OugNbNmM0N7luI5Bf2uvBXzkt4MJx1j1oo+oIm8
yMXTB+OtUntjsUhATxXW25GgT0vHm4MJczqdVEvqkyuv1qAQ4xhCt+zE0TAkVSt7
rabUd0Rf9KpYr4oOhrRvgBO3KMwf8F1l5JYLodAXA6IB9D5TISF6Tu8PKXPGMMxJ
n7qGB4xynYbweqnkFYueqyY83q2SWlrBaayuXA7FhZJjYCBDi7N9GSdmDHaXtvb0
iFc7YWmZbl+mq97SsGMdk8G/FjQtAQOQbP+eMCNW28ZHhjrRU2RkSZL8URON5kzy
S/VP0BB9neqC15dW4VJoOX05PjYqptjct6hrVTfWFkkhUiQpobyTiRRaUTNVQ1j0
KfWQVQjcDjldhR6GhbgLNLFLe4o04BioQXoJhbz5e+eRkYO4vCsFKIZuST5K11LF
63gD8AFEfBsCyPIIrMj/ZNIuedHCZxv2epUFi1coZuIuxSszX78mtTN2JLolIxLk
BWv3Scf6Eo1vqB1urzHd8K+scKPiyh4C1mKzjAq8j3Oh8UncHRPd9kLgjidl7AVQ
lnVfpdlvQw0kA9vJD5zlKkffzCpzsbm5oXEOnfiwVSi8tWVNvyFePBNN07ZEwXZX
xlZK0rCL9WBV4BeNXiAjdD/NkbrTLlsL0cCWNDXDdLQNNUCd2MPXX29UtrpvOdjT
4zWIFFpcAbQlKVGqVZH2gkdRnwGRqLMY/8e1XJ0lvRAQIkD6syGAAeH/jskCbilf
mJN6V6kU5kGVXUXoaTTA8sW1dU6AjNMqA6Tk1f9bikjNGuxVp9e3hOQVUFLYV97o
OESwPsYRnB30JJoEJzPwI8W0D7ZDYZbo3zHwZYJbrH7cwmPcHVtKurzGuS4DAdie
jxFmK2jWf/PiG9FN4bL1ISgHXwTJhtufVzrTkCyYglpx8KGncxguEmHGY0tsWzGT
GwrON3pZ8AtEip8hzfRNOAmKK9Vd4Efu0Yg0nMA1gmatRldzBsLQNeNEYZ3njnpu
q2yYv3jVQSKaVCNXpXOemHzEl6uvjR+BvSnbZcJKT+euuTdmWDfgTV2rW1FdLTd1
GaXepmQUozFLzfqQrT3EmUDRw3HBUIh3RZEiNRilpaLfQrhdtEJvHkC52NgtyC6/
kU5F/4zIxRSvfs/Wsa+AY6m5LROTWHuOuEPHMFrye8BlprjWWdOh88Ph1vaU3utk
VbkcQHxWRAOod5GHEbb8JTUxSDTWtS6QAYtgVOvTUv8X0fUFgVpvl7Ad5TZ5maR4
l9r1hiSWvidJ18j/RkovO2vtGqxu5sZ1th+QKE6rTzcTW7u1Q9vdmmsr9p+d/6/E
nUTlOVlUM4Y6eyj5nkwC3iY0kwdRwVskt4ZCMwrGnmFfdYgHdvDO9RWlXciHxd23
n0uP/v5E2Z+KGDQ/MTSH8HYspyTaVBvV/x+LPhb9XkfZaWhjEtGWL9Ovb3o0db6T
PdtAVBg/YnnHmpB1e6veKhceJFEkC+c8YH8j3oisUBxDWgHFLPtoHTvUW4W2cw8O
rjpU8PeP4OEKKtZZDeQbbIHy8T1sFuAb6K/xqTb2t4t6sTT8UaLtRY25HqIo2arT
IDrshqhaD0EVXSNHtZWD7jeanpd1qeACVYZ95D4uZqyXrY/Fl7gLFbJNRSnX5p25
lR+6a9wXnP9uNoMuMi7TikGz1AJruCa+2bLbPsn1kENwVdeulR15IozRmcZ9WFDc
c3rgOceuRB8RaIAJ5glfipjsWJp45Dy0AfXs7V0p6XbHwCkNHWb6aMxuTUFNcuQO
4g+q01enO7XbJx1MFazYv++1Nb0wZiLIA8sgoOaVf4lugNIqbLTxsKPhNF9H5obH
oTd5Jdzh0G1tEbNAU+ugQnz92Wae3n0A7SXwrbqGYaFt4yZ4Lv6GUmw2Y4l2bUPr
4Zbsd0aOO2+XgIOlQ5j8i1bHACz2Yrmx9Coy7IhpXIvhBD4KgEHi525I67u8wvdB
7X0O2qC063iWgMvWg/wVFLxFm+ieFTxhZaXhmUBf+//7ygodIIV/fxLTzDdMC+IL
eOAt0qsJDFYVOPCQDmrdj1ycy9TscAkxvIu/hvMhJCch8yUl+3yDd8eHRl5QH22b
I5pwr4cTKx00W9GT4wHpREsPrFajhvF8kd07mXYV/LfvDdki3FiHcKVe8TubgLDe
bBh8QEZpCMiHn8Tudlc9SjuRHD/hMt1CR8qiXRG5tX0G0WKJg4s/6KSGRiInDc7m
XQqptpaeoiKtXisF8D/0od2GE+9U92wU3enFjng7o5yA0Ho7QNA0QjLVegjSfq68
JpiZg7mW6YDdtxAEbFuG8ZeX4M9cZe7eJ6Gu7DAZChB4u8PH/HMo74L5Xk8tRrRk
0pyeHWg2nuAw1XTrYUTqoiEcoabT7dBRVAizGPB8E2YwdJ8bNc5NXWELt7atmIQN
hX8ZSp7JR8DhbdQ6gJYLgRzUWrckJFAL+sEYSTnGC9M1cWVppY7yJiYO0+UV5pf5
oYky1vBMjyukuiskSTNBORg6kMKBwfy5u7B9Uhr9WNRHVLIQB+H4HaMoXWKD1//W
bXTT1kuhUQGAnQsiT/nGKCydjXi11Bwz+u8/6bB3ifOKho/3J0ULDuugGOzGHxVF
qBOMyfoe5uiUvrx2eKmGt7JH0pMbh860bIc8T5LSMraOuIcTsbvXYS4vgT/MGTEl
e1QI84FvPs9s9iXzWPfOZiSzMaWND3WUL8R484yn+AvRgt6lA/jY5QOd10xfRyNU
7kfoZ/qlkU1RJD3HZZKmjfWTUhpgwep8Cp3N8SYInnIPsP2FMpweg1vhusNgQM5O
LP8Jm4R3Mmh/uxL7DTYlJZClKC0kN0tdLKTPan5aERBx/FxuxYeHHEc+i3k6HVEm
X4Qqt5AtGn5wJLQvmCRFx+YgTmPAqL6JF5PoypgZf1pZ4QAMBw7QHKvAPjymaY/t
TbbnaUSmaqISCaNuSqST5gaLQABXthSf2cnOpXEf0knx9AqwjPuKsxFGGfY2opPk
x9mYsJLrxRaYcR94nCZmhcRTjbgRfAEH5AgHj1g8OhEm+zVbjHUPWhhkhfgmHbTR
muOluPP3PVXJQcw2MbQzLXydK4k0V84fma9fu+pOPuH/PbBd9RRpQzBZ7U9STSun
jN1U/JuHX8XeeomtC3S2bvyiSJN2Wrp/GSGE43Wz3mKqRv/l70u/+Uy7F2iRgoRv
ghRyzHT8Ok0FMtxDuEboW3K2NNI56SvwDILitgDBd7lE/a+NUkbDphIkkeZJ/p2H
msRfDy/KIegkFgHkZD9NVJ5jhO8ISPNilQGZDOljgbrs6+n8DsmjwR8bvV/1NFJw
0BTRBI4MiheA2RKocKXLifmi+lm2/GUX7BmP8pmZ3eRI45DSFY+ak+vZZeCvHR7h
rLE4IfJwFySEIY7CFteh7w2qi1E44br83zv8uE99nOWuSb3ryId3L4izQX5Cy7KM
sWF/78TX+zc+yeoQSIv98UerhlTsZPLJednP1cRBaFvb+MsDZtsbWulbz6WL1IeQ
rcgdWAeNNKSCdCiPISwmbjWgafikLoi7J6jIMTJLAYT86UY61SxOjTw8jq0fJLSy
/W42TxDqqihZx1QBx9/S7mij5FLV6ZdUobgVjIdJrP9nTaL0kn/UL5Z6XF62PzDY
jh7I6Zaf0RU6zUkqivH6LqrO84tB4QphaxhRYh/DKl/Ff8ePuIK6uDY8IFTM4OcY
x5YfVTt7Qx1bgxAjJ9tVaU7q7OMJlt0yNmsBZtyWZsy9FoLaTbhPUFO7fB6GFUCG
bGi6T+Bs5y5tO22sENxedCEpT+zCrrHajE3MYM58Ua8PoA27Gokaks1xhTNEjhz0
xCOg2/y3EVL61XIwU0Mv9WzMFB0cpwk81xVmOOwNGb6MYcqPdSFnn04gJ9bMi669
XSY1Ekxxpyx1/ov1yWMz/Ccnojycy7WuhtDDcBaQRP+UuFIvT5weL3nCqFjaH0ru
qgxK88EZz4Ykk/X6vcUZWsTavdaWScjtwC4sNrvLEpFIPvTDMz2mT1eaPb5hPER2
+PTe8TTWWQBEBBVYvmeUQNFnwuN5iZGnApV3jBQNrl7n9a3tS+lsQzvoGKCmPboU
n92Ortyn3JFjwNrISasbo44LF/mnIXJM3QHc0104qUYsA8jhcDSLevqM6PGAzOXN
QgEi73QEhD7o+5qXWyzZtBXRsjUBjjAbYgCHgVyC0C9xuBCVElPFbkLPhhwwcM0A
DNz1SzGnWI6vJMSpV42sdoNToWDWYpUBKuELKHNvqtAF5SV8TEFzAgfi0aVgPsPw
cetF2FrrzFV0NdCPTzP+Fip333kq6GHPjZHFggXZq3fLVQdo5zMifZFWxvVeOJCT
cV0pZfRTC9gV4bC97+dw3oYYjuM3EO/BXYkN7o/AJRYdjN/rm8rv9i351qESOqNr
XAt+A6+iB9lNStVVY95vHR0kOhHd1viySBRX4Dz3OEcS4m9cG6MancJ2m/slIY6/
jdhgTeVMcthrGd5b9arZ1TiVFuwojJpRYXGcg6JUU74QlRGkutCDXAfZQAWmeNLI
+AK7oU72YAj0lSvzKV2ypwruDfiKKbo1DRV7DLK8242ZFRjUh7pi+2g8yEnMjdez
dPA93jzeNGJFQgVOkSHEL43AcSf8eRrlrz58RlcyectuJYfwAX7WrCmyJtiyGhnk
Xla+2xpbhJVVws8O4grxRUqRrqPyLRfTDz2cXdZEDRJH86rURM4wu8v1GVRs+pvS
6DWRrsRVT32QWnqJ4Vp7DHaeko8aw2W/UWv4DHrkHy3ppjAhJ0LCy+GFcvVKMrS/
vmD7Y6AHL2TbfqJNS1A4BFNPYtAQqBllhIpryG6tCTx3eU/YMFemzyRrvZt5sum9
qkzlDqojAR+g/NbEp6sufmOwDtcOcAqFsK79lkUWeV4r0dBzDPWDDEH/1lDSpAh6
DA8eLkdRT1GW5zpXWC3Zzozd0Aeway/RLXc8FNpHxS0/d11V5sRc5HJNBAqlcaWR
P2N1K3KA2+5sQjU1YIH1G3/1J/9it+uN3voNj+tJ/TUWXM+RsWIZQPkJubITMAsk
9jY7Tm5JIklG1VJ2UX1PV49XfKv5LuyJjBWsM99ZIgvTAcWQHTqtYtw0nMO6+gyJ
Uan84T41d15j6/ZFTh8rZPRdqHsXYyFhU0iq4OvCBxAiekIxwkUX94OyVRT4Oe7F
KWjO14gJn+FxARQJvg7eeJBz6QLa/0/xwrHcYoj+VtxOb2dsHGHguC1ey5tsM6s9
LB2ELia96TETjR66GXlkAx2hpsCa4pwpXpoPqruxacV2dCV7KgCG69h90prcAxZD
CoiZVHJfHpP4zTfLpOf1h0Waz5H6zCjiCBGB8ikIyQ/MEtEb3PZlJ/NhMCHDByQd
kvpKDap/GZXFIEpZxcicp4dDJtK7DYTOFNGGTzcyz+e1oWXEHt6K7IJcCmnWqS8K
nQHQfmwEabfoJtOChV3Gto7zSarcDj7xYWyoMfwPkNkrMeMVi0x0xhabQ1GQZ97v
StWxgyitZQrABOiuRRKA7//OuraK1BLmc87ABM2sp4offUk13vOOgLrT9aO5zSwX
bCeq1Ktze1lBdj5kfiLyvSwov7iTZ5kSXWyxNAvuVjDhSOaXaSnCgooPKKCKRNsJ
aO7/fYZUnB7OVkS0rbIznB8tyfpphkVsd8XB4wsKumbeAzdgY78df4woxF6d3yyI
Gb/0sFsepvaSDxbj4yQHAoY7AB3beaJhPYuGLMTOXzYUZSEFZEVLJg+E16KkDDSQ
0vWqyiffdGgQPJw5SYmWfwC5RaN44L4nIaAGgQhOD7W1HXvsiWZ1AhZ21Ngz19gp
mXrcmEKqS1u+EZTWokU8nqUWIYwP7FO0FM43S2MO9cfBg5cy81pq6UGg0tieWIkI
1kzMTbZ++ZLN99xgA5I4m4ZwfALblWLk3CYPIwWwh59cjLoJFVQGYQXo6gAzglOx
BGsiNGTP+srcRXilHbUyZ1jCNUYd47xOsvpxLOc09SjPVRDfZYu/BGxZBKa+/O2C
1nZefeOiyKRZbMJkRQWcoQ/kugAQ59OlBx8lPpVa5GsE/HOZhheH0OeMC1mm9eEX
6p9QwOdy1ZJh9ZdA9HtZHyKq4OxMVvQPhMIOqVegNRqUTuLs/dShr61JnSYIBE76
Xid1Oa/HjB06w39nntrqiYIkNmeHk5JrTFdTkQB4KFdCY1uw118tgCUVq2qW9UiO
wyk7qJaQ4XUGd1Q/VrEW9CTVPQ/H8VdinRkH3ZnHFzS/IAqqraOzd7PV2qAee8ke
sP+4lWgWk+0gfYpEKX5z+uIRgLP9prcedMmJhEkZTj6TMg+biKcCX2NtPIH3M9Bt
u3FjNgDcbQTxQaeZ7T15zu1JJbDwPowJbPqJ66tpOPJt8puUXg6Btyneh0R9LRF5
LQ4WBI8Y+pJUU55doC+CF06zugIkuMRKZLtkcIoJiqfSeF1VqM6MnZTK3ELd3wAi
3G5Y/Gi0Cg2PrKtJGkc1pXwhKmEpZSU33gHRz7dLLrX3IPhYgLd8F4fYS8HhrFjR
69C4eqg5JcW2FYyfj0uBV5x2OIGzGJMZUjzW3ZwMGKpSodV6c4z8OIinI3n+HWNc
xcJtIqpEfpX7x618ACkS8Z6XLgC1MKj5sICVqYegqD+NETf+uhHDWkWxjx6INVsv
nRbxxFazG98Dn652bUSK5PdFQepsJkYGQ2Fg4gGMN79HU5mHofB4blg5oAdODDOK
TbcoiV1+Zae7P6bIId0DGq6X0f66KL/4aBcaT9s98e1Zd7ip7EMN+72kVeYk8Zu0
2SLtEGDmu9KQk5MnPjZS17/HWa0Mc0CEGUrybjLTbD/aUk00iOPthEbw9ZJLZd/K
SB6kahC9qmKOhn7p7AoQdWO4uY0CQdlE3gvuBBQ7SPpQrNcbzfV8qvzzkfPWdM+H
rqXltNE1GyNL/UkzErz4U2XCPtBa8kvieHwCR+VH36SnVmWAj82Haptg3G3b9u97
vyGUG+RlhoFV1m9oAFYWPDRazi40tndcWGU57K8yQywr9v5Bw0hFdlgTsTpzyac8
TOuW/jzeeB5kNYh/P2zRtNlXFRo2T3uKWGUOCNIFvtdhAWR0gBNQKoT1v2wWwEbm
tQyYkhQSi6qBXEJzM6cYIiuFfUnDq4pQGwmAKcSH4uExYecouR/hvAYVRSOiQAem
VoAz4XXPRGRhTf5iyVnXtQJkgURMoi50aUFb5fuJw007QpIyYsB2GOC0AvBN61YW
E3Pnt9uLL4OGi0x+P4KFrZgtSsmOk5Hx/k8bN2p9CVg6fEznyMq2mPoYWcQdt88b
3XhObLeXOJeG/djN301xisHqnVcP+X/O5gDfrmhAiC4CErQkdD4/Zg6p6wf63dVA
cf0OpBDIxDgI6+zUD+XIDb/vSrS6vwOF34gd2h/PfPKWZz/qxGi7jmdkJwImLL3K
1B3HqOA0aPLf6l9hbMKihhcPCrk4PrqV2TxxbJ11QPUR2ei8nlu/nnyRdtfVbojV
1qL34yCSvsdEnyjW5HqLxflswBcNQzluq4OMSpLUGRoKDbYwVlTXTa8hF5RzeLxl
qJ89Bf9+5Gs4ciQmPBYFyCInL/h9PeRLJ5WNNx0ADegmDXuBSMjWmHFCkF7CeWcN
+qMtnoXyEZo6+Y4/pPFuy8IvtVxxCHT9ta+YUbamdeSDxh9z2bpvah8j3lVsiac9
uvctP7eIIpMNSnYAlXDtNI5/NqjJrvBoxWpOv71xD6SOUjMPOlwzEGJlfr/LSHxP
FAb0gzu1pOgFVIgoAFWUkjVRP0vrQMoHoaA9fDbkmALGRov8wgriEnNwkPIPDJWY
Yv9Z6XWeJ9vhNmtwiPKaoMkQ3dmQ6Rehb0KAkSsYz7VhgXdq+r7+3HzWBet7iCAy
1xhoCZi2wMSudhPoFQQfulDbxno6UXal0/QJDY4fcEZyoPD3gqympDdzm1tS6SF+
CD3ogMozD0PVXMPnDLcfzENafL8btu+QZrHjNZoJbFFCV+ASz/hAs1IkI/YBrbIn
J2zZ9yMjeTkHNn6oFcPTtw33jkqE6lK0IcX6LfqXkwNK1JkB77dsn3PtZAsobhcD
1SFJFFWT8XeezgX02mQJFgmqt6zTxnP8IES3rGCtrp/0pUHL6BVHcmaL35JPZrU2
LBJSQnsuiHiZ2cDJhVIFsJzCWseouF/xfEASB4u4Q/qVG16Fmeta6xru5VfcYVAV
D4foFxrRAvnfFZpQF3mz1VaRxGZoLQzd5CyiO0fjgoPp5WiF9wJJHeBQ4n1v3v4t
JZIvAPlfR/R6ia47yaM4sr+X9JsHNgBKWfGh9Lkpb3giByDU0W+iKVPYGegsao2o
t40M4rEQDziG/LofOZ7xdHnVOYfwseKtjDMzcW2EVJFYawpJ4q9lRhX+laoLdpWe
jULOo6zD57b1xkYIDR4CkdSryDimDWmK3WifS3zRVG2FUppf8U1K29KXR3OZ6waZ
cz3ww8LV9/lP7M+IBxfQlVB2uWrMZNXefY6t6W9CZGtMSeFQyDepXOTSzTNbQpxC
W4cU7dr/iUFbO8vqTn2EVPLp5DHo8EQUnw+QRpJJqfUfUP1zAH2EPPradpn9Qbgd
H4Y8UH0Di9I1xauDKFTEPNbOyQlz/LXTsAoIpLmv4GWL6I5Y04TJB32jPjnWKNcG
QFO25eumXxHn+LOqLyKVfOoM/5mLhCjSL1EErKkx2bp1TEeMTWEIeWn0Xq8kEVNO
371GzAn8tlZSjUBdkBpiGzsNcT6kWdKbRqPwRFDbvv4gidE+BswC8hgxAnCesJif
8YSaLzlSlCn3fbggdCTrr85ekUgKIiXDGv0Q/BePyogpaizvNAM5MqIOQ8pje0C1
/nm2hmtu4KOUEij/IbLEFAodE6rCQ276kkyKMZpnVRNrBpFMi0EPcfbYNP/5MJ/t
EmfYgOZBS/uXIeCumrJ88CMcz+4yBh+EjdaQ2yInRlZHVWzQFj6uBt//j62Nkryj
/Zu0h832+fHO4JG1ePKh5cvTYh/d9BIm4HqvP0e4ZhAgsOCm8UhDsyjjJdEi5x+P
p6s6QP9gZHIZIyJi5ki/HmNjtmMGOaezolLn8ofO9MGQe01rDimJ6gSYoGS3jNDl
ZiRtQ0/aPTWawWac+NpzQvkS4oDX1D5D11e4A237+y0=
`protect end_protected