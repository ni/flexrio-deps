`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFTH0lSaedAGrYi1rCPd+iJ8bjr/R1hcOl+Hl2U5Yvzkh
4ohiBG160zadTw+Watg9lamx+TakjPN0Dpuk1GvKqP/x2pyX4M2UwUiGgL4H6/KZ
zDAzK8OAqR2pfjnqa6Zxty8mM/xArz0+spVXs87osnQeOgOdfEeDITrrnduPsCoa
zhkUYrLHyeZtUhInKj0QqfIWACv2Sinv1P2ngfOn3mLQlOSwm+DhRsRhkKJCdMg7
edLP5ZmycChec0XzzYAyg72en+s/aXVMbxgY6zi2E8UCYPRYeSQ1wU0+xxTwn/pa
USDYRw3OS0NIwCyzUFjX8KiQZmc6nxYMaPhITOuHXSrM9cbnWqoICP25r+batQoc
iSrjIfovJUfugPVdM36ekSvGIG+7g7JLHmDCzGU98Kkiqry1NFgD09o7HZhtZARZ
8iNVUWK1EgQFTKn9yIDxvR/ypCsbj+6hOZpz+ta5l6D1D9UEp7qcwumMyk/FA4E9
WYYMIEVdt2aJ5cxMVcLI5lNJrLT/v+p7v0dFVKFnvm4hHDlQQCRHc9Qv5mN3Lz7+
PL7+OIoi61HhHqXFL/Ru9XhkUkIkLtaVKtJlpN3iuo5sBqGuD64qDolzepXiEuKe
l5gwL4J0J+ZhGuS8JkWsjLIT9RsNPWeMoMXEWt7fEB5y82toyRD5vXcBQ0iJ2SLJ
X9jx7IrvCe2GuXgQB3Cwd+38NzgVLkogf/sSOf9j4TDH2gxcz0YghA/lRirYJkhi
LFD27GjJAWxev9pxfTLDRjlFc7wlrIkM0OL3ctUMvY4kQEgKsj5abn1eRFH80vsT
ZuHawlVCZ2n6kZjuSG0yaqaIgIDwJg3vZLY7y6bCABx6sxVy+hOME817F5zU/9IG
EHsTXy/95rZ2FY+NxNdZjl9JJdCS+SGUu6agv9DF6x38UyErp1d0olDqARI2B9ua
dyar1KcQzBKviYzI9VkE+kADdc7LlZ/IK6q7JXg50uJzbtAUtMDFzsNAUnUUWt+0
2oZWJyLr4V6WKlidxCNQX/y5r3RJ3SsL8R3Ycew9C/QqYr1b3gnYi5BYy6R89KWI
1m87XBj786zNuHy0lShkeEDfoieuZeDnZah5zBirCsOxm6NMuVZJQx1+wky1NIsD
fxa9Bx9NDEw0506hyOqb3LJ+ksdJSd5tRmk7WiDrfgBctAPmoJmEd+2BmMeR3o+y
FbiKgLf1qmOiD2TsgVGYVjo3SS3MiVq0S2VuvZjwIFqCA8eV0VafGkys6ba35amO
w2oKCCahI4CzRxqGqWltgW3IkxxUzhirvXutC1+oSwIUS7whjBOBjrLhIfWzbCT2
XkGajN/3hB/WMtlmRQLlzbekAHMoXqqkD9iq+w8IEetc5if5GVcKtA2azkbtGOae
KY60iqjTEUg7+hfXxYM3Dh504ALwTaxiVuUHh8yGdJ6Ekex/8nwmtFPi6jx/BKd7
gBPhc+gYel9aRafQp63PZeK4SGVLeFufdmjwEDs2psMXDmdFWeE03BHnnOlPQfGh
wv/HX9+s8b/Onbs6UDcigZrv4sJuB0rq9sJSc68f51USM6ZOhBMwdlWWsXJdIZ48
LuecAefaqLaID6uRw+IEovHzhLjoM/quV/BI+SlfIep1P6P7wlG76V8GrORbSWT4
v/m3gr0HzfDb4GOcmv9d5L5dQotFjkgV5WwMVQ/xjCDzTQpn8M7hg0KVQzcclItu
iE3gXo8xd+jIopewe6NfBOcJBndArb7rOmcirurXY6+an5xDQ4w12yAJIzctAf+V
jPxD+RMSycZyOOayf07VGMG+j7yGgb3NjctpMo6eEDVjAC4sTgINs6vIaO+RXgaY
HXKJ1QDVRYlWkdX0r9QC2VwfRWzVQRwaXt7/a5ixiQwcMO5yGeT+iMLfN4SjFers
CEqU96gzWDT4C1AbvmDjeNc9oH1rwUx971ljmxAP/Y02rNiMYtAtBYBQtKy39DQW
6m3Qvs0JAm5A0sxXz+eXIxYFi8j3uY8+htN7wF3TWr3/bhYbeYuKB5me+r7BQKLw
15Tkjxlh0Ncurm+nU8eplGxcxJbzYhsIB3v5xMc4udZSXdC9n8J/9ya+W0j4M6kh
DS/V/n1cfSPNxwdukzJLkxVX/XLZKNuVoc7vqxzyLrbydllq/QeTLi6M92ZSEXmE
QBrwPhR+RpgIRmgX+OCaD0Y60kNbuE56McYUBkzhWuEom2D++CXJEinPns5XfKS8
8N2HOsq8Fzkm2ZzxuGXYZRZFdYB5szhzq6yRzRr1nvemH2vrbOYGjokuabI2rLP9
O4o3OGsRqk4qIcSr61MeJLi3w14R+YJ99+9MVUewYlu3ya1jc7ULZ9k69bSOhfjO
IequwkpuNT6timT5WBEOUcYvAA+o06HKqhoi1VF4UtSjV/iCe2eGQmPm8A4Uk4BI
TDi/rD8tfGDNIGkLelbnC46M7IVWoZQOmg6ptM2eZlrCF/NyhmPZX+aAcg+Lbx+O
BsjIgGm/9gzqvhOGfL58+DGEB6wHwfX4Y/SKESN1gXX4bH9pBcjy8T+EVJHhG7Ar
GYaINIzPwM0zOHOS/2YkG3MKR81k/wrfktcFVhT1ib0VQh3/On2oj8vsGdDtOoeZ
fbgh4/X/XS7bq+Nf22NDkDKUNlCrEK1puUKixOJp2C23pGpFOR+XB2VY3rP/n7CG
gPYxia8b0lrDs3rnf09RHNJ0LolJ7OvKYcYPu5mcF2U6bagyCJ5P94ivHajsNn5y
7l6pN63g0Z6Crag/rJelAkurbFaxzpg8cFvFE81kG0NY0dKQ1+VemnMdIdYXiNA1
nww1T7g+RlKNQwnAnOMOfuL4Po32vWcJW6G/1/mwYtlwGaRxUIawDELAI0fGusHz
tkxgqYzx5Jxg8hCwiQc2PjQDaKa0y6mXZC39gL0qiu4IiBjMV8vRKCtoO2fQne9B
SIqFX93bVAZT3v1oZEzJUk+G3Z9KBKB5Ph/IQO/OsD9OH9NxQbFHw8dbuElw3Dmp
n2h0ZgjIimFTgk/8t+MmiRimfpY7viS49+LzDAiozSWsQ4paq3o90z7CXOAHl2Te
IaQXtvcSTza+gg6mMN9mLzFin65z6M4CzzhvugXgtMPI2p7MZ0/03dIBJgKYpMSn
zcMm21D0iNpuBCdKTjsBoknUqF25XXaXw2lypPjbrf430X652+96W14bykqOPH5J
Tb6zgqKw1kA3wo1OV/vrHYY1maDs2cfHYjfTtP1KPZE6vn55cyiMoEueA3KKmNba
8K/BbNXF59KHFrm+sAejFJJ7WkDm5xZYxGftWo1FoOE7YtI2kH3cu9MEyUbMmIc1
apUwLGTL6oUly0q8IaxpN2C0eQXXy1BWACKyLy8lgtERh3The8QdOXzyqqRU24aH
cKtpgnpv5ge1NMF4azoM4r8s3ZP0QW5XXJ8S2BP8SWQwDoj12S5f6JPnJlSWVc7Z
5bd5R63e9LRNv/tD4Onq2jem7x7pcIRSL9Qu8qfgEywYx+rqm8Lr7I4k3OL/7cea
2SiOeqEgxSH7+DA33rO61aRJwisQqnzqMGFuPzq/OWfhpJvpeSinBCbMFwPo91PD
P1dTS3ubUiU8jeIE8hThaJYroK+6niB2Jstl2DSDbO7BhHhGRWKaU9r0tURhtiCC
IFl+m25Vopcp4mDljERUO/mv6nfPpjPYB1KNN0aVZtaOqb70dDeNYxhjVtcoN/6o
ArC5Zjm6snQpTE000LSp9vG2Owk+Q6GlxevDu8q1N7KxZuzeeqpor1G6+Tu9Fitm
2sQDwNCiZaCgZYqpHd3eSJ4YuRjDQqGZat2fE1junDoXNygAL5+QzKtV6woevJWx
DbpwyJqLVtLK0F7qnLSMg/ZKULo/DthsWs2UAL5UG6rMW7SmTcufHAc3741bsCGl
WMAOU4YL4RPTy9/JqryvNJaiRNd8zX2oQrBI4yaE/AxXw/fqLNtQALtFu/E0LmEM
WYEoSnirm0F6uQXbqiNK+KVYTN9DLSJ/u3PWFIzvFoZfD10tboW7qvE9jFhWxWHq
KIrAUV8Br31PpE47oYmHMwT0zZx2z9uMcG3ur7laU8j5TC03N5nLLSQJ0yaSO/9o
AjM37t1/odDrxxfCPDNwYdH3F19b2lKE2f2PbJ9Mot7JV6bmTvXi4oOULMPbsIxo
k/0OIJURD+IV4WOlWHDQnHCzn0EZD3AMFOvCBFb+24RpXxfjVjp3lGlyVKjI+zDP
Wv27f50TinaymLNKR31RxfgWRp+VnYbAFSMiBD3pgJ8aIbeTy5iYjbokglnzmv5v
L+xROL3NI+0eHfteBjf6t+pxncxANHxr+xOz6OxzX5Vwc6TnPx0rjvABTXSTY71N
b1neXKmlygrfE+UfmoT9Q8/HBQC/QZlYzRkQT/DHUF7D2XXzLJDb9qz/oNyukHhc
ZcC/L1WdlODCw6/2otOWojUqY3sDSUcdhuVuc95ioKK9WFq6KurcaT/4a7QbEIKF
sbYmpJp1daUep2nUL0SUtyDVrQEsfrt+Tct6suB6sYO8LR7dspYxF5GLnsmK84c4
+KXKV4bakVmx3IKfmRFfBNSP8EmwSD2yFJtTYaktG0bbb7BkeOcfJYqwJxmdodCg
i1KhubvmSBGwEP1zY3p4Ju1qTu3M2Q61l3QqorMMauS0WMtHzQquxPnOfvlUFSlj
7v7XjJM52blwcKyBE3Kzf5nH8yPTRucce75/uhIrC7GWl+rJT77GB3zvliBgDxpQ
nxS08SwKbugEOaiewzUS/rX61uzkT0wvLaY3uRugBHqtyVLvkoFZe9hpX6kdH7/U
KC3dy9cKL3cGEFTkFpU7xAKCo5vv9Rdq70DEalBm85WfGvWXdL9977MprC9p7Fk9
C1+Ls1yLtGFGrg49h4eWQC+Ok6vWPVA4Gg5WnumlG33ZSMWDGqgAscH5jF6YyoyG
zUppzginDgZew6Qs6u5I8QpAEHFYeJUw5nSGZwH9+h9XeAfjeZva8gIpfFunO4q7
0Hi6LOBqPC6NjOBk6PaEfKx9rGYMnRjqC1p/tultOThbU33MTjkq5tarsr3fbRi3
WfziwUoBbQdP8onM6LJljLufteobZj8tRtwyL8eqK6ZqoKAWGpcGuA24FpEQFtTN
9i7TRo7AcBNG7SpJ5CoVKPXvIvByJavxZM1hvXl9w8n2yXSusUHacArfVN8imWIR
6U0kk7b+DlADjTTjJH1zTKsPFC2IlzCK6sVI1u7MVRHBGUuC6NMWTQLzj5ZVodWf
ZFTxzWZFLufkiP7pXCQAPFJY+9bthRLkZNtiV9xZat1xBWathTmbIi1jsH8NAMJs
bBvcdx+V+DAsT7+GEDSoIrK/HZZIfZxqBOLjwVmsK3aoHhvn2naskumEEu0sivKV
/OH/W2hStVGyNeQERJdYl1rC7ZO84HUgEkyc1iQ9c+es1DWWfoSYa3PsD7vU2Rk7
1ToCFV+SMA11TS5AxwP9JRzmN5ohSm4miwhIjri8FhYe03OLWVuITjI2+i9sQOwK
yczy9G2NAXMkAOcYz1kH/1X2wQ4/ctsKpeqgwkiR4fcEBqyADFAO6BeWSG6cmsI7
Cq/GJJ1geh5nBNVpOgu6Gu+8UENKycGTsajCMWqjI1liNrVFaIo5rZC3dMqjUspX
GDXAISZi5HhkrZv0EhV7q1zJ5Mg780r8DGkPzPAEV1UpRnlpuj9gLpXTdz931lbY
bfXcQmEccJX6RE8cmHB5E7DFrORL1ARThOQzbJQOXeFHYpNSTPIQLTg7bh8k0+fj
s585XOjxkAq0CUuCQ73/Jin8RIwD+FxZ+Zx/H1DWTkJjII6sz+9KJS99MvffvvvS
DZSthxkvR+XPdvaQ1YrCAEB6yeu1rfuiJBkF6hjHpATpFBQVSqRQJkDg7zKdtbtC
xLCqdxYG2QdvfMOZnh5emfjkSkw/kPO/gyza57nYhzN5apZrLSz1xIqzded0F5V+
+IA5wkJ0RtnVc/okpNYy1vixpeIfBbayjXfyVI84ReHfk7V2prH/KcrcBvWvwYOE
OWPQy+ygoScuhZ06Ev0M9dl5vb/kkESjgmXqzjequoP5RY8ihEkX4/V5uheeqFHE
ssZxJXHwJKqbcqT/s5O9QqFYDyBbSDSpBfPjltPaWXCa1uCWNOXGfIya8MlwCac9
BW9wyCm/ZPQyldEIFnpMlefEaSTpXTWtlkEVrvpR2Laxu8/OYkQRMhnIvrrjvFC4
/lqeKTH32/w5LeHEzBRMEmmggIHYE3XHJZmz4I0WgCYcY4IinGTb4mLx/yaWkSWQ
/AM3073wzbziBrDpNvacxrYVce6Tlen05oGNenRAmktSlviZGt0QLhoPBE6YtjCC
GHm9e9trqW0V8iuuOiHGF92MlyByEt1zCPRM52czyd8FUW87O1R6GhV5EQ+okD0K
+I/DshvBoaokK8RyBzUakQU0mIv8OmWBEPUyA1GlGvQBa4H7pZermuDstJeYAETj
IS6f9zvsticoWwa/7p0MB/n/E7A43Lp+jl4/RSNWftru8pjZXlay0XtICEBwv/ry
bsvtYihSh19B7swET82fCMxIBA6RdAK4rh9d32AfQqc3TiBRGb1Jeo1433OOk5TM
bXOuJXonTjwfkuYhW0epEcVLS8u3pYsClj8ne5vssBJpKJAQxzgE4UtNRymGO3pT
8Jp/i3s6suWzUpftfzUWtiM+fs17lp6d52zKXuGXk5A9Ux+xietie5Srml4y8o02
wjas8fGQwT+1dGn0CSpIRAOGgtEQo9PIF7yJvQXtCu38AHhEl0jJ6UMSKhJn6oQ3
o8rWNdObffAGE2/IWcQCL81pscQ/9EEHpGVHBzGLWrd8OZvX0gs7hbWNCFEdH+L2
j3y5laTfMEgLV5UOxOkHr8yEr6CRyKn1ZQ8Qg+Jtqg0Jyp/DMIzrx3DH6JNoDguG
Y/gcEHr1UeFbA7zVlYkZxmTn/Itu0dGOl+kInyShTPsmRQPeaR09wmR5uJ0S2CmK
jaqb9NzwhPLuz818YlVUOxu7gwmpDrGdnyNaDExCkCl0d530aaJ/+gczQXCB0h7i
T8QSk12w/XIHfdPUrGbWjPe6JpvWFJiG8rp7ouDxbMHjBi5PEYGCqrd1JbyleaHl
2fwvOLUGt2O2b0T2PPZtWiid/P8CgOq5dMm3jFmAuI3UijHJjNmaVPAM71sRXaAx
+Qo0MAE4PTs3SY5p3G5+nPsWSf1pdC/A/g4f3OEPksKCtwReAkKVIUNMlw17s2us
jP1b/+ojBEyy/iwZGKgFTd9x86r/F/n7wycXoiHyQcpzIdmmMbXxrB5+yqjNgfwk
3FOzPmTwylhWOqRenRUGBEUKfM9nI55Gbn/lxrnTY5kw8snpp29YPwhdmyY0n4iS
rdaxQHwHoPwmY2TjyS+yUTcqyN1URglwbAU0Gz14AzwuRLi7vtb/C0f965m25tBW
uB9Rphug1+IrvYrOBduB6GTXZMuhRhz5d/Fj8FXCqPAnSTIZFlB5T5IHpALd7xni
NLULFUABGMNkMdE/mc4BzA/Q0cvy3mjJR22NGOONcp4nhH1eobMPdy5fMYzT8A0O
E8tQUtyIecF/Qa1dR+2yYsmJZUaljF5Z/CXJWwyW6qL9NNXYLi2oeHz2oSflPWXz
xhQOLe9R4a8U7mW2+xs2hrf5MFMTJ+yCxFe0twwAd8Imn0gusBen0qhOThiw9+B9
j5XTScwWOWzAGHBlVXQmB5GXyj66925Oop1PEFs95Hm/EAgMlAbImzhsSWeQKHmV
CXQEncyt7tY22A9JXrihuLdRtYR3W1B25jfEb7kbTkCX/nmtuAzFmByWYm6TYmnR
mJgD+0bfA8hd05lS7yq5aw/mbyPIglr9YF2k0oH+HaJmlSWYT10Wc1GjuK4pAocW
BqvE5B5p8xH6sRPkL9ENqMl0bC+HITTWKM5mp7FDOrsAEyU3TcK1bU15tRalYhTd
NelqjAs4s/aP2SgKTLmbXbrv5M47oPrdUwjt8OSy4D2AH5oVbdknb2iSlXjsYnuu
qGFvaCBQdjv/mppCdiXuHiPK4Q08awjdmBDF2l/9SnhKpnxeQ4HmvHAGw/JMloi+
kjaqRUoBSi7gLflEjdiGznRJCA7dlPeTQw2aGldJMLjI+HW0VoF4VuDLc7G2QIIp
HjFVBr+3YGGaTCnD4ofxqdKir37fkggP+OsbuGNma2LUqYYdU3hHuvfiCfnUQgWl
KqmEUKF+YLx+qBl0/pnYeAD9AwUrjaN3mFSawcDe5zwJ9Y2MrPVCVQoStbamKWOR
K9JOHI0NrV2nEnVLBGFVM/nf+YKWpDFEcvt1Csqr+DKfsmk3vBPg0zp+kcTEVFX9
MsuN2ObD5xkdAfZdG72pDLkRpJ4q34ceKQGPxKVDMTBAKYZo8gvUQWK5Pc+sxeZH
1gET40r/Blj41D+KsvjXVXpMybbZ/w30q1/ObuPntPxcCWcwkcXgu60Bs1QFinxR
kB6j+41hRU0QOZnKXy9w/7RuvqAZh5VEzQVwzdX4vYNDXPabTwB1MemouLOLw02C
io7MZxoNCEMDkebi7iFFag==
`protect end_protected