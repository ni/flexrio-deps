`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvc7d9OZOUYv/Ydd2jVhg5pw1Oky4yTg+qWvwQ+XIU1H
QVFP5lLKmhTinCRRqZj1bILLg9pxKJJpLO3rrIuAdaP98xTy6zOyNt6Eu93KKEfU
zkwsPMi70wePELRuhEeCQcnOLy3LWqkRdwguQs23JBxNAdy1hHs/Cmeb54yLZLI4
UHGBaCI+N30EtREpUgIhmrgIX2SrDplLwTxPcu+xEN4lhTlE2PbZM05H/jJUy+7G
+L9HB17mTAxW32G2UsC6qO6nerNL/PT5uu40DOrJZMWtRy2ZOAnskMovBC0yOeqY
QQqFr3dXk2MubtL33IaI9zQmnNcjVt6zjo0mRmTYimb9QRXjW2zx/V/3X1Y4lWgb
nfjcWbahIcWLORY7RH45hfCVL42ITkY3xE2RRcsMoKt/dpFiUavUhqaJ53ZyVjCW
4M17EsDPZNWIzevlAQHmQYQJ0Pm1AyHAnRQTONT9uXk6UV9R7QDByktyZS7aYsNp
G6CzsfneX78mDJk435aYhd4OJuCz9Z57cedw6XWmXECxta1exr7Y7p4Spz9NVQBA
wNuEL4cnmUNliDapYmej58M8FBMlI/8FwSGJjCO2cnnmvsbkeN+df5c7RskNEgBq
P5zA3/Sx9Kd31yq57CNrjzO9NUHhnxOainyssNa7M4UkBMGRTdSZJWKWlZ9T77Cp
yc6neN/OMIJSuOvwAWO6kzEE1tWMwy8mFKqe3UZhjWXkxO1USTAwKID7MgkIWhr8
xJNf6O+odH1itD0QVoCA2QJvCswIG1PenBBH21xOIGv3ELDPIeqs2J9S80mRhwpW
Usl+c6XKmfOysnCwXyxe9vE5pqxQ118UGSA8cGOYSOHUWpWUWBO+Buurznf9yvmU
YRgwqY2b+EcrLv+m6dDcrK07GHdDyPYl1b1TFK0Xf24dlael88taYaZ6VS6KEXFe
/m/naAGq0PgeBZBt6i4zngbkWTZXSZBw5BNNrbLQY2MZNnPSZCy6jAcLANYbA89V
dDpVDt5cfYeNe9iFyvqp9Gxu0s357zq6wJ3DtrdMe0xTSnRS0L53E6De9iyjg+vT
dJh86MMSQcBVMLyaHHduVvZizCoqtcY/szaawPu4FnfQQTJNO/2WWdAH5fa7X21f
I3Tt5bEU9+QymxXq4jqFXPnh8fO+QPebdLdpjfADtnrTXZFbETKxLAcYmODzdgE9
5IMZKia97IT70ZLZ2TZGIOipKIKD5rDeWlnLEcA7mWciTmngiIXq3EkLQhzHbIke
VxPOgSSjaTxN/vmKCgf759Q52Wh1RMV/J1r4QYdRax63UMZyQQltzDwGHol8xtzh
awTjiCr0jgqEaw0DALodC6gcS8pKYG09DF55fXUkJCimh7+f+hr1fRI1XE/bmimS
VAT25Yc1YkfEULQCzUVkxnlWrBXsSZb7UDP9D+JbL2xoveWvr5671GXkXT64KBzQ
wxqTW23+PGvg+Wn8mMqKDpNJISEAOH2JeOcbu23iuZrzgvJizntfMmejzibf+kDz
NpSJHhEDl5oEiSEyAoWFyjIKb0oQsYaFwRqcxOJxcSaRVvdgk7LY299AqLbykgS0
Jm1MJPzd97UJgyws+D9VfKVVnopqF+ga7/l36UuYjyN1k0FuPJRRgnIC6msrrRnw
oDCcpBieBM7WMC9SiEASs5X5PyXfy0F1IW8sHJ3iR6XKD5H6h6KpozZfdsGTVlzq
rC8T/7f2RkZe4z8VplGaEuYiTiFRB0Q3G/UvzK7D2TgrgSaQWsXyLTHzSqwNpYUB
hrmnJAGGp3V1/ux5UEJRYtXDdwXIVqRn2ZD2CA4c9nllYvSiqGhx29hGJdg22A1z
TculoBmAXAQbkFDoQ2ba3t2kWskFZRSaDsb5lsKdk/HqCaxRJZW279U5wOmuDDA3
tX/pLrv8CuXOcQ6qTvvfeVQRQaz+kvSkhDHWkqY7EepPWN+I5jm3Lm2HVncuJXD/
QO57PQBn7Le66nmEBt6kwHnp2IcnvlDVmjOLjwqD2/QXHIJmhQhSg5glyTH+wp3N
bQBG+eqcVucvTgv8jPuRAZBQ22L6ieHmPTPheGPoCH3TuB/U7dWGMyIwGyLQkZ7c
CPCeP03GtaJKytbDgNPV0jiQHUEfiYXvy4BEdEaeWzYoWw7E6ElzHlxa6MQd7baQ
mP+qDyFGPUdoH+plW33QkkXMX5dWUQjVhtNy5J+xY0jSZ5+gSFLEUrMpbQIQtyxE
2TBCSR0Fn+0ncpr2JKytDVB2XJ1HzUTCSdlSrc56vCz87vM6D13g3kYpM1/16apQ
OudD7ZcyAtOmRAQCvEk+MDkdDcuqGDLNCaP08LmkPVEhWzy275gcv2Cf21opYjmP
zebkZTrhbzztlbPXsmL7JzGCFP9rg3TxvktCIWb7ETmUVK2T2ySR4JiT9UGcgK/x
hFnakgCROjwljjmVSGcf+2eM/LvRpUN2Ryn5ZU6jtM6tS6j1OXVFxo4LQSSIadYd
1wEohAfZotkvlH74u9ilJ5xwOOYD6nG/7xr59zMT66tKk4F1vjok9bbML1t/W7qy
oOr2twBFLMGilX/yYLXMbw/VgPoBiVsilCjoLnZUQl1cHvtOLi0aiNm25FZu70o2
AzEwanpgN9fJcKTCihulN1/cRXtT+tX+FlApSZ5oYsbDdNF8nDpc+cY15hjVepX1
1T7YPhHeT39RFdYxfrZ/NHB8CabBANfy7slpBPiTwIvvTOZQiQiYSSgNq+eJ6BJ4
4QqieNRYqIt221DA0hdW7p4Wzo1oo7+6ZUIarAfTSoo4dlW+Bzj9vAv1Q+h3qBzX
kzitpq5uxmn0rFV2kPXwbV+nQludPkIUgnuSNGuK/S0KYQSdc/Q8luQPyzQaCntF
r4KyNqrl1Tow4aI1ALWBOXO+xeH//JUPCyevicSp5/drrZ/OwZpum7ZOvzZIJmqk
msWpqPGqPaUYTPw+HIZm1g4ciIAeDB23BlZJtAGAs9zZT0DZtCMa2sMM1XUgRmPQ
C3/LLlZSbHlsIgVA00Em61ggImaz2JDJe6v6noQ7r/Vb1MciCnFcJ2JdLlnX3m4j
8FOt+JSon8OixG5Z5qtiImHFY4/zVQ4wHfIbkHFwcgblgx9BXWoI5F9aToiIURax
AQOwBH+iKC6r9U+GoQxTiTuW3UhZfFFnlC4SqbAn6R70/HY+i1yOC5VThbCZZca1
UbB2fMkvjEFPq+as0QoBu04ldfthFFbOvTFEwqYzeVAjXiZYnpfIRpYUqNigJ6I2
4teCk4HqOZEROEy/y/IIl1lm/EKiaa8Wvhhyb9jrpejF+4/iR3eIjb6a4KK81pO+
mbOgsQCOuozoevetPYVFvjG9LDzaxYpo1YW1x9rgxB0o3JFnZk8SJvqW6Bk+TRns
Ls19Tbcelkn/huB+Psrl3jGxo+/V4bh3P+qyiZhdJpDqrfXjR3uwk663/87aAJ1Z
1kpdfVhGb1dOe6l8fQ34NXqRek4yi1sLNgj37WegCkpnj+ZEPFooHbSGW835+73n
9P6seM/lb+09BZFbIOLKsfyLK2AfdNfJFapk3UDV+pDdoKkLzzEFCAK5GbD9OY5b
SnaJBT35C3IeW3wHdMShp6h8y+r3PmYCUssL4KoDpvZr9yMF6LmqwoxLdZ3EVME6
9qptDKfvYgF999uY1hqHuQiMN50MC53KZqFZIoOuSxkQtU+qoySmb77ZFCA/4cce
ZR1g61lhfgs3E6JBfWfTmlYfFMythFVTbqvet0Nv4deiHc9e1Xvqlj8UJvnyETad
dT6qEFx0jCJJ4cQPssVrpxjqsAux8EGxHqq2eenY+N52xdq+PrNOUX1jPNmjujPf
1qeCZ/Uw0CXnJOcDg8rDYGR+p8OmAEs+8rlo423yZomItDmPvYJ6lVUD8QFUoV8b
jqoup2BQP73E7gfdmkAS53Cgintu6TuwkXY5JzdEHCdTK6VglsBk7Q2IAKaoUaLG
h06W54ujPxD2B1NT5T1GEvjFjcFPq9++MNzbN4ALdSoqKIMJEJCxiU2b+fNbQvvK
5lS13woMZUswtu8w/UlnObUjU3CZXAcJIVL/3QuAnYcYKQ6x/j1aczvAQYOQxltu
X9fKmQ7IuR7YSk7I/iy8GqVZuaHyKEQSU6sQwg2kf2iSv39n2b21f8vs/lRDXad3
25x0M2D0cim7z9eS8VEAK8DaFfuGfEF6pDjMD+QkF78fsqgZ68c5N/L3GWlMgxWk
V2zIkHchuhnQjVauf6j6dRamyrZiNJOiEYsboCrZV84VCXUg1EyFm6QdOL4/q409
NSREPE+gMBvUT5NSb4haaCD0yfwynaA50tVRXV/AQyNCKYNNWSj8o2Dd7JIHkZo+
v6l6xrIJ+XELphz522XDCa/JNrNivrrCwBCAuz6CEB9Xr7WVzgLsnWnczthTGvQC
kKb6yZ/qx0eJNRkY2xP75eWgFAwGhGmNJFzFyUi/ZfKveWr9zDZugf0h4oFNdY8f
La2NhAqhiKsisu271KTbO++z5VLjLHRJ3pk93aqLvoDmBVII1HA5sIZEH6lWOF+J
LOMS6HJwvzFafaqbCzKmd3lFk6beOIBMPYBfDi1cTRuFaMbaOJi5MwAwTjb8ypTn
5q/yJlHuzQpiEVkXC7nYHOv6oCykMged/gBlacliRs3ZzUzxOWNTleFUMn0ZgAvG
oh8wdqEt/pXyQNFZo4i3iiJWW/U2fgEQsSgcxgJfkiGSCGMWNO0xJLdclZlds7cE
HbQTr5ck3HVLfqT6MezY2Gagqtc6AOxRcM5IYonEdiGMKxEnd9ppL9uk8mDSUzVP
Hs1/ZdXvxbC99v46GbhLBAESBAD3wTXFmxjwTNJ7aRQjEJ9qmjiv7DZ5+1NQ6zRI
9rXx1mMPsnu1HntHEWej6d7RjSALGcdWF/q6HT8ZznXAarXxnM/gpG6bsaEJ1u0k
j5yahpOJ6/7pCkCKDsPLnrFSU/3LfPj1BSpHoRwTIq7h5UIVhKq9Yxc4SwLkAbia
fuZx0/pTpyXJUfgSV3v1nhBaNtx6Wj+xqzwZXZP63sm+Jv3MBgTPT20yMYjBycFV
E/RasVYx+VJmBaARTB3GRvAagzE+/83IN72Y1ad90IL29I9mB8BkG7p+Tj+tiDbl
lxKlgv4639W5hDfIbI5PUPy8SAo0rsEidZl/gn+HJrWG8W3pDumBVBeSyL9/gRDU
pcGaF6J4P9nDLGgio8A29SXXHI1fsDdYyu6ufBrOPgVxImptcy8JCxkPfOdp7+xc
QDNb614fmf2drKNL2NDkDknJrmru0WWQa/u5eq2m+bLllN2x5lNEUqFjE6fDyWcx
imrtnEIbwhDtfPz1teFbm3sOY38/PsH70FvUD50k2PPR6RWzM1RjIsdHKZICKv46
BrnT95L39hQpuwYFc23o8auRpLWaz67k1AbzhicNmAqbeaGHfrGRfKk0L4Jm0coF
GF9Cy8rLq40EiXkHiprAlk6rYFT6mssBwl8i2GdZIHrifkZJCTO2O2M1dNdRg/FE
kGKYGICMYKgQprUhI5M4spULueM9DjnbRKbMhf5CpqhnNIfvSgVpCWfIhkiZJ0/z
BWddHQhOYiKJHy/HxjfpXy9hOcmLGTJ81P7XOIdDSz+FOpBN2zvcWovQIOPG7X4u
nkdQeZqNG7Ge0a7NBPkNYd0geiRgi2b0C0vS9Z8gkY+xVqoBKiPrwTgiIA+06amq
rTASuXWWDwrRNmh0vd/qhRjWJuURa4ywrgaXNX7A1IrEQ5g5ypZfWpn4+PWV+FcM
fox61Q3Z6vMlbcsoO7KC546LpSzkGDR/9Y6dBATi5xwNpRczYhyJ1J5bpBLnvai7
EWvuYg+3UZwIOgF8yArNR1axj+yLWvKEMt52vJhquORQ6CCMZPZnOMjS0snMnwSc
p9edXx2nw+jtPcmzOUnVoFXkpQrlKL/svF9SrKFjmEYCTQLrumOBpeYXE44Ykozr
2ejrDOr7OYuS0N86FuWmAcd2vTYz7aIHvbJUxs7g8PxEgKRUrT15K520H+TjZ7K1
T6UxPi+u1V+fWEV0xIvLEEOCMCexlhbONeZ2Lwj2IkIzqBZLdrr73ey0Ep2gg5q4
3giZcBlHot+SQzuJHnnKKAGyF3HX5FvoPvRyFYDbHKYJ9qh1i17V3mIp77kYHoJ4
fyafEhCqr10d/X/aDmM3lBQmN4mlrhaJrgwAluRGa5hOWhGI9l7f8XEVVDl3E+uW
irCIC0EUFLXhBsmLb75LjyN6JuEehSfnXw3+4guMKkXqBhmz686KRHFKicl0Xoni
HXfBvvxtos57abO2iG++65jJihbTbc6DPri9H8K5UcGD9b5u9cbLexar6g4avweh
lXbRvAZey0H0dHz8KAhMSzX6bqV3tYkPMSC7R9rjdIq9wNuzl4OPsxxs39hOVbiK
VbIPYZyurMmD8P7wPRnpTyYZIcfi31QZG/dDZ4jilmvYh1+QSxRDcgtutIkpyE7O
bjQ/UNpCTmK8hnG2O5LSJ4c65ChChdQsrGbmSQcnbbmGiq93jKpeGM3+7M5OUMVh
yXz5LHzPNHFhdOGd0/eg03XFbaW2rWXJshieeanzjWBCBXul/uekmYTNuAVGm1/h
2JkxS5YzxkBYmd7fczZpkrXeCkehantnFu4JJOXX1Hy7lWUlAhfirb2rhqGqgIIm
06giFEvrEC+ILyWs0MaXw3/jzy4Kggo4kDKqDkDoMKtcQ90Xiev6TVNTGJqLdW91
XfZh2TjyDeBDr38x6KzXANCexSUtT1j/0rNhpHYa1XLh3suJ1DUwft2DBMxJenLA
a6UsT4vTUq36xLF1prWSNGwt68Yq1m78DgEuEUulxafehvDmyFC13yzZIB2nTXOh
OLvR17+99dhvqjuauUYu3IDJqXMIpMw5eNbQHET6/eLdR3RCVP099JC+RpCJUF8Y
FkWUDIPq0BlBkbOfXThU5R5gPgiMBONZth5SnXwGtBdhVcQkFQ6+iob4y0pQzlPj
TdED7afQR9nc/EonOWwML6XZXIsaIDbG8Ih8kQLCsF29gazHGn5beyQxR1KIXvfR
KLv4QNc7lVqdS5SP+wTrA+W8WTVshq3fLEZEnd7LmjpeeKfWAsi0UlVZKbTGnzMe
Ef1tU/UtkFVURk9FZbjd1gueSCJzQzWtnoYs9SZWRo5pxxQPWxpCfi4Tb2WdQ9N2
nNt7t5GDBospX+KpXRulaOjQ6Prxraesgq1WHkGhWpr0tKG5C33lPTasKa5u3h1S
pUgfepDJeZETAeeqkVuHR09v2heQXmoPjxFtexFD8d/nL2ouQgsjNODvlCp7C3f4
MkmFIEI7zVu2gaMxhIcLNKRnKqKzrKirI+/TCKoOFf6B8M6/f7VoDYJlRrpNbetB
1twNMfhvGxRTQ/Tp8NjaFQAfxXUoo3ZiR2zZ39kcuWhYi9dIxIkn6ZmakWthAiY8
DCMSa+Ork+vPDTGFNVELgIIjNeKP9XK6NvyMDgxL4qwAFQ4JE/xAoiOUwR+98THc
D+iKvqP+gbFlET9aKde1rKmFo4ohgGpUflOKXXlynQPmFQ6OjSWCYWVxKoujaRBw
a2J5sx/FnWxcBHCBFAU14V1vvB+WUm5+7fDFTij9W+N+oBloz13L3NUkYebJSJEr
iGHgxmXO0BuPMmFlQYzITkftT/1BLSAqY5Zfy0z8DTM8Dya4yHRvZZgptFk18oAG
IKyq46Ie/FWESkyVd2klqhpmwwcDVsEuuHXDpcZvdyVmiDinVbGsNRqY1uOZ+Xvw
WUezlRW9UJa2mAqkja6Ahbc9dCnjyzWWSc01AiHr9lbR5TaiBme55AH6wB6PyBpZ
yXdqa2F4jJ2dTbMS8IwPd0iZIZwQWMXWNim+lzB5f1EEueY+qjzOqDnVLaBBTXhc
7Fl2MiEAB6wz/n9/DhDsdKJPYyR56O23ienl/SX9g6Hc/9uTE2iBtsqRBd0+0P6L
j0ockgs2CSafknzg7sciyZUuyNt+ClA6gy8RbtIJIzsx3g9lmK3Nn4plA6u+JBin
GhP92ZNtv+wagPu+UvKGuzJktXgyErq1h0k+E9NCSPf0GCIoSr3D1JCsFgbyhuNO
du6n76htwizqUOyTqmIvB8xEjySxr0gfXvZDFrHSstsSzhVzVJT31stk/Gj38Cx2
JTx/prtxrcWZW/jcZ2wwOtNu2eS6qfAubAsgnPtCyfkQNAbZ9fiCCVy1aHkXWs0Z
m52vbG6mO+hZql9YuPvkLn/xlBcYSNPRgcuDwk2XAOnkE0H5/mtZlLqFg9SmWQ8g
9VWD+NqdC+pq2dvsoAl8yYbP81gfitpEq6ALqTz64jDXsSlLIt6Zmy9WJuCa0d8C
DeRBm49tgsm6xZEU3yZvWTldneLjQJHQVSEuXziU7fdUQP0H9oGj93CE4r3RqNGc
T9s0z+f0Rkih25KSEg18dxF6omRUu7UEjoccRg04nEmZ0VcoQ0L6ZBCGU3M2bBp5
8xEyaHzeUqsMUGCi9eeTPD4UIDWjwZA4AM/SdtIANTWePFtEtfBzZxtePAq+AhZP
fb2B603Tst+HBsNHCvWL3GQ+z+NhxI+DSudy4p3YjP40FFIrfD0yInPmeUD3bsmU
FcDh98maBcxUU1leWOT6BGXCIsBMh6vokVuK/hs+a1OYTLvZh7xJGJdwo+3OZl4f
gKzvHe4KsnapWNAW7lYuN2stcbozC86xdT/QhmsIbKCslWY+L+51W7H5rGrujgbJ
PCOhRnU9eYvBmpAJnOaNq2LwTtydVaeQKp5XfWqxaijtVKP3L6ltfC5AxhtLZK6n
0KnrQwTZbrRsGZcrItL1DAle4gJc9K7QhvneIfp1Np6y26myMHT3r5m7jfDm0s91
3cAc/sJeJUDHhmR23NOEkNVkykQqLtbjU6yc6desJIi89Qe+VcypET1/zhaVT2dy
0Df38Vjl59kntXWhsMWmYYQTdcQhGe+4ZXTKrNvOMa1q4vuc+JHcPCKNO29MokIa
RakZMcXpc53RLE+ZUqukaB6NUg0ru21Bf/eKOfvrvdnbTRrvN/kSKO6J8/w+DrSq
2rKqGMAiE/bCdb7gLxT85uYTQtlfc90jJckuyYnTBTVVHdfMRJmvujqlk9uJUnok
oh80AmQOTchVW2oQS2es6qv2RCvvjRoRa4YtAF/aJ7F2ntrHiyqbG54bDBhLHfRJ
buMfDLNGgaIlH5/BIbNHi5leu69oMKbwdXxkRGHLZmNs9frM/5mGg9U/6exQrnac
RCcRXO3aC0qWKDbrykr4/eIugZnE4s3+ITz+FYT3Zs9G/UP9MexxnaHwrEJnzo8E
9dA2HOJG5D7F8PuvamYqQ8iz5U5AC2gZfIP6tUmF4s04bxSXHRkbmMtI/bicOxU8
I7BlaeSfqu+7bfT8uNUebS1FPku6orX3IFMGGXChkA5kPE5E9gZ3QFEZNOGa1Ok9
BR5FbNTlv7KgQZYmg5w3BOC2XYsLUkeOUWuPpIrhwAhN2c/gTVMD3SFK/2O9IlSC
pg2COoZ4Uysqx+2W0NOOyZ010Q1aQlXy44mcUJbLEiCtEruAudZxYwO4uSC0IG++
r7IoPfPc5LuIefZJ7VsXYxTyFwmDq4X+DVKs7JQIIZgYiW6LB8XZYBeCF2cQd86k
qa5a52kyY4sM4W+V8d94agbQMFmgqBGkZ673wWvvBGI8AYAcwORRgz1+1reBYPNa
xa18nfJZYBthkqudaAktCWEF8602b+SjpTDqZqd2KdEEFq+Hz+BTk4eLBKDcrckA
oHZwpBZjJk7BWxP+uYYGtq/NN+ZanboicmYE/tpEgSg9Qwq/30dr7cUdolzodLXI
tWyknpHk6bccNOadHFaI/U5Db7GrYWUavViM3WUqC1TnEb+nTIHLXfoh9cJykSld
jyu6MYDfEpLSl8qOgQjHprHslcc17rgrWvtiA9GDnEdb9VM7hc1Hz7PggX8zZMsO
VUwPpdXWiTC/yLvI/ftn6nVswKiMIv9DRY0mJ5kQHaXkgau7rk7RCeiOAwny+VQ1
illhJSR0I5d0iLQO+bOHHUJGtPIIQI8eRpkCl+x08lnb5U+tcgYWuLWQiWHG5EB3
3WHeM7IbrIdT50QW+5PUuFtDlEVCadzSnwCj05HiYN50eOv9BqEhPY0gWr6Zvmcz
+LgAOYj+27O1t/8trDUSDat6MTAOfbZDdj3CpHU4OLyDc8p4sFmF2HvOAvlNck8/
I8UpGwZ0Z+kJUPqOx3qS/20S/vTZCuKXdNiBcX6AGybmvhoGrYbPYnE/JY1P+9eW
x9iRZ+QRXBir3E67XSm2eVrzQpRuO3Q4IcR0KqDLInE3NP2SUYIdrj+YB2Xx5mBV
tPKq0McIAlAmqC6ZSmWiVdslzJM+RXWEba+ohn5VUwBJRTVzLn7DZDaVJbYURsAP
Ke9+lajMuSsD5n31dCCR7tC/6W7qTmwk+n+gymxqRsp3fIPe5OZa4PVv8qtogt3w
Ry0/zKH3EfCMAVE+uiTKp70vWbXqZJLZfwAbdbyHotTrGMkvEmS9HCwjP3AzoeP6
VU/1BxsqmF3qsPPYQEZl1hPJxLp4EpqEeGCJhbU9zBm0aQZX+0hEaklRuW/uIzSt
HLRWZZKB+SVL5FFnM5FWBggn6s54t34holidmbw3+62QzqtwhzYu/K2roiSU5jG9
0jszVPHFmgbfQCFHGyp7+bLaNJhPdSA+LYBIWJFItpzvEIppZH73E5S4PYtHrj+L
fTcRUjtphcUY970MBf/Q7/g5W3rJcKjmdAop+/bRmIm1HmTtgMJPgSSXymuTc48m
/EG5j1HJ1Y+641zY31rBn1Ke2mMoFtoayaLRsIK/wlvH8X7rkM5E8pQfnaHHT2EX
ZDctU/RgIA+XiA+VWwsg3x+tOZEl/g56hIXKOQJLNChXnyOBytKlp7tZf2l4uc1L
g37xXt1M6BNzt6KwbhxrGvz0Tshdni3GHLd2BRRrHXBjGpLJFoiFHWOPRG8i72sL
sLRORwtomHptwwJPqNIZTlnumosAgMQkq7Vd0I7b3DLgCO8ohN9gmVBVPu/r+PB4
zCTnj84+cAsanaRy0nSFdKPzwZaU1UZSs1O5Lk6ZZPLUuxGaugOdU803CglplZKN
FIC62DT9c88k1XdH1WwSPuguqcqe3HAHz7eCmUpXWJdgLliBt8j9O6TqtgmbCTvH
WNUjaW4fT12pCtrC4wIAT6hlS5PU9OY7RBoBvZsip6GN9+mbaw8rf72Sd2f11Fmz
Quex55JwbKPQjv3JybWx1LnQLIxhh5u76sNCR8+2A11rps006+faV/yTH+N5wAGO
DPVVuGYShR0/dGkU5dcPzK82cT++dL0e0blAm/UoqSk6yw/Tc4wj6WtltIMny/pz
LfMTDQYq2MqdfNFk/BxyFFDP2VMDFLaBi1SaLfK698KiG3WN0tl6Zzbb62yy5n7e
T7JZiK1oZXQuLCA1RTPA8mYUoxqP3LVICZlm899mm43+4qdM8ymni1DGkVzelJCg
YucxejcwXt8WmbmQZr5nD6GHIyi5K1Lftt2SFIdoKx/ATsToM2dLcL9XFJ5xtB1s
j/KhQrHvWbT7D7sEyGAxw8Od/vgNNAz0IC4ARombSs87wgF6ODCkCTp71LMm3CA4
pJ3DhwmurmnVce4t9U+rV0CQPl29L3J3GmTzgIFJABd+1wX2w7H/bzD7jAJJX9nk
C7/Lv4vM3okHsFDDk/ZuXd7gzh/uvbGLQW8RwwoQlnFtIbakFsXflN6O2HxaN/Ip
NEG8rO+plmO0wyTo5XBe4OwTeOIG1DW5eQMChA2ZB83tVqpVYGDDd8zh/ufYmX9M
a5uJfDhoZPjly2drbwFVBGsAU1wgMBab4odZTEvsYt2gr7Vk+b0TtWQb4SwSRG3p
x2285g4D2RKWXKbHLjL0AdN4c6kxLFq5JayXVY5Hn3YUIJ+LAGc1uA0jDOxvvL3G
8Z8nh/VPwws+0gxI3Uj/SF7+ZApSGQfJWYxd7wwdtJg2b00m7XetSDOAoJlloP6d
9fHQoPyPkYdCHQt53rpacp/HOlLrcdda6EzGLOCnA3SM9pp5TQmbYU5rxLd/1h/R
PkbAN05GRFWy9xznXWFCbSSYWt9uJZu9IlBr1eB5QNv54xZPc/gkSKHp7sZkNlxB
TpDhrnj8QgvidcEmKfFNE82VpTlaDCulkbZvIYFgJngfWpRWr0kmy6NOpYdS3sPV
K7GwQdwwAK2WKBRFnHhryImDNXf3usUtn5969Mo85pXJ65iBxlPCZTsrqmbUB5L2
QOdfvnpZUsmHpxp9fp5f98H1vLH6ZupV5qz/fjSFxWK4ddGbOW3UmPaNmVKq1BQ3
psIC1XhgFSpKSnZSXLSscuXSqL8cdUO3rck9tWzCmMZyS6y28xCf3DmAYfHC7Vln
kjK5NS84hC68/O7wl1bF1Mltl1QcgyMI32rKO0oZ+4ghjAvsHyzjuHsDOrFcMxRG
fjtd/8qe+4UuNkjp1oGH7VpoB/XP0N4W8+YrUBSSPg4OK95M8DuTARa1oMVcjV/t
UccGRsHDpu5Hf38oPlyWS1Lbl3UpIiPKFYa9llDT3NvzBdVIr30ZXoNc/vevi2N+
u+MDl7rKZa27i3kpDB9vhK0OyU0bNlYCuevxSimXKpqcvX/F1Yg0rev37f/y5nN0
EwOLMm6hCtsx3JLbDgOcvXNJxxFuI5krE1WWt4zin6ZhhNCEjX322MMfOMD6sGEV
2BuX/CGwTPk42z7cuhX2FBaXSyNU2cE3VKjPAM3sqGPQeNmhu367N66CDF8MRQuV
xEMAFQFKFakt66RsvcqSr4MLgWk7F6Ba4diLjkXNnpQGG8TP/sbxc4982lisZpUO
V3c2AcLYqmcXmg43FaaTIkqQ6OKzpHJWqCtBY3OAMhYMQbx/YzYQPTU7a/8yzpWx
vXTVDl1ZieiY0k3OZCCfy+37rs6rXpqdRZpjfI+JC9lBkXaK4waTSOuCUvbK0ll7
AQS6nef+dqz47bV4DsFmy6J3lIovtn0nhtBNtoH/VZDm4oWsgkrPht+mKY6N9Zk5
wZ4JyR7AWesklRk9jHa+3/CnHkIs6AE+1vkrY+5OIFoi9ENfNgyOSxXodIQmMnjc
7F/ti/Qkqo2iGAa9d+OXvZ74axpQgDZSOgUjo6EJpLpUEizNd/IK1gH5Q1liPkQj
YJ1B6CUZXFkDbkX1MqNoujjssXmuet3iANUHSmCd0VM9BNaTRFouyR0nRfxSGwda
m8B8MoQ1B2i/KFaTubS+G/e/T9umVCNmfaxnv/+mW47layIjMzLYO1dGadgIlmds
NaIVp4aZuJuAz31OOUmvkWI7Hp9yDNH/n6XmlpXdnUxotWZOH3xMqGVBT18DrP3Z
h+xlRPb+Emzc/rqDzRsZG12uFZbHRw4jQr50Jq+jcSPOdYj+i80x6RaCx+VWXO+r
yc9t/C37V4aGhGwDkQMglmIKwCfmSGpTqnyH6Yzr/tPVGEImWRR14QzTpUExWo7P
BVua9MwTKGB2RLHE31Vk6zw99j7WR9Jq2+IQ9+aA0izUxs3+bIDxyi7y6phBTIcR
Ahgoh5zLfMyiSLJ5Q6xD37f4kuIzI2nPjrczrCBa5jpV9Tbrk43zhNV+Pa5yEnLq
MkQYt+NvhXVUJAiWmwQ+2lx82HrGGuVXN+Xtj0mUrPmOxPYTqHsgPlLbF/Kix7Hc
L/u1bzbmttZ8CUnBq8ejrgXyQtFj/M9nUPzwfjiOjEoNJa/MrF1P1dmb0usLpTyq
d5ox27W+b+viTGldtjK64Fbo/DSddad0JCRJw530i9Ga90BOIzdjLcSy8Mt6MMRc
py4yBhT1KeN4A2rZ+usrLijjtwCOg5I5D9CHHoN6diWqwxVAi/yhP1bavl82QqF1
7fkhXbldLNi2KN3R62lLtOurUTCPJpZXe6mduxBHxoGpCeV1Pw/V4QnHUlf3VZ/o
MddaMU79l1neKt6EcTGCtCUgwqMIXPy9YqiIYc8oPz3K5TgdASXOWHNQ3tjz4GC6
Yi2mLI+iYwsgirGkCOFMRtEn+uRPDOcYO19osY6gsu1pkt0g6azE16CH13xtgqTT
d9zi4HTZixFxOLnG0Jy4rxu3Z8qsoT3Rt5y6PdF0QLkFUuLctcfAjR9ElVvxIWyN
5xStdTTv3L2xNY1IVnjwQZhE7DiWpOHnkCvLc8EZB530mRWySyrGys4UZD4IZuUc
rveqFJa+aoZKphsYvzCqdM7vpXmRUdkvT7hsHBtxLEx+hfOY8abV2+kAaWqCD/oE
sxKsqDkT/SJwUNMjtSBOnBxEhSCPSdEC/1kUYRNhJ0I6TnjoEdg4TkgVpmAqYzWT
g+uYGlr1Kpc1FPO0iLrX1nNOy/iB5np2Ew5HURQMb436dkoC4pfC9E65ZlqO/aNN
6ptMl53vEQg8yjrY3fWThBX+rQtM57RyKOhREChHr8AkqPbKoqdFFlRIwytam3UR
vtRBMuO79Dz9WwPuKjqQKKmE4o5r4jAkLqI2H96SKg1BccotSoKsEsSOaIP0/RJA
vmQlSS/lAtCT4qlhlOfR/wKDlhfgTIo4772VDMgpnv7TWOzpuXUVbZkumspAfigk
gtxZre/QMcby752X4OzX+5HuF1kX/gFKjDgfQ2JNY+5c5GScxPcpeTmJuRSELx8k
TzbSSgy5JXMcRvIGNGjtT5lbdvqP7EvOqL/5AWcSFgy/GZlThZ17rTVBdchppIOr
Lm9NS+Vb95tjMohfJIMVZNdgyVfV+SbOmpNdPpTl2RgKhGXZRDU3GmwoZ1koeNPN
Ut3T0K2/Aix7UcE+OJfqYzPlgt5IPdybMmwB11PauJ9EJr94NNq57AMWd5mqoZqW
BMMNbIVeflG/VJ+YToXj7nYGB1MZdR665xVaSrVwkuqmbWFMuzW/NhJ0L4BFeHc/
rLRl/Ldn9iXwSVnZgbquUL2GaghFMgkIVfgyffJ5uKHClfeNz/drzy6GZv3RnG2z
/XpXNVh3qyfmw9xuP3aUFJdtSoNtlbRmALJhWWms2w2HkJiaqxGjP8f/RjTNmGRk
Tn2IHeA+M/0ZGkT5m9X6PmZJQ1VmndP52QXIvmr8hNeMFFozlOXgv6geYz4kfNON
sCEBU5rLJWFLx9g1fgU8KKbFF79G2YqF6B2F9guNLF1m2c8Uk5L9p+DkzeFP0I94
HdQA44AWvA9sGS7oLjmzfw+gr5CbpWId5ulIcqtBN56YIfRZfghz4sJWmS2Y9fjG
rVrWDQ6fJ/eY+xT5xcMqzzElK/x5tZoQaUoGbs1ya9AV6U2JcODFdYmweFhi88C1
T20SCm/kQU031RtmMTbecS4vR6gUyg/Y5l7oadOg/yRLhNcMVE/LG0puyTpVN0wX
78mYV2C+t7+deBgbDCOqzgVehLt1HKBavak0NvwLlOg355PUygStWGhTUhXZkE4i
0fbCzSTLsMqrUPQfNoyepZu8Wrg/P0BJEElLq+J1ius1JkxnEHe0dLTvvpalCN14
oOAC7pHiKh9ajXTymiyBNqNHedBJOLIvhUV9a0az8bNBwlThog3AFbHIivZPv5V5
S5e0B6G7r5wNNOyeNAqFtIc0MjUf3e44wuKH0vxNLBv8unn6vG11jpGYIOXl0Tlx
rskwtzwF8A7/mBNxxrdOvshCS2Tl/W1/BKxaJyGPjdnVqWn2QlqOmO9OPaZyS1vn
upd/l0Q6KH5opd37J2IXK0fu6UMSxGV3OSuLmrFPJjR/+3MbfS3zBA9Q2yqDHKUq
opWNps4RbZEjBoo+mFx11KfJkwbl1BACygB0ACgJ5T7R+M+zihpp6FSqrh8Z6JeC
6aQ6zF2l613OHsYIjYGrywImztkvi+ybeI2Rixx9OGnhcTW4USkYLik0QSLJ+XOv
PND8HkxHeudIWC/V0RQHzPHvbQUPk0GvRZd0dPGKEQOJ9qikr58Bp23+gpaEcaiW
OcmwXNTS+Y2GTqnOciEocbroI9dfzKgvU2Xres4cxW1/GGh3tocEeeQJM4m01ZnN
wFbTgXzQhkTooVM/2wMQ5zAcjJKHHzrUceYGNOgiME4QAcnSTrK33aq1RIV0ZOWe
wpntnxfRgm3M/Lxb4crorN+cwFXnn7y08GBUyCTR+4sbEct1SHjFpeii70dCASoe
mw3ag/5p42GZ/95iSa+mQ0S43UsQxcZzi1289lZp5CIE4L48heph/U2EiqPEAi0E
QZtzIG1vZ6gkxcHz2GKDZ6+gc0Rlfu/jgszNyRnClR9/lLcB4gh9CexKqWNv6htP
3Ut1YgaeOKN5gv1/U6u01do6K3VZetxdexS7ljNYM9wvRbxm+1stumcmm68ayph1
asHCLTtxQT74XfqQQFg0T4NlZaNGehzo+FueoEx2+syyTT9J4NNzYTmNFL2u9nR3
svR9QROPsxszdB1tbjRCZTzlPN38kDXkeeGDpTxPV3RbQCAbIlSUCb9b0xfGKPWL
M4qhnv4LfCsIquAmHwN/mWnpKzKk+/cRFeQnUi5D8hexJNCvTpgRAKvbqZSDjSUG
Ze1UM+LCoGjAgGQS536KcIEnvdqBF/kRD7qh5nFsjit9d/jQ4Ja5OJO21df17h7k
4fo3D0MNE//8Nbpo4G3zrkVjrsljY7jCgvSck5OStquWIoaYGq+DMFICgehOAo9a
rgoy9teErXiUVlbBLIHK6mGQARdd3eY/S0PkiqYycnUXZoD/vsjU50JmVM35nkIy
REN2faHNvyGQZhZH0skcBSblaR6HfuoDyfJEILbNuTP2k5cL4LqmPstzfOYnUv0y
A3JuF8PGq64YmPiVTx79ggFlUvPJYq+01aJCDO8bF7LLCndC5OyjZgqUkUUqjZZr
nySSsGNoL5H99OttjaJnfSZOEfmxFVD2m+hue9Q1WXWwGCOlUT+213IYocFkGymr
srDHRtwDjZzkhE1Brgu0OG7LXzvOvABetfOODEj9T1UJsuTrpGfwUU0BZzW+VcLS
BzEkbRQ6P+1gKegMMJjYdgNhKf45Y+K4lZrzOftwCoNILEmz+5CE9osndrQOQ5jQ
s3pXdQGFr3d4hpYo3okaCMXjnl5/Yb7vI/+3fKBhnRpAAGk4ca2fmcje2Fv5F+0z
MMc3Gg0ZaA86WkibRktU/0w1mPM+AtAWisKKEm2ixZbGzUn5msSZwDKwbTBjTKUG
ATpvM2GlrS0Plp6CmQnvuB42aBJxvmI2fwjxk64MFe0L/kdX2bHnlxkU9d5Oc8Kw
K9u1e86l9PmQgOmER/cOurz8xaU5VSD6QHaN6cCJMZQWufA4c1UVZPha4n/dCV10
NVA74VdXLduR5BuA5kS77PugpCBcNQx53wIe8qdBrJpdQlgqFGUELmNvScxmk6Tj
gG3LfRsMhmcKWFYUvbmIQKuVaJ+FkJKLDLa6/W+BnkQHSxy/wA3tHVvl/q7yCbqw
98BhpjGgp8z0Lm9jKEIxK6om4LijgleHgopj2Dz9dz/fjlbhTZP3Jv6m3jIpZNie
OH3lBH6EfdtlMkgyBgvm2y/VsN88Atz6ZVLPXyBBaT/b0jJTqRk9LQKXLha5g6kc
yXQhZT8mzcN8wpaXKh+gqaqaTb7fRppOxzXLXbwVIr8rHlz/zCgkbmU8GvmI+yl9
KQA/mb7YjrIvyd1CQDNsHHvTXjBkZdphl36QjJKnBpPPu7joHOdQhOejCuVSQC2Q
4h7PJ523R+RPCC4T3mBU0OP6QOv2sDvN+P09jW70aMINUiLb0ok+ZJ3lS7SiJMe7
eVOHklGUyKr13VFb8msq39742KWUubILK2Cd0MDx22xE5j5oHR5HEYkCGmBych66
/UVfriHhuaXTgFu7VA1banp8NYD3lz0b+4/i2ZoQnEKicc8fOxh2Ew3LK5X52Swc
w8nJ4xhZNEj6hG7Wi3GxzxAxYE+lCAe+Q4saYJszJNMc1OfTNrGYosSqSw7TWrQt
e5a5d+cppE2EATRnmuxIZL4GsOiKv3Hw2KHndDpdMqpSTsDUZkwGG99yiXKKdorA
PjL8YTBJ9TolxGNf6R1Y4ArSG2q0bVb1ftjbXK/rDiRqOyHYRNJ1vv6n82dBPO5B
Jzr5ObbPuf7PPYksikTdEFbFiHlEiben9BId/qh8b+hdP87PchkeFvxC1Wsy21pz
YQpIbG5E3MVZ1HV9wqR3Qp6oTLJe77Z9R+02cSS60lhKzo2A8sfFiguUbkiZH7x3
3iP8nhWigLwFf3swwgwVF1PiJ84rDphMKvHnfsaXtQlixRE5pzX3Rax93BYu6Cv3
eMOWzQp+DePmRVwblLLPmJ8iyWOXo07dfhaPNszCbr/6/SLw0WP6aYT535j0e0ct
DddwZgEDacRS5VnsJGQ/zHXLgSRM7QkaKZMLmqAQ+ixGGF8DSinPK3UPoqErcyqa
3MutbdcWHs3zyPr9bEVko6LiXq2MtbeGic/shZHZIR4Ughqu8ol6cfSqpR8u8Q9V
FG2O/MXxd20fYIdHsKta5Vdn7lVgHQb/ToXI73QwSFxMRrbIH57fFYiXK5DG0uvB
2W7XTSe5oRBa9gh2b90lJDmlayX+wIEyG+kiGrXz5JcmZaFFWt5PiW1fHHZjJQDd
t1QkU+rcT0S1uM2d4FEMGEq70edxrQuJ/Npw33jD0crU3CIIPbu25JzQ3JIFlaI+
bA999ep0e+uptYbSIsboy0RZWm6jAuvMyKUSZs/FER1Qfrm9QJFKty0tfNlIl5h+
DHqsBp6420AMYvPTzUqIdi9l9VutEtYkNcpJimy96F764b8f2CiFb287ZJwVP9uO
B1VoAU6Ug3VNU+F3KBzwCnxcPfs4k8lg0PoONwVvJkag2EM0MOwgWFkAVDX7uhdf
sr64w0AWsdz22A7bjb5mH3yT9YYti54ZO/0er21vanhx07PObZUrHpU+iGFYXryg
X9vVFoo9KvhiWK9/MgOqQm2Um5cQA7AmEQDwghOf+CrwFN2MC3dB9leSrs1Z42ZE
3SJUiJaRUGXKQUZOVHw8BRfaKmwk5x6oLcavblWsi2VxSDNwupY4qLLUBs0hMkbx
Qz3+rTegX4oKQa5HAscxLlKavaPWDagehqIE2ukh1wlV42lg8+EufgBFhQl+nbLQ
aH0xI1JO4w6+dMN8p1kf15YPCYcvwTESTDIXqLIrBPBm0hQgWmbdnJreJO8b+yuc
Op/bX/yOujhUjcUZmPQB/RYgxZAM7OjAchnSZg0t0aNq0sAN1gaiwcuWVa73jO6+
Vl5GkI/QlpD69RUD47cFGSTUBfg7qKj0qsQ7ZVImZINCBze0fW3t0A/HvuOmxzeA
gZtioCI/h52rZe+N65W/SIdqBYrIF24zZebDVk/Ryvt0/jMvg8Z9UugS5v1nSGMA
Oeo8TuNLn6x9TvWF0yGZzCWwmhKGCfi4PvyiPQkxIN01hT6oOg9XNvqbXL/MbVeJ
m3a2tLMtDhmQuWeUDqo8X/rB2eiEod0ZLgHAbX+QuLdr0GERMIZLdGueoTGZUWAU
5ltyc05xFAtFMwbOgypP8UGzgOlmT+KcATF2ipqGr8nmi8Vmt29rEeRpzQeXhm5o
rtSbA/kAFKFQMDTjI0giIbN7HfiAlowPQg00wLl+3hbodlBvpwaAkK2fbhzG/+J9
TVjGDGbArIuMWtfDRBCiZc/jG2PegrvYWc6kzDmXNDuUwMeEz6EPtQAXD4ZbLWD7
DkW1JhBRK36yoYCwfCkafCJzUQgajF3KqRwpd65NhHTambIkt/sudVtVZVL4rbIw
AEehK43DbV9Zj5ZdQY+RlyiOyNaFnJheu1fjTXDl/E7d6yg9qgF2NLnTTvqNuMev
0fOK6sVX4Mv5PhwXpQMnM1NTQGxADZn0Tmbakv9PcO8iKqPAmdfdd2NlM3SW69u1
Ql3r83SU0PotG7m9pEPSuLutwwYl2qNCHWfd0j/nX0U7JUepSZpwHVhHnW11Yqgk
BLm86Pz2NfXdz9zRG47arRI34MFp1uy/STUDJVjyqhguDnLMqPCZNuuZfrEHrW7p
G0KHRF+PIR6UxNaZBCcxFIDTatNJa9HWW2dPj4SkQCyry112vPs66T8zCiOvEGTw
VIyOUpEilVnf6wdJxeXL/DQC/d/oPUh8QcIVhBEvQ6ipkG8OVBR68RSN2RGc6XoU
EsCmOlseYwYuAVW23D9kxeYLkFrONThckckmXgR6a15b5lk99aDOZ6fwBCFCAwzZ
1DLmi99IgYa6BfQZ/jqIS6yHpcov5d/064VoTzNhiupJr+/BlOLShz91aMOlLN3O
cAc92iG02TzgJhsvy0v5h3hHROB/DdgFykOW+faBQW1pLL8X4BM/rVNuJAyJ1bIm
KN/Uh+HjHp2cqM+uAqO67y0S0kOkLy3ZpOz9zlXDv2LmyLR+C0PKNyOFRrfw3yzq
yRrrV0qF6KYCfEI/LlQUQvV/Fz5VVgCsQu0xUYXIk71wSBeYdVmbbMI9vWqR3LO2
cElVwmfpjnN2JRFM4lTOsR7HgQpC8NUy9T4830CR0XQ0rnAh3RST2iC6/hbFuowP
7p3m7O/OeUvXkQbM0Y5oE5cYTEoe1i+ZMgOU2cHaVRe0l/pxGuo/UIrZKfHYutbz
QUIAfu+xVyogebW2jmGZz5obobA7bk+G24M97wVfasNFVs+E7KAVgJ0akWDahY7z
jy2/QkUp07NAHOXgqakPHD5Uf83C6Sf465flcELZC2+jUasHl9Wd7/GttkHrna2z
066KkLH6VuqMeT4EtTBDcCyU/N0ue2TAI5uLid8maX7jHJrxQdjIlvp5Ev5/x5s3
XrJPaamrcPT5a0M50yGwEkyLwMJe5TN+Xwi6RkAQljQaX3lvTobnsqqE5zgcQsH3
yXoQwBrwD3rnFDQ5swrUNWnXXAMW3VNnMPkqMkL0p6JS3f08vJ2eCb/DBSHk643s
ajE2rzp+WrwMwLI4g9koWWqNFEir0crRPhBjPs52ZKgPqPGMDFNKht6d5+ieIwue
R0u37Nl5k7vVp5WGX9qMDH+6RBkzuZen0rRkNsr6hVHBcZrDFIz8clnwkHL193wO
R9UW7T82W+yGMrWBpjdSZi/vhmuu4qkOiA4egQ2uJzbuOaa2egwYd1KGL/g3CPRt
l7zLiiN/l0yVHh9++MBkmBG22UQxXUzh0I9kfZYe3VVf/+ebcbpAYPSGkPcBwu7e
840sScsAVkhhua2SLMctMoLKbdYXNQx7UqRjFKyK8+pV170H0UUzuKL5b/NSCXYb
XrwGxBnmy7fcF2/CZm7e25QODgNWcT+k7SohwAc5h9IDyYs2ur7fjtDCeZ2IR83d
M2fj2LtxzZ2IkkQUiu7r4GcOwSKkTROiqV2U6IxavtZNFCjkcTUTtWFmm3zrXLLw
VGIPM41Si8lt64aPp0K5Cdea1WAuidEB5EkX8orZdIrE5DEOVcNq4eQY4gzbW1WF
kK70gZeh8ire/a6WbB2CVe1BbFGLbNTzyjA9xIcLr9HS0sZrp9g9myWuVN/ZDA9Z
QcuBhGU84WlPA7fIZiJQYiRy55xSHADYyKQzUMBueNP9uqiKop9mQ5nmnvN5DCHs
d3BbwqxWW1pNDpy1ghTHEFhpb2GoZj1J9cO2yg//hYQmOYeP8UnXENMZxkdLP1hl
QzrZ7x3Y5PJa6zN9OL60ewcm/Mk1ms19zx1TwnHrq7z8USd9MgAZmyrpM76WRJ24
30qLKSyvGN5RDY+LKaNPCWTerBMXBa2RVyPH0jrnt8SfoSIqfM2BX5U9iCVC3ck8
2+7PM736NgWq6pJ3BB/TbWLcZjhSzzOJeEeKjb+M7k/kjv1smqNtfnFQmmeEMGWu
jJlDkKbXTMrGrPsfSZ4BxUGrF9XuTWcCJN1kQzs91mGzvTNv/oW/993uSERmYjMT
e5oIZRRBp69KiMdVlX73+TDsVGh0rkO3Vg0aztkwrZvN+cxbg3/7D+ezeB3ydDhu
VE5hJTs+8pKSe3lC7EFm7OUZ8SRkb4e7ReEQEKZPh3JZh8o093qNhqoNHyfxVlMN
GdavVyt7eq8/IHo2f7fHzFcWtiay268IKoHpK7owwUyBQ0VCtqNNWGAh9QC2Pfj5
6pwVMlUt8Hh/N7pVn2qkMQ3n9bYgOGFsZ0RAJB26jJb5kHU9Djergge5dcx6ZBur
+WbGR4zWzkNlM4FFFHB1gWnUATCoeQ3BFBWRknotsLjlN/LJx/1mIFPgySWavfFN
Wz27MNpp6bbOJ1zWEkhlM7LzZsgcQw50uV4IC0MYNNdBak1djSgwYxt/8reiI6mz
3GuuodUbiqiaYt4cqP12bBsao9WxFi7+8H5pxhuQ7OSXZToRSxkVZtD61X41aThP
O3MtJvLkD/B+Z8MVA+1eNDZqDaKY3tckAE8/xhpUZ+2ZIp6cN5H/qXpgZzq2MtS7
opHc+85Rvn2ONvF9CPB1cLvtkxYJKDDPqYAnxkt0vDy1PHse+nt2A+DIBNzXh0X3
gZJFxF3GpOQv9yQAeGG6bF0cPHSAFIAlOE4VKNiFuKPlzSYD0I11gU/TBlKlXr7B
W+cndIFVeumLBiqYgxWBp1LLxSZWth+qSANIdmFOayAhn6JbcgBh2TGmay86DNgf
Q+Sa3gu9+lr6UbGgoDhaOaTE5oeEuo0mM10tUhuJ219O8uuptxShg3YFncf9w6tm
U2ab5B27fnkPGl8x+lUiRpMWy81VNlDChDbLJ0ghZ46T8wIg50w/uYrVNpQYJ3V5
SkRaq7N08lvROlaf5Xnms/oRYMdZPi5Qp7facR0HU31jxplAWVN+ijP+Kj86hE9n
Op6TBFasrWRQYmrI2vwkd/K/hLpRUvAu6q3t4csbmVU20QVjmT7f0857HFwqycNd
EYN1h6FFWO0kGU2h2TlskX5avXX92P0z1qzp+Xmhh5G6N9Vk2yL9/pjLQXMEZL2z
/QNQs1z0+PJdv12IpyQX37t7vKvOMvtDaVQO9/0fT6nBx5uxgg1+dE5oqN/bR/To
WGA6B4ILOlyRTMvDMjkjX+jgpsxKJDNAJZOAns8+BRk5yilz5mFRvZBrCsTxYJ91
pASnml7i89HDh+eALfBSXCSwToWm4pF+zrIerTbyVBiiWgCulr90KpM97s3/a0my
1DryyDD69DdooXOdMMJoAc3sgxaGYSeEyo+6i2UD4qebAvd68xLfk9ZRnixmgkKL
2ekacMkfwtSrD85OQC1bFn3ZC0kiZCi3uOXMxxQuoUSqouoGpotXg/YkSfekCQQ1
aDjoCivGarbyVO7AAP0fPs2M49cae99wmrrc70zT0W8I3C46O+g8Jqk765YvVDOw
tsB34EK2l47fA5RVgbCDDqpCK84sFDnyYWEHQbCM9Ko3M15Jik/qFloDeIivk/WF
2H8rD6RD9ECqaHEz/MsXpkcNwKWyy1YzTA60P2ZMASr+VueN3lPL5ysFysJnzMTS
gnDio6IXyTI0fzhE+dIWOOAXox9KucVnIHlbgNf+HJbZ6hF7gABbsyJlMn1DaA1r
zOdp88Ji33P9+VrfZVinynMjWOcEyNy82D/0vX3YjTLqMTgMr1vnLnV9RykyhUhA
p+h9x/R+xx4omlLGZVx5Ho2xrHGJXJZqObi3Td9I8CHaeJZon8r3rSWE/iD8j4Y2
CYWWwoznK52YKqoRjX5ObwqQYoRmywfAP5L4UIUG8IBploqcQqQ/8nNHj1Li32I/
XfHO6aJel7NDqOaQia87rIHlctJj1OX3wsJHpg1RCOo/A5QzoZ9Q6UnjqjvDGfOh
3WslNCHPNOMwlRBggCFkwM6VGYfjZjgP00p8fMYaBmQK8iQUi8qIVb29QSjIhcMY
YaYHHu5gElVcIoW4r1TWlUkaCE+FAcTOzMVTxwPj7fpL4zaCIGKKB7sOBNu/f33R
Zjenlzq9XVW6OwQ996793uQ97zhgGUUjmkRVMlbELkjYJPZTWA6+BlyW1cS7w5R/
B38kYGKvrBHeUrdkr8XRWN3PlcO7g5PBfv+6Friyffv2/plUig3JIayPxsOjs7tc
sVFnuDnyczEQlGKV0ZB2j2oG/BA6upBcYkTHoR9qN+WnlNnTzcVi/d3uQkbo5hT+
RoPruFfCCL49LQ7kwGmLzTB9lIUxAI1B47J70eD5K5ZHZGoljyJ1I4tRE/rcaFxI
gOxLk/FqKvOntOFizJRcQq+Zd1Nqz4JHdpc6oV1Zfa8K+EV+brg919JQ7sl1aTb6
jOrEiiyFXFYOI9LqpGjrg0DZjqnb6wPhWLaBk+8oUTRwqqmI+08iuu9XhcSma3xy
75FcMYbZnks7FSKYQCf6x6XzAeWE9vAcozhVG/AlEA/9jczIiIPpJ4H2Ojm9YmIN
K7j1JMKO8uo+B1cI0f+nXKPYt4teAC0D9x53zcdeAyIGU+zKo7/MbRMf4n2QIncn
wFUe8ZECO7+065KlsOUS8YfYvCowc3zS9uJXgcWX0Xq5yXUn+f3SIAeQQ2da4mSb
81bkchg6dvWUcLFkMqvMWu3OHtvqoShdNeUf30rSWRYvxpc4u8HYCFICxcYXNckB
grBZdjZ8+E7MUNv9IVtBL7tZ/4UONnAYKq0mH2lxt9n6rxremIoRKFFgoFyzuJam
inJ3/NLxsgWQzboFOURUB+XfYcjdz/rB2n+pxwJYp4td1ouDN+gF09ZsFSm89TMB
S7lioRh85b4Jlu8IzlsgDMLXtb+8Y0omDbMR3vIejWlCnmfBZjKm5lfGQw6Sqh2m
2YuaG630r2gKFvX9UHIKOLM2o9wQhGR220R3IgS2/GttcdJKsOXasccG+qiCjKkY
8gyUBiikvPKITYsd6lJikxIiSNrLmdAiHYyAoe/4I/7SAUzKXXJ9fcVZzY05q0EP
uA5aQOBSif9VDAaV5A8mhi+24uqvGHaR7fH0cW3r/VVS251InlAR34+jpxNNgvKC
N7VO1TaGPcrsblFvcKu7evieQO+MGR84yhUNTa7daJyRn4cAIv0Sn7ftBAw11g0b
jinldZlpknQA0WMs3lXfYoRTSJ1TrHn6S1ziUcs28pXSUofXQCeYgQxFkADdZ9Bd
SyhxWmj6/h9o2X2H6haups33aHvL6dd6TF1LIn7Qen5svIQOrBxmn5cwH1OkyBmS
VKics1qntOx7MmeMx3LQB7XCZokvvHlbUKeXWSI6AMED1f21cAnBPBa/75wJd5+2
+kDl1C54hP+NBEM0cZJdQvD6WfHDAERZUPmxfDonuTRcbKLWNIYw6KSbRnHdJ33Q
DlSsX5xIba0W6nVAo7+zum9lyHBxqP74OK9F05ljCApY/E4STyiIslOJI54GqakK
2cdUUSwWTD5B9c5ZqTDrZxQt6NrR+KqWMIpQC42QA2K1QpclUdUY1McPolFMq+2u
dbTT8GDrhmLulDlVPSKQfkxGcZBw4e0Jvl+AVoNhrePploIVPiNv8OeWOFrPI/fm
l5Ck5T1/z5AiH/Fm3xw+VGT8y/veKS+a+5SRiMtxJonHAvzlOtM8+UEvSTi0Yjd3
3KDZmS01sbwIRkX6R1CebI3y5MNybODk/fCR/ZVLEazyWKMgK07MqqE4dW9Udc8P
FE8mjQ2ddjgOzyXA55faAJ1nyIafTRb1NQzf/tr8QtRtYEtzpxN2rhVHNAnhCDFd
Vgat/5SUKCOcEjxtSifJA2wmY0TU3A1CpmBag8OSOXBVSj/Y7/jCUWN1yO6RnweH
nUa3epPjwSghJFUML+ceDGdvj6/wn1oBeugKZEK6vheVlvzcQmWW8PcBOlyGc3fc
UXiFi2c47yxMQprwh0pyV7fibKPiFOqg8UzeNve344cA3qhr8ZAmgytbrBykJXRH
tKYS0/qRjtGsc4doJHSk3y4KWyL39eZHkZYT0Tjrfy67EbknTNtEBWK6FpCqhB5Z
AC/s3Y+G8r18ZQq8RCdwEYbwjKpkRlXlLWqXER3bSJJ57g5iSDwE62nZPaPkk47R
2mMWat/QmW+BUCfWXlCf45VBexsdjv/uB9NvisJEeu28bstB0XrXTbiyj/WiOVhO
8R7U3cotcf/4oCNumEu1bEH0rcOWNWb1J5SZ53OjU2JXip/EIxsTKi8tmRyUUR0G
nHFBs0HdONepkoPrI00EfH4CS23P4rosawVC3DqBcYYFrEV7Q0Q9Nme14re6//zY
TAKvtbtYhsezisy7jb/Q4cKRxKzgzaOa+yS0fcw6qSczFUmG3JY/coVYE2PQrxG3
TcObFYCVoB+mftIaV6wsPiBjcu4ty44rC3zr+NxVoq28IjNR75uULKvDPcKmZMmn
YdhpJOR5y+aF7pdobf/4KKM35xtrusWLhJQJzZ8yKYsz8HVd5TazTq97adB2Gq7o
WFURdw/yQsMy/gk6lN+nt+hf5Ay5EuhBYe4b3YAe/XfFROFAXMQEjcCgKif/IUxb
GVOHOzCF/NDMX6G7clA1v0R7KhsAEb+RDjqaDJZ4yGw2ALmDiudKVoIlqsnyokm3
UcZe1JdKkvhw8OYKzb1JIf1AafWuM1jFt/mwrkrWBneIEU/RvTlfMAfyBHz0HvTK
4FvWAL1s/82w1V4zowQBm78jvdi9M6+UOa7YkMcijBa9/OaQvt3/FVIHUwdA/o0B
mHukLk71+6s9YXnqRSPw5uWKiZSa+1sHCXWt0EgHlGTL7ybWr6TIxqxeekAzJ2rR
cxoeUg9EJRw2IphUAu0i/DiVjnbyWpmXOMpf89okxBcImjRf7T1lfv6w1iniJjfa
b+WdrWeZXukMQcmK/EwLD1ItGx/jbC2uI9ExqjIfuGeMOzMQuYVRcMKlqdEG/3WV
fG5YfccjgDpnLwUrGKrKUgM4Zj+qkJdxx6OwTfK1w+wq1iZs3h2LqVFZsNZxr8GH
02pAyDBOHSoVhuXxzUbqSTeBlEE9WGe22uvayDnFyVjtja+Etf3O0ttmC0jG3Xxs
y+2B/0m2VoOTMwe6yrdr53sfEhxNsSTKhxSMFELIsWW9bryPA94GZzrbfHjxLAUR
qAd2EuFEs4OnW1Mee9vuBjLINTBc4sD6GoSEtzciSBsd/N7Z6wz76f2DAgXKGuz4
AB7tioKEbkJI7dXoUhFERkvz1gslOG/3k/bLB7PbZy+RGHHYJCpiVOkJBtkX7423
z2RzMMaxj4Qq7eU4dXOw34WzaMZ2rp6x8XhUDzbUr5sopN+43LdtpaA1WPeyeqWd
3xt0mtah04C1oMbULdBoab9gBvKE9h+s6bqtGTciZdMI2HPPCXTka06lcnTZYAp1
ZwydekVtVlgL+uZNLNqDwcZJffd4RNyd28yO1H8hbXvw0Ahbeo+2cgsyUn6jbrK/
df1qBxEz7er13TiKdjADx1HdDaXrU9huIDR82LJdjNAY2VmOvO7htmzH0xFEF8jo
JFh6rhnNjwTfYXYt3/rvrdeePtpchdKpW1myAowpNLeaPjFyxaXhs0KDo9Tr2/cb
ON+et5CnYz0K9ESj3IxJ4utVUlNrVSorn17xKaiuibW4notJBxAk3CZX+iaB4BJH
wBvJXLml5bw6IAkiDYhzYtbntm3usTw64ZVOf2dKsCqQth3cU09DLSou2mJs42MD
SCYfnrQT0vtJmTIr/mUXWY+m72Fex5+nGxtmwn7RjCMPnv8LNh0uLEGEt5/jNrsw
RL5WYLJaBPowHyZJvtg0+UA7BnAQyKtSE2z8dgkHwJhNVVJNKYNaKxfcKp2J1dgi
hlU5Iz3LKjVM3VVk3oWEr9fuM0T37F3KcLwem5uRm87HggDDLS023y+xGLk4pY2h
iZAzGLKVBJcRN2gz/4SY4YBU7aA4kTflAdMFoOv0kbPicmHx5eGmqMIm8u6i00JD
BDqfqzuhpikQJOlaim5Rh922CdPTVgjqfYb/z5IXdDQgnl+SPJEgXFUIZXpRME6L
Ha5rvMUy+RtunIFm5+6WJrhUSLp+jLLKWz0HKMwM+QIdCc9l9NWdE0qlj/viWqg4
uoGoEI/R5nSbujRwxF137tnLnh7R4Kj0tm3vQzcWrVNgFa5InqFSHb0gJLL/fEZa
lyd6Pdpa0sECR2IB+s0ZIMw+GGvsJS6Yg/bUIwegOb72G2isO1+Xv7mj/xT1Zkc/
mFlh7xi3BiSv0OSOBTk4gUOSDGgwhAbjmZ+zQpZ6nBtqerga3iFLj0lwuZJ11oqw
FjDNg+g+EOMfS4tpmNv5ILEZCFHUySPCOjx1eSRnxFGLWQAfN8XBk9c82k2dqWIH
9fhBxWNQ89F/ng/YdN4MDYzXOt36uohiuAtYbxPa5NOOPA8UaUmzIFYXqLmubJyr
c1cCey5Croz1MXRF93LGMwHzq3qS/KZvwLQs2yodrSb6qv+m9P/8ZGNmrcbVpKTS
BhFIK8TBf9oF79FsFuwDMjb3FBnGHU0uO+ZwBjbIU9pKU7ZXkrcIjWfVZjpVnJwN
38zcft12qrXhSEx+aVUk+ANSI9xQl89JYbBgPERFySdoZ1A6SiYqdbUSbacW/A0A
0CmmKfYA4+Zoq0DvpIiz7QGqWQ6w+QVY8t+xug8+cnO9KOzAXQgYvFZR+IJ7cSh8
Qj1b4Y24Oe3c/O5r1CJXfok0tNqd3y9gFYVeh+IlgrUoxTABUnbALL5mAJ0Imqwh
L+vlEdh1/baL/7BOX8Ai8xvJsnkSEVc6xqVS1K4D9/e3Va2ZuBhjF9gEB5TuZhaK
ld6veNMZa7Gb5zxeaNG4kT+9rRHpjTUT77VkGXdEgZ8I2qzerL5KBFT0cVdzDlgV
BIyMbHfiV3EJG5jw+Bu2/nLcgnpjV4WubzGkyBInwC1BlO/mhURfwXYZyTkBJP+e
gRq0eNK7FxZXsHsw0qjMX53NwXFi/wIFa/G+Xy2bEymaxUk6RrD9WN149wUdarsB
/Rb2x7FtBgRwNl4hNuiWkDdVlArMNeRc0/G/xobYX+6d3wojWvNWELpycXrxCFAU
+OQs29oW6KzYwKs6qEuHIUEENDne8iJvVSghlsh3nDXo7MSB1vhnQMWZwPPY9aqx
EanFT1CFEo9c83W0awa9/MsBDI2jMSPOlvkT0KMjoAsM7mFkP3yPpZFPXf0vIdx/
m5vFIgyiZReREatHX2Zu1a379wiC39p1uW4ufLjI7exS1ebwf9meyujRVearG5Eu
vUNYVH44Y4Pgw/SN2c19QW/jQ1e+NXhA3TNba34ypOuuk5hKvbbTWHK66XXJk/4n
4XGCheAiCNx43q8o67w+ncaOOFu5IhgTkh4RiDGwe4Hkx3UFuts0KC1PWF5YsEF7
oQhed6JmqbQQF9jVC+0G674tXLeDaE+h85+FCGcf4D3L9MKceMzfznu/wI3fK2ZP
wfnwZ7LW2fQ3xnB3xPEXZRKsVAiLuSDJjJ2ZZKxAsI8ESnVJyc970UkHVVi+j8Gm
Yalib0HHPIykIkScKKEMEStp0Ql3hLQ9mWuP8REVC4ivxf5Fy6q+ZiiFN/KvVCOp
G2jp59Xxqg/UlSiV8EDXqitPPhhEvuTWCuOFDa8Hk0Af0ZXBp5UdXY4QHvaBVEZa
Q+e3mW3ouHqq5r1c009jlztm0OU9nzxwDpq9AaxNr47YPIbgkZzFKrE/lfHm62GC
zA1eNDg0BNhCqpmZaevzZhLPmGEom1uAbNAvSpakjsBkbdwbppny+NJqSQvoOI15
0Ho7DFdNRK0XpWLY6tqSr07PQi9NmH4VQ/ttkzz+/vZnRWSZ5ud7xhh8tRVXSMfB
CExVzQh/ZWicQDxWgWYVbqd3Y/2IOaUvtDPnZmMT/zUQz8rO4SQNWdo5Eirstzgb
AQ9N3+2ujH8kMJ7spaFo3ZroIUTHGoUWv3t0jYYzZBnL5AEJizaNufk5s4iKApli
Cv/UxCLbixQoUUI1xM3eb35Xb3OHmWltevfRviOz/5lFpRhqR550cnP/d6aPtLs1
6oGP0JvTqV34mWOilszQpDUyGPjMzuGzCsG3OScVo1xfGOvHlcnd7g5CXIVaSIak
y2H6KmMr2MHSJ0ws64zPSzjmxMDC9NvOLOL3phMfL+44xnbJfEopF4kylIzccnaA
FLaGmr6HDlMD6kJKqiEon740srRFbwf0gBYZ+vABdrDkKVBC4wlpElFTFPsZE/PM
OCler6Y/8V5cqJi6DQVtalphftASp7eK/dd74LQjc0NWpsnrioEvjxFZ6ZEoMPE7
jVjRnFfVBp3VGzv/SX3LF72ErVQdtavxZMGK2c21Uim8zpcQgqi1W56D0rIA10qS
2b1fiQTq+7OiyZuB6ojm6xKKnQS4Ubc9lrPKPC6SfGCwWhsdBrkMa9FO3Zg4rGhh
MBQaYnjkAdPpL5NgJzf05SsrqCo8qqvyDx+q3sodV6mfF3qNo9Wrtu5X0mXVt1E2
E59UXtmniCMMZlxUKEWrYottQN0NAAbet+sr8NE2KhrhOfrLT8nkbGzUPpjCrJ6T
cVM0Co6wwa1B5xq0aacf553MgYLRRAOTYpIE9zX5Sdmd+U0i/0Ss7MLm4jfUHStB
hZoRGKEkfekBzniEYn15oPIh/+iuQPvvxuFDfnDAk73oZCL7V1okwrVKB688TbGH
QcZwdKQVRZI03gkKWdODz4qsq0Mr29PCRNorfjvGW0JMSul56H9lkKz/i03ZADNY
/gfV437DH8DkT5ECOkDS8qT3A2vM8f50fRY2Qr3Le0xFGatVctTCdL0x7uN6CMaM
A5e+p1vmF0gK50o+7aVAeSEI6XeZ1xA5CTGN2whHs4gpgIg1MMg0VCP4VMGq1ct8
iOpSF0SkO3H7mKynnavOjh6hYffeoAX+wCc3M/Nec0rnngOSlJ8ElXmKYnGtQFgN
gelzvVty09dSVsLpYA2lVYvse3rxVZKebn3XWtNI80BGKLn4ulN9JkMXHzfw4u0R
s1/VwKwI+4DE9VNlgsl6VznXJMUQuTgeWwHb9A82Zwng5Wjx1dgvLuqKmxw0RC21
EiIP3PpwRKNy6+W6ydaU/tVVZNmU1MlxC2uJSLFMdsQsV5/IJnzQJrjQ5XjgB28v
GMc0W9Xz2Ip7KT35J12yFJeIlq+aW02/FY5taDMyF6U+cchFOFKxTHwYzpExNsD8
Tth/bESEngWWxlstmzQAr92C+AZRigayk4rHFnrXDPDYZEl11uIJUpyW7RfQhQKz
sOM7Fz20zsNSjTHPMwLXtwZZtTkH+HMb+Vlqw/m9YdTm8vafArSXjybJ9XA0VrJi
3bdp2YQDJhRhPl/n3jOIdBD0wCfPSkGKm2oytLKMToDuDxZ64pJ2WoLfagQ3ULtr
m6J9WOQa8esDRG3Hd9/tlP310uLac6HruN35B5T8PcC1+QTcCiovKl+jhrbJySvL
vRqC06E9SzKvZOnFeSPA9lyHTFAjc3JydMvgMiQtMRocNUyOP9x4PR5zP8GxiD4v
4SzNV/RkU1N9GpxX/TEpM1A52v4ynwkiN5GBSR5MBBO9GjZ8rWU7fYddaj6rOmCO
6pN99HQ7uhSd/pyRexXqc00fx552WYpFIWjagoTC3FZCp3HPBxZx2xvY10DzbHu5
VjcALCb/NzyN68K/nZi28NTV5VZQm1Q5xDsHTZA5kgoKkNbPTvFw9DUC0qG9+tJt
XtLgYY+Frr3uvmoHZqknNCRCjADVqvTA9MwlX/Qvt79rLv2uhpb2k8zKnBjM5czC
Y2yW29NBosRyZnFvD9RfWOACcZpI2NIxD9JJ5vrAkxLY2BCVN40UouCo3KKr4yYS
yFLOOQnrJxwX3hYIDdvGPFyaIB6hNygp3ABygrqF3+LLhLULlmipwByAo2qM/QFb
QRZ26an7BBAdJYCelf/oQWa05Itgzw52+zajcsCFtA5v+DnRntxoqxO42yreKRdv
O8s/yJvZweJ5Kdp0ZD/7KHF/HDIDYJIp/071f9eXHQSOPw+DD1iwwI9wDZag1VNu
pZpSHDINsat/YT6cc0tCqC01e61T6zZnDmsY1rLKN1R4hMze8TwkOSEh1l7frryj
yuP1zxa0E5NZdLbPmaciWSa9pv9I1Q4w0u5M3ioNAsRxoCi/45HPw8oks7NPPhi1
/OUjsCF+dIBU6N2L5tByLc3KX0QoRI32zE5QH9VTjeY7mTnRBpEHo1Q9kQUdiWbm
Cer4EpirzlHA9zZ0TJwF3Ib/pdNgm666STpjcjyfUIJDy9SMgQiBtyrho5uSLRtR
V8kBV+F4nJB666Zero3rQiMnVK1cjqgfhCZ74Uu3vKKYh6wsR0+SrirWEcjk6xr1
eKAkZ2O72nA1PvlxDKl8Lf5GneQlDv6tPFBami8zjrQR7+fkN7ml/ulsn3/UXFkg
LxHSEQzV+er2vS78bnFsgnOK5FzSa5vf+RCQshC2+zs800774uNU4AG1k2fkLQxE
VY1VIlLOmPlmgaTP279ZxWfkrSlPTjEAXTRULkuyojtiGURXmmq6B9hR8W0Jwjh9
uXe7eZih294wVnJ4IRLauI4FJiRbQe/2ZuFkW3D8Rxmh8yToaZhs1hBEBBfX2dhi
Ry41AAaw+l7Sm78KKjelHogbWCZgg/rK+nriWj3YYE8uJjAbsxHuVVV/1TkBtED6
tZ3beeiLKk4rHR3+furh1PrtcwKNtolVt5tFCbwMiEySvqTeC9KH6g343B3MndE6
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aXRbrCcpiJYnaFnZ0YzCYQAch8Xi5WwqJmkOdMlLUjox
eBLHGobJ13agaBHRKWJreRBO7PhuFfaWh0V8kLT/pbhsUngMZne3ol6j+0cUfS7c
2WqTCHHu+d0/iBGQhKR2V4oVFuJ2g1euTZQISzC5V2vn3/DUrpoQ5++w2Ty4aG/7
87PrT8mtoEAclpvfAmGhpVe5kPeBVq/P9QNiUup8brypmhBCNhwcTaoB58wKfxu5
Fa9IfEGhm4biIM/SOVK1walDe2+p3WUObbt1D9dN/mlbWjp4CgiG6nS/4TPUNYND
3JWKx7YLcR+1ak/fMRirWtT90CKMwDv3kjNAWfDwNEzfQN0nVkSj2if1UliPqYK1
DfjjESTBosAqav4WHIofOvjOsOjxFdTJVHbb0a5KbAUtkxkuGbWpSuN/jzNqWQNe
Zel1UcfZmtp5bnxuucHZ7Q+NKccVYh3MQDCfou3Hn7y3UJnWtwnpuRAx4Qcjpb2R
IaI4CwrsMkLBjWloLbK5UtxKJCJBVol66Vy53/a2OqVWCLEWOD8TQKnH9zRm9qfP
JwBASbVrV3m68v8fJQNTr+RTkaEApDamX7YNdaE9H/LwgDs3efsZyK+LoCkSmAfj
ubOvd+oJvl/NCrE4wbwV3YFTv1lZq3Iz0VDiu/+KzH1/AT5CHv6R/GnW1rS7J1kI
DkI+raxDyIJh/6GpItOa4aunLt73cf1786I/d5qVjjNZT6PRXQTB88DfpZWio+OA
KkDuY0LE4A4AyxiRzna8iUnlsTzgFJSUc2AyWwhPdANzb9r1d/VnvWRmFypQPFrV
wQjvMR8ZQFOIHNBofPS7Vx1M7U8ueu4dIgq5ibFwTAZWLHlgK6kC8r8rCP/HsISX
hSy28OUIrfI6F9NHW0GRuCYFoNSyuGzfewidmTOMw7UUMqE/C3Ci/sUIHgbdtcdi
MpneN7bvGI5kdc73eoETWmFhHWSBwPbotuPmtKQaO4gvZfYjL5b/uKNCvnrg2mH6
CMbkIht0k7AaRGvdn3V+OBeOQSL+syQ2TGU87wmRlsDgJbMLTXyd09m+gNr3luAg
df8YfRZirVmpsdoqkloo0j0fF87Qe57zZq78gJS2gp8X2u/YkkMrtk1f1dWnz2SR
/jmynWiGQF6EpgaHRv5v60cS+s/DkCOG50GSkLGeypdKXKA1izRCBIp9j8L6/b98
VMvEK9Eqrh+eg4kGftqX3QEl26RXiujXR7QErthlQUJd5rKklKy0F1AkTpKC2z41
JrpeqDhrtbF8wwAuSFqhnNlumXCVHOVDSvaIIjC6Q5+yN9RwpfsGxE/pt14II8yf
GW8sABZCdLOf7Q93Q4fUC8tCdGgxR+4c1BGKrUPsjdr6sC0s7OWnECYotQl1J68e
MA7jXb68e83yLFzXALmuc99RQh3BcpO2HHSKIuy35kZsyWkEmx5u+S50i0rc5Xao
cNh/IjQEDcYUVL+BMLlCrqnUrICA01MrG0GBBX3GlqnPv8zwsx3jTP0IjbHv63VP
0kwhS9wTYWNZN04//od86IwgUbtgXdvJDql84s8b6HZzE7v/K4OozwR635hrExs5
6nWeZTr5iRLJknbC1IMgjGMSz7uXzrulZnPCQUO47x4vSpAdUUmiowP8KNYx4Zip
3TUjgr4G/PIEygBeWDPCGQcL4hgUzyhaBQmcABhYMH7e3iVGDrpRCMsPSwkdXvH+
0fsKY/hMG9U6ADb2OcdziSDTiyYswfrihNvquKt2kcYE3Wx/NmGCXYloLNtIYUBl
PA2BmhEq2TaioaJS4Bzzb4CLjoURVDqR8JmwZlkxf8QwwLas+vl1wO7C0RicB+tL
mNDBWB9pCwdewy3l8gBrgACJsmVkEjRsE7P71ZO5tJkrtTDO9dnIqdY/DThNISCs
c6liHq1lTGNTM5xnKBDw32C219tpBi1MrlMzo3DQ9+wM9NtF81DVn6UyW9vWI/WO
G1bUDZXnIm/2buolanuqgKWHEJnn6C8TpQYmz94PP5mfl3SDd6xo/Mjv3RQQn8EX
CtmcZHXvovxYNggeCvKo/UHbVOnVESM9NZtU9KnDHkoKB7HbdSsHcwbj1TnKYmFO
AwHMo4H/3thIDeaacSd3P9WenmTN2PsN+sVblp3N22/71c/luGt33ElnVJCrODg8
6t0jk4MRrs5mUso4L4vyDE7lLPotkj1YIfCs34S+SK3vhvt9EJ2nUPD+/WYkgRkU
Ilw/C8Q2Xgytg13wEmFlJEcoxhinelpJtY2yPwQlz1iIeQkOS/3TYeEDbrm/Rbtd
z6qBeJ+Ej+H6hgUt1TcMm66UzittJl3YB9gCoGTNn2cIOMDz5J+RUZAcIcIyXzAA
hk98xQWXLsPFR/NK9SYUIKIglqUEeNzYIJJw4BP7SY0O25KmeChA4n6of0eVKk0c
Kg8B58SCjkC26hdU7/jNbVHblNFaep8sa0JOIp9MJxxp8L8IDYNfanm+aozKVKh8
qVB/riln+XHzk334MSGapkTrxPTPyrnNftTQJAQPwE9kYCUHsE7atiYhmDSOHHJy
5U42tnSF46gd+QGL4Q4bTOXlrKX8itbdFbuQjGjg/oVv1nZCNdcNccinecLQJM0E
DYC8tW7tkKbCjNov5NVFZRDUGNQiu64yEt0SuyU5hJVm/6cPpQXIKuVDpiOmbnr+
vY/Zk9M/+FeGGqeLBira44HIuOSDXZpmejsbfgyXmB3DbP5HBnXR4pAXL60qbk3b
6aoJP0CsJVjhBEPOCjH+b6B9tH+A4L775Yl0+FWYIJhNBdoDCj9tilMejPu+6O+M
S6GdPd3UfUkXHDFRPUJaVkA9WIcUG3t4fOrsvKld5CujR61gPIEeZD/lnt9hNDWI
wDcXbKDMQfwuBr1bpISI9InP0eJ7qfW/164ulG1I8zNW+OK2AvZHpWRRc+YF/XgS
/F/muhMTS75hFk83l6kL9qm8HHmYN7tYrgh1tKhqJn4wrTHtwqGO/AG9Kz5B3Srr
9GAw3l+xKtO/pCpRut/mHiCRwZKCM1+Nq7x/Xxki6Fsk/fugNKGnBXLvtwM9LHnt
7K0nhIJZe/eQ3y7oLsFgJozl4MwA+ijQ+/RexHuOCdxoP4Bu1qKLs2gPpdRvZj1x
95sHr1xEidmFwj+iNHIcz/bwfFaznaj1Vo9xLNz8u+I/naTQ1xUupxFgQAV+pfWd
VArqMtsBnDAZafdcftN1OvakuPsFZzMTP2e+ybx7b1cc1rO4yAgmJxscJ+ERxNxW
HOlVrd2qA5tjzDjVkEEpUxy6gk2BacU0YTqR42sBI7dsJWBGAR6Jdhv/4leKWCA1
v7KpqRDKRQwtAexXSk2v5ykml5I1ecZPz/eWFJU29t5LvdH5JTNCGqxFtkMd5C7a
Je9ZaC7x8kxhQDzl3HSR5Lycmsyd5X9yHvrWiQj6YCaMnfW3yHlQYVNVzL6dB4OL
pmJGzZiZgfoJ0INslob4Rku1ca8CocsnYwo334d7y3b+B2yRs0KG82MH2CmE9tfw
QT6GHToKRxzuPZKUtQdoyKW6kqKZhsWJsblG5RjaYQ4Ic1eZjkIiROUQ6lSbY74a
j16bhVaCHDv0G8EgaKIBoTQuneeM25+NI6LteXnJy1Igwf+CXGuMJuKP3qlScXPf
ySCRZ5Fs0v+K14N7+CWItKR4NTd0steAkyVPtHdermaq9NIqH/eAfrJQjuQl6Mg/
5zfo1zHSnaj//it9/nWbc6ghXnZZMDmldhuGHBetoqnB4ROu3LPMgcklHYQvlsIW
Y2LxRnqMy8X0YUmFqzk/Li8HZmd44+EviXRTyt9stIOeKVUy6iTCuoNApaOsMXE9
TTjyDWlIK2jht+bZrYQt6kCrB/q+/UlPgRc6V+J5i0a6j9iGPihmOAb2t18HgFIw
+1+NNM7bIx8O2f26ZRvKXZoYWk+fNSDtVo4nEvlv90JKlAWh5KkabkJrz1wwBj3J
82vXWgPsbFAYOeAV5R5JyxdITr0R6LDL7Ml+ILddIN6wvOViASEd80Xjkto1/QjK
kRC5F0kEEZ2685NOQfP2ou/wXvhy3gPbiPgAY1n4Eo42ombexNv9A+a+23R6PWyS
xRR6KykQUdSkpKzMg1wuyNVLzR/43pKN3yfBz1PYgPy5l4z28l3FW987WHumqjWs
IVltRb3LMwEIUUtUAAIcius6/oDEUjTLUAqfSfWVoNFCcSxFIkw862wRIgMfWw9b
spJ0M9KruDPqnz9d7ZC2Kg2nre5uC2R138VOaW0MCY0jXG8R2N/cak2EABq1gv7B
OAegPqXZ82+d457vKq/cXKuXmao8R1pphBOnBzjHrkb3oIRp3ch0YCJZ5L65ohiX
tb+unzYZ1y76KVBK5l8Q/Y3BdZBdqL8rMTrlDj5TXYqmu83ceqrcfVWLw7rsasvu
6vGIsze3H0lUhb6LgLihE3CfKzD54VlzOqEne/qdNWesMAAYHWNjitOz8OktV7H3
OP0TeXNqc4t5pRSLVlHxYWu9v4aZCgU2hhNiB+x8Ga00cvvWvm6XJ72+rmhkBKco
3g+Sfpva0+8HFU+Poz+PgdtN6MrD5yO0zQEzwP17lNUdkLe/9eiiRQla0juFq5ke
EoK2dGSNg64tTHlaT4IREISOFubQbOgKtsJfolMQ6csos7bP26i5W/J1CXoyrz72
19MyQjWJn/ufi1VQl29CTM2ig2jK1lhAr94G4WJ/OULH0hn7ooc91ftGeOYggOsA
Pb9eerMAGaZZf8wx7nFZ3FzgkN0D0qr5JD1YQPJ9d/kTw6Wyiw9pVaaAef/TpI5y
xDIiRa5rEhrVQIFRuG5zIXeSaZN4WXo+Ua8hzEgMNpj0F2SviqHAkvEqC790/zcF
D+Z0OE0o66dCfA7GY9ApWaIlp83UtY2DqnwPlVQsy4YG944DnXrj+FQZWq0e6uD2
roigGk8zNqQ0CrvNaubCaZUU93/VjAkW8K6krk7MAolNBPZGmtQxx8Ymz1un2uHY
7s2ii4XEIpcnH/lvMyWcZixrUAUh8F+5YqFdBTKzDUL6SugIDdklxpuKXB1Pn8ex
Y75H6Fq6PWacRapNO0V5mRVGExWUY+sz72qVWs98l9J/y4+nbakGeeclzLntUCba
Psodc/xzbkqOzvw19s3e/dODK6J9CZsOfi+eQzS4FgN0RA6QXX2UaEv+/p2pbZ5h
ianwd93KdiVorqbvlBN+Q6eszkkpNwvXwQSbuOCWi81zGs0GQaY/pKbyRbSj4YAg
h8F5tGC9gbhwqNcCBd4vvfOjQUx3Nv+NMEvPQLz6JzWKPnJ7z1FyuRxKpqK9srQw
eDFq/4p/yY3WZ6UtQANq2Xuve2CNu70keTZzf8h94k4dQOik0QWSWXaOQY5AQwdK
HmBG5gCcRpQcyN8+8FckVCS0ccZTzNFAudjnTCcEKm6KPywJh93lMLrC6uMFs0Fv
0oMH5b6OPh9L4Kr7x+LdKxbDKvY5oszuN5sW8p3UVWhmlaGcsAG97cDprNxXGt3K
ejIophGpMFkMg5EXzWFen+sG2b47ql2wS8XeZEPuypMK8rXlR4quotVVIEU5V3RP
x27HY+E1JYgqy6sZ4MoV9Py3zcb0Ax6csofgIMVCPxwQpXnGKWX2Xxh4mNbiC4ee
I9/X5GlwzwAr3ag9kaq2SzMYVcVyQWeksdV1ghAL/Bu6hdBN9JL1SDu7VmL9YPMm
dC2i/DeVEDNr4ysFJRp80MnU+AYPk2ImyOXKRKkEOHSe+lKSj+jiIdhIxAUlD59E
rr9eNKVXFUk69nDmBP4a5BmZmm3D5rJa5Ax2ABk5jXK50Iej+chr23SbNBTfRi6/
ZT52yqFZm4J8jE6qwbSOd/2gjMGwxO0phZgDWQvSNDFbaUPTr2CJ6hC77wKnQlrp
jT40Xslqz/tYc2IQb3iYW9ymSG5hIcD1Xu0yqz0TliOItfSq5hU1uWg6tKZ30yNZ
UIUiunyHQEi1tHRBDzyZwHpFM4G8FTTKFHoyqclTpqfQDFKM3qVjHNla6NxVZTh0
FDYnwkWpCitVYNjWP0b00JetXxBrq2TK2YLGA8gtdHmCNw1KqRwQtpf4B8hDz7ZS
9NR+Q9ArdhEpzS5KIMEd9VrScWwNR1TXDT3vzXtYJDhknVPs97jN+4PKA7qL9sBb
im2bbt70txEPUZfrzp1NSGOTTTVt59/pAVg48XXrm+Bzqgnm7f9xOFdto8DXnh2U
jvZ6vAVJfSyseH4SgGcfeOcSAHk2capNLcln2MjINmhWJg/YUUDVZsutO5f1DXic
dzksSArQIch/YcWbG2EYEIwFwsaTEd+KWRrAJ1nzHwUee3fZ+gTYrThde8stLsAy
DoIN+qDLb0bULGtN02+QOLPCsfXc/HXYXJ8HoPRFZ7/S+BuGTEEZn7eRdk+k6Hnl
DW4Lhyt4QtsFSPgST3mlMAE8OWl+XhkN/d916QsVWWds0WeXzRSq1tGsmnF5eQaZ
DI9chHTwdAuqjS0sc0+O0b0Oq3iGf2oWP3+stu0FrCANH0O5DjXTRTpkABFIZQpz
gdePy5/sQekshtSeoxoe+ag9/SQtyzeutlyWnDhfttR88+6i1dEZ2318BiZUzSyJ
Q3tFgS2AD9pFCYmmqEQi77DH1MAX+WX0zj7XelRqLU6kuDlTuUYB6hZ+gIsDUan2
0wlz/9auYJVwfbJDtIFt7B+3cl87cEBzEs7ZSqwYocPhQVIT+TEY/eFdUGMNpo9D
R1KhA2OVgXTAgDA2TRyp/AKOpU8HDTBpj5A7tyhzeoDduDJbbQz/IQPwW01/dpDw
20raVkFq2eRgXwPMCaPaVL4bFxptHucTUcG+TiDqQVtf1N6c4NPnOwOxJ2gLSYOF
zcvorcKRnQh47bjcVo09KPx+G0DlrXj0kW4P4HVmhgB80i+WFisZjGXT8TuVB8Zx
kh/4UgnHF0lgsdR6Qb7fejszFsw88cYkp622SgNO9uyl18dXlpUR/y6pvZMIcexl
FBjApOLOH36dMxsl2VDfd3ixH0oi2DsuXiZdO8DEaafGire7XVjrMz/TXnzQmUCI
VnhPlyZXmvC5DGb51pcwB2/nzserqURC0J/2zE6D2SssWhdlWo8DImzDv2l8ZkWX
mPKEjU27ZPTA+/xXABkJgVykgo4LqmmXchfq1WjmYIv9Wom1nmqPT8Qv0bqsyR0r
67KZvYTLvqTwoeHhPmGnOdlQiOWI5bTCU1C399D3dsgeJDyHRRXYGKfZR80Gy+qQ
uKw4QWu6esINlrBG9biCpD4qPi8R6dCrcqXK5stUkuC073GlkkMy/3sRVy9zSn/z
OrU63Lcri5kj2zEg93aDzCIAHQkDy4hV4CFY4pE1cwzaiXAcErUb2p3zETJYG05L
omxavPCqS2lDCoWfrG/Zu+FQ3SI2ggtGQwUHJya909RTgph03w1zTwg3ger+VYjI
52eJNa+AVYczDMMkG4pEMYWrP91Sr0ytwtLxt4Yz02S2bXvhzvQkXqZ1ws9Hi2pM
2915+BtbyCl6gJqd4di3LOX86QaKul1SOQRI+E8wHfLzLbyzceWc+bpZdB90lu16
YGse4xNdZ4XS1Env1ADbkBJEjY6j8cYf+GEi6D6jkDKdVims2T71d4YrNfaTJOa2
9xWoaPveZPn/7fZaXslpr28OHgFzLLww/j+/jYTaxoZ2SAyga/iH9EBlOZlnInYs
6zfXtTZGftHyvsaf2rQy0bi2Xd32TFKVXMIJW4g8eh7OyzDHbO8EjOTcu6d1+Zcr
at5+eEAk8uMxlgJGsKHhzQET0TmzzaClwTe9eMoxammJwaBwyQ1uWfD3TUSZ8kb0
1wBby5cGmAbfhzQo228o5LRxGmZncoQeuhK9HgOg5SCiJ7rmPQfWYP6dbgXm5PwE
7JAub9j5yXVclZdwGNBSNpfp1sHCN3r2wnEJTaKC9eMkqPI/nO+zahdFXBMEitJH
hcPzBx3fo8ebZpkGqku0wESANOIB7Br0sb0MT64LAQ568YRWSF4YH1n280tJWvY4
746+su4dPxGHDvDTMnErQogPu1vy1H7omh57Yg4ybgBtWW582JCRWbIVcItdsmU7
P8un7B4KlpuSULx3ksSERRBCmgY9IA+tmRxH0Od3aLO1pfjAN5HQDhtj1vamXixF
tU4+3/RYQZVsl4NpwHI5ZNaNLrh303knE5HTE0GLpz8Fuxjgch6PDzfIM1FkD/lj
zFfM/FpS/l1b7Ey1Eoc2JfhgAkSQ4z0/TSVm03aKwL/SjpTetk+vuz2gdkbUffqx
wDckJhDV5yzP340JN0VCf0+mozOqgiehGbDveo5kvn/YxMUL+46MN+K5L0Hg2ckj
AipDR++9dYJmg7P6DtAFJEvlr9XF0+DaKvfkvQs3gqmn4C9FB/Z/A1AO2vamEKT7
H/mk0PptYqojSFgoBi8FH/b9mteoD3+XOi3XxdKHIwr7KHuoNu1hNvqHRC9EbaFM
/6F3MLle/FAxVJ8IW7aJyY6tnJqX/jp56i+FXAeEbAUTp3QxGenwTnnbIRvuHRE4
eIuZq+hBkyZXuWyaY8R5PWvoUEixn7UqrYB2sfgchknhlbsDV832lqDuZ5ndUbVt
SadP+yTnht9Q5G2QoDzRKKi9IonwRsLfhZz2lP7jOPOhKQg5cWRAQQG692xSex2/
Xb2Dv44qwAHhrizuTwBH5FavFpCicB25hHtTQc03g43mbtfncQtEs+/3/gUPx32a
g1OAj0pVgAUP4+2HhhuNHtOge000KV9gWuHqOLisdAQAIkErx6EDe1lP1qPnuGlD
HO+uaM2eEK3li3C+psTyIRd/eb/YZkMgwhP+RT1LDtznd3QzAD3A8uniAgrGb6PF
qJORiwMucjHOrJO4BPFWmABX6YwxH3TfMnOZCnHII4NCZBK/4smcggn3EAiVJCSL
FZn8ZN3+BFVk98A0PuhTEySrEPX1QnzSvqZ7moezS6vOQgdtjcp/06z+flb9BKXB
NqYEuw6ySlPkSxrV+5R5yqE/ProJtlDZQWUCBVqQz7VIAIHFVy7GKrkklqdZj2hH
DdW/kPdggP73rq4AcPYl3M6MnrXy09RBTvp78vdEaDAG3q39wfhGYI6NEbiuBA9I
snNC95/G/KG5S4LO+SXPuMVFiRKJheeAFiR7EdtCk4aq0m7elY0eezUA2I8b+bFh
20DO9fgUjhE+iDEkN6YZA6+yT9WAYm8TlR8d+naOStmNb6PUohAEMg2dt1lGSrFA
hTfGRYl8WefM8T1ThR/BiAe/zDUEvVavarS7f+yq41qEUXxcJ/HTFZXbzT2/HqBz
N+STJJ/OeXv9z9OewJUzktoMAXESBF2Kx1oC45temXmtCtODsNSCzLc8WRZONJBx
9rWFDYEj9A/BSzIW9K57WX1SZk9+qk7WKZHglyX/Vw19cTvsuNnQd++jPp4SwoDR
ikZEBjAnzjMUdAzx4OdhkX06FoKo0zsGGlnIEGOnId1YLSGyR9Yz/FBgHiQokSv9
BUspKpS4of3/wVTLiV9KJYe9Rnv3wb9Pa4lyqeQiC5JWBygw12KFSAVBf2bUU9za
u5fXh5Qn504bu8imu1cY+bQuNbUs4Rpg5PED2OFTysa/TFu1232W30l2byHFSCG/
HdMl9ZJCXGwjqXJFIOIQNjqKCR/Hwfj3VFMzm90XpCuinoQ8+XIdluBtTzCKDMJZ
Mc0gFJyLE7tiPmQJ1aL5UFHigOIgWF6PzTvjusgRMhySlSrRL2Y4HzfAV+7bHzsW
WfEnW+GDNR2Eqe/OrGbMA19DYpDFww+2Vrdn/TGG4WGaMvoSFjGXkyj9yDohEJRn
ImzLX4ZbLUWjVzx2uqbgW4NotRq3UHpqxMeDOC3gaMI/8RPFUiRgz0T8XzSY2WVg
STAicACuFdVGUD15KxtmWWez7Afdpe+kQ1p+eoOutzJ5BijXus5XJZYPfOOHZQGC
H7UUU0tPbwwc8ZSTk1Zi98+P6tCqdQaKi8AJrwZx67P1xXaDvuJ81jfFAT30Gd1j
beJYs3gqPx0Lymvv042ciZQjihl4aEEwpr95rWTJJWS9ZEw9iqLfwpWLJ6yoUr7c
rjad8u6o3klzhPmIClQJRdOiUPTxi3Qs9RNNnYKjZN7bYS1kXepC2nMXXfBn2tQO
jer+PsNQQQZ8ElJG0/Xphlz242hAyB86KjX4F52CAjmQiXHYVtgWzWa+XtFhKXLA
u/yImQnu9ct2TjqIRI75t4szVvcU22iqoQSZcJboxb0hwZVtvKbP8nHykuNy3xXm
MCF+jgpxIokh6+GMif6KE7zcgbaM4MdXdOQSWq3nm66yHx/dOpqi2spOova2Yjfo
rM6sShXOFfWg7VluQBTI2g1PtVs5x7Dyo6U7IXJbweQPXAnZ0uLUO0f/khtllbTw
vsC+xSgVOMGFF/izjhu7K4z3OddwS5QkaJ4Xs8KodUFRkmFKBIrVoNt08Tz77kTn
B4MOYN+tZsxZpb6Bo6HESgDk3hJI5IlCJeoYSZYEA7EvV+1rENUlcOBROVPXdAjS
HBoA/W7xMZQczQ+7nQPc52Dyuh5QFlZ5A/td4U37MKF0MkSk91Nm6bYWhAutPqT4
2WB2XLXs+lJ4iwx+4mk/rUntjsexMBRLY/COhHXSlHuZXSfQw4GSPhgbP2adJO8r
VBfzcHS8n079nZgIvYkkh7usK+NYBmqUmM/Mji65/lwB70uvypj3orTfnJhnRZ8K
6upXAKFSJ1mAhO4LoB43KSin+ICWdPB2ANWLXXEc8cKVFhWaN5eYQANEfza8W2Sl
CGlHiKo0Gw++Xs6bNydPF4kE2FO0Quephz0iYslXizq82q4vzWhVl7g+CmEf1Gom
yckmcQjexD0tTiF/lKUm6htos4jt5lsqnCOFI2pCiFckASMy0rdfaYFHImonegTD
begrYt7wgL9yBzWMj4vwR5uRXyPt4IrWg1uZfYKfy2ACmRIkUEWY+xh3JfJ6pAC6
M4865mLoZbg4Jds+PlvEx0xMZ/AYt+/d1TFRGyGaAuy/igtkeAuuCYGpUaPkEWKz
6eZdelPsEsEX3S7TQ0bPpeHw56Wfus0aExA/cLDA+eYrToklZ3m5YJvLyU93e1qu
bDWSVz80v2zkMkVeu3GubXHFaSHeaKRHX2xMTwrsJCyO7F+Ju5Wd2k8Izu120jTR
hKharE0Gwcbq3EA+rH5DC8YUfaguM2MWAOSjPZtPpvBsrMVgvMckji1pxuatsbtt
m0vNOfIpfhPNDm0mRoVXn+UzW2aUL+TJrDLrwhAjaiHmSYlhxVD9rpW8s4VQ+ScT
nOUDFzsfseQ1C86280M/ef0MYNxPVvtU67/TKEUsRtH/g/tSLChCgmXrLaMy5NU2
iW4/EUKkZcRoOwA9bN1SDSrT3Q4VY8EF6McDgevKytkYi/3XXnoLzocSWgEwhzpz
Recq5kXeMv1IlmxvQHU85cUs1MaH0wstKRxQz3zfKs41GZ1swQ+t2gX9Lo+mMHuO
0H0A8xB64gUHmC29Icm26aDeIcv1fZLdwznwHHUMzJCmdoVCBF8aMPHlzGFBKXfm
TStRJr62kNLjleZFiDvEMz7SrA52HsfgsEdtq/4UQww/nSACMrpNicoRSUgIWvyh
rGvq4OZsIAp0C5ZFqRDP64PEPoJVnWyT4HoX6lEjbnrSZ1hLWzTao3bQTRnsXhTW
x7Eu42sVqxfhFji2AsyxTEy6SSi67evDxQ/ftatQoWRaq6IBfWk0Zvad+PlTAe81
oSQ7r7mrBbehwHLUmix11grT/YimA+bNif7bxM+twkwkGhzh9EqH2yhjzh5DQpWA
FcYfOOzKF6t1Nwfr5CEMXYG4dy07UcJAQDXHGXf+eSfHi36wO+C+a9+cagTws/j2
/ajklfYmqCwyC/N4ESBtKOPC/yFi61URK0ZcedsbrqKSjZJenhVJ+nFfqp0nDVGT
ToWeLHhMn42Xd348Iv8QFh+Qh9kD/+XIVLpqg6NwyunmrClqawsEitJN3cI1sbCl
GX+Jo86gkGk8aAxNYmbPk3WZPQrD6vFZ1BnG3C9rOwkE89mL0p+O5OpTVdz1n9rq
qoAepGzb4EA6Qn7riV7Zz6PP/CXV+dcZv4PsRuhJuCpMeBLWjkpGQK/ValXv2irt
ISbc7xildOEkqujkzcy5O6oGrd7cRE9oXztgWe9eXvY89CDFS61M0+I3zOEWa0rz
nKkM2nkF7wUqJJZd4Lml3/hQomWTHD+co676GaoT9Tr4TkfpxViv6vTGD0jlBWLK
aHSl+fHLxN5foguSNijWbI/lQG62oWLAHoM5DvBJWuQRteIVkmRtkLV8rUpSuf0+
jsLu48cgZJALCvtHRGsAcrkosx2ZUFSTtT5/dzD6/+YunGmcWnN3hyFre0T0y11t
bvSPIban/bH3kGPPPetGCaYoRBCkG2BfQNKEHgPqfthF+es3Dt4NXyninwX6Hi23
dyWPMsQKv3Pe7VyuQ8k54/BO5Rcp5AHQlM0MMjWbAmteRWpyy7t2EvtTmiwQxR53
w+kvkoJ1Scvcix0lF83c+PPlx3o63HQ191VezG1SRGRCtL5x8KFGZI/p7y/eLJs7
JQAVG8bDuotV2tZgaXoabjf4bThfUsXNO120ZI7jGecf/GB32eaqsnyxq+79aehf
CDlpDOrI2t4VbXvzJeAnAnAbTIliy5tcZuCIZaZMmPiu9PTWcmd2GyX9FlKzTz1h
UxaYr4yEFqbO/nFMpGjoHdInXwxfxbicDdxYub+PbQCB4ug3Z8YarnIeRt/XKynL
6zC1QEtEnt/2IwCsotD3yj4oSwg9EyqS+jeE7JigsxrxjbTsBJQMOgAABomhBtK2
eyJi4e9lUCKNVKJ2zaE+MwVqCHbOD25l5QnyNe3SlDEc/1zyzy7w+mEjPwVhR3DL
xpCDjJk6wE4KgpA7l+nti4UPQ2Pqar4eTRPfLi2u5yKShEYyyCz6j6GAEwjwg4gN
m68Xc+jO61TGY8FTR4TRT+bxn1HU+owsWW8yWQufsItEJWqWLIVpdhaHffUdSpoS
Zd6ACnRDOxZPEZIALG5Uo9giJKN3JNL0UfMih9wsgjEjuqWILKLexTnC+21MDQ2Z
61srM5WW2UGhqtDIsNFnVtds5pYUFI/gMtIMUaH+DX13l9S3UVdRf1kfLttBlYmH
04GEvSoaR0NheKeWo/cCQ9d4BNU4v7dtbqhTERofXSNUZAFZZDXO1jx2N9xqDGjZ
+DbgxFId0UaNeOOm8nADukeojcGA9+fQtw9ApEXXt9VKzvnjdRFFVa8siKXaxKxS
kD+5EfZ+tjByf39j0+v0pqDNDLw11FYngRodOBapFcx4jNShRUGQXOCTUmXfsD//
W9EXFCdaEviN9KS4hkC6BegaGzyaooLmT1Z2T8BEU5YuagZ5Mb2VBP9eRyUor06y
XWg4wii+cWEkf07seuQkuXeuhLxB2nGB25wwBY2c5QPpE9nxv4VS+350gz+L08a1
3ooACFQpgZb+x1ohlJMQlfRajf0RJLhgtVNZlGnIpmxbz1YEVwFKu/Qz3osuk0qg
NUU41Id2+amUXLr03HJ3j0lJ90q8oqEcVu1Pg3RYN9ztdZ4be4KG5Z1Kvmg3O4Fg
xxtSCVdQH9RxiOHT/OK/8sOyo3lPAnML/PC1xNU4DVUATyA4f5W1DWXssHI3NAVg
R7R04sPCU7fwFN+0OSTLnYR8qkcnhrjngnNz6OCtULBpbvFhsmFTAzr+RamNhwAF
6fy4A6kc18KybNNSY+U28c3wv7HPSlPP9X9ISpKIoA90JYmOHb3TfiZ4Dr6k9KM+
hFGsRiqeL4QJQTnpmElHzlArRO7hBcDz3XW8PJoDi+KNHchXE5lCuKUWHO9DIBUT
S7kyWdWwfjREQvtNTEJBxE8hmxUZS7bNMFQ/8pckXvW4/l0HysTp5vEajDR2c9io
uUyfTzH5QBBkNAa0dBkGTc9miR595PQMmP5o2qS5zh3VP4YV7ZJLOseD1FcXHlVA
xBb3Q4qVLASgV2Z3fMz5tPMN4Em5yYYwMz8qjRB+gWR8TXeXWDcPs6Z41AldCDyP
nsmP3M7zpXgiVORX23yrRYC6K8vswTwfruQp2QC7w1RTQP4uAwWYF5aY70tOkJtA
9HHlW9uGBYxjLXxEl/Z3lM9hqsXsrs2jwu/NiK7m760hcf3FGmsshQEBJ8MkcFe7
k9olLeLlTFhD0hY1S0TDNh+i6AI+CbOMrW7XfM2QfzHRlsfxhEYO6+i3cpPqwhoC
YbOs8was1mWIXwN1RTZJ0Ws/7ABSPKBCJPtWK0Za2zpkK/e/tbYYQA/W9NLUj0d+
yd6VSGXzfovjqKGhy5XAvHhByUwQl90otp6oZ8CPxJOjBYahmKf6RpBDfXZyGiKM
l78FsDOVisOorV5G7fRdI+pr38eJayUXkDDd+eTxuBW4PtzyrgqqAUhYJqrm3veY
h432QDluYOfspmN5pG4NbmwWKa+ml3Cl/4LLd3Cr2hDehUMxd0MRwg6XWPr2qEXC
634DGE/4bsRc2oVs5yfUWAjmbk0NgZK+bvMVVUXmSddxoPdaEmT6JteT/ypTclnG
ItZvS8k0EwSkOUG02vaf4C45nPzY9aYnzn5pX/kM36q8ykxOyvt9+oUvpsEtWdp3
18c+Bye74uqAN3VgsptLmBMkFlwKTBnJOFm5o/UYJ/wjOdbupr0DIqcFBVr8wCKq
mZ1esPcO/HK5MyUuwrZ/BEwZiLeqxc4nQojLir5BQHFTP6CSR6LgfvRC4MYpMQpv
DURrGXc/bDSfZtgk1SHdyAfHoATx5u+BI4AZ/1BXQhtSrwJBjo9JEk09/huG5861
HrHNw8tV7NWb6p1nQ/PXl3KT7lXUU4DMVzCGXBouzX7xaLtAdUHersA4LOt4MqX+
VLZUPNtqt4oYGmufAocc+g4Kb8RauAzs7de1NeI+jL35NdEWPa12GgMP0+udoq/L
0o5mQetBzjIB4wgJbgxrau/B8K1NlXwdff0S3DL3Q4rxRGO5hLOpnJvrkyq2YHNG
jwqy0gQ6vc2fzIDna+1R4KdMoWf0Q1xf0vy9OtQaA3g/IHIK1p0youhDiqBM3mUH
dhI6SxJ4IYqHy2QeMesEeP97+9hOqz1qPMXtSY/w7FK8mc190mUJ30xhNYcfywPb
njud5FpArz4mVj4Hv7FccBk3t41wxw+uwMfp7zoX9aJjnkQUId1De+z5Q84foA+4
2h2sypXnyiomENB0iJbNoIwuJpzCgv6lWwSIz9A6fE4NTi0qvQLsoHCtvheccUJp
umo06LmBcYyX6UVvx778NQphl9X3vxdNK0hqOLwpe+yjTC3S7i0Sxrtigcq+o1lq
E9TIQMmlh/7amY5qyDqDYv797IFE9iJd1Yt7CwXQtCTQt4/xv9SZKgvnoGRYZJHN
CoLqWuO7yqckwCcouT/ctPE9h3P0+uFRcy4oWiv9HrH9BlhEmBbyBsjvzlM9+Bvm
JYTt/8+q+EiyPdJRC0ENF1YMf3kR2DfR0JJHYS9LphWxzf2bVO6UaRFUcDiRmgNq
YHetVtBBWLxwcA2FxLajBdFLofcBx1Ryc9XqsOv6md+oZyu7w8GhcMeaZWmSe84A
kox5sRVSI1dahBsdM0uE5ATZbGGemdnmLQRwThTQ7fk0ANb3Gk9qCog6z5Hcqi6W
ad6oYLtfPWv0LqdtfnJEEWoFsLFn4OTKaIhhjfytunCYyR29Hmd7hhn89wbfkNRB
gLVflwtEzYPIXIRARFFrbX1cB4kiIqoeqU7fxee7GJbZp4ovi8RmsR+AZnqGQ6UL
eRwVkE1fuyCMjGqGYXjDp1ylpOx6f1VajNbjWpFQu3eZVAi1FLKtp27cOgGyeOxN
8MLZUnBnieqkiloLj0W83EYjbxAawn1xznprJPQ/dUSnKGyf4MtxPEmkx0hNOTBd
TwFMWW04RRjiSuAbKwvs7RCU+qHsfNgzU8+bCFGOsNsQ8doWNtGetCeLRNxiVKzH
mrQIdNsNIjeQTVLlQexDbgNFZ8xpnpzJR1WDEfrXl53Jp3lCCehGhSOo2I5sRY55
Q1pZctK4Ep6QteVYfdAfSmqDRThF5OgnzWbkLOodUhF3fVakJb93xbtPARyK/08W
jXnVgq8E/xxFeplE1mXqtAE5eQL5BN+LTxSiZhdUUQXRboq4DpG/3S+2fRdeBeTz
DfP9MWXiLqEdr+Fu+aa1h200qlMd2Z5uxmANS3KqPVFGfEtGJucAMHO292Xmxd6+
9z/SIPgIzXLYUjrPLe6R6oGYlssdDHsfYMliMGTKg79Ab8y6nelzIpmjYQSZboh5
LLonTT6TFBog3Fn21KZzOOpuhGDEWIQ1s1gb101RwDIFzyosGm70Ut6B16UEeN/l
TR6iyq3aInw9yiO8J7SovEAINZXg8Kwrv4mRXzneH5nQtrcrvwsQrxoqtY8VuL0M
9jhJ0Y0WMMJNQzF36LVpWt50eXM7dR3dfEzzE1EzBnmUDG4+0MT5ElJx4z309BS8
3PZeFlRM+zEyeaR5qlB+4ndZOc+1MW2DW0c8dUxrSK7i8CeYpYNvwFRrVQAOVkCg
K5Vn4hk91j3GVqiFr5wPaY8C1t37HIeLJulRN7lw8MRmeBTnjcB6g8RiC8p4MWa0
WCbWZJC4vnVkV9a68H1ebn17qgUGIditnYvgQb8ZC7qTPIxi9qXDEjtlc6sdpLGF
2nV4uy6XqQKB0xBMxRjCZyau1Oas8CIIPyct+GXW2VHt0yRIMQu+xvVgYyEpQj6d
fHIvHZ49JVK93T3Q4TxRSF7MrPOXz1da0jupXtzJXiHg/dY/UVqLEZJ9mx2fz+Z2
nN7upu0/k1D4k8evQk+YjuWGZU3ku5Mg3m37CMDnlAgQAa/O+Py9OExL7JISNu7v
UqAfj0iKMGj8I0DohBGhFEN5O9HqYlv64ogj3O3JedaUDQhKdrqjP7fTafkOGT3g
dK2cYnPft5ePTujobuI7PeJG/iAXLunCq9KQq3FNFddEXSlfykzdllXDZinfBWy7
uzvnxz2wfuCXAKFu19sreiKaBlQs2c1uKZFyICfA7uQHgb38hPyt4i9sFRs5DLZN
ewhRHmsZUY73YSu7S7m/wsT64QxvYaX3J8TPkVRHZyBPH//GQNtdPAqkSxXFD8Dd
2jOP8M0nG9dUwaK9S6CMXQmBEdYHFaDVAXBdPXuTLlrYPr82bPSTmRCBuabA2SMa
8GoQn7koy8OAgBq3UL4eXp4faLsi9vGB18GS9kEbhmu8cXxuoCLURKxm7nSkblLu
T48k8/dtHSNC0ZKsW3dyM01fsdJCfC4q3KT8pIC1UEcxC+fOf6VtNMfYl58j9I1j
BfOAFfqVFuqO2jXAJgiyt9O3dERvW4P8DlgLd6COi01Y2c8ETSgg7fOkfWKz5bXu
m7ef8pjbn7PFgaT+hRFkYUNtsbf1hgYX7HuJz7HHsxHlOEg5oUlsBC4ZKH3awEXC
ij59PAu8LmIpDb+mg3kUiPDc8j1PqSYPxpu2EpsRsFejarA0nrXfi/EgVRxDnEQT
R1nmuq6SWFZgKt7knPbqqXgen24aFM8GrSqHQauD2Qs3PthwBjluXNLlH+fYwe+p
Kk4YiU2TkpBMSiyBqcFsrJhX0iZJ4DUqv7fkYtArlBDy+a1di8IszNwnyDicKrFP
Q+4rWIezxJlkTkCgoHrfgmvjgkHZhltPe7nxtaLNhV3NWOOZlY7VQ/ASVdKdbQZ0
L8aW4DC+AebHHgPPy89BA0ZbdST1+uytefaBWUD+Cs08kFEQtNwTtkTm9Vl4MVgY
MHA7mKpyiR+kiYTni01xY4ZRWL+giG+aQBHP1KB5B8yg9P8URglGmpT5bWcMqDTj
UWCt/Ni7QoxtkeucXslDNvxlcc/I8v3aqmY/HAzZyuPsu0dPcsuA1tt453vH02ph
es+mNSqHm7BuJRnAols3/pHeI462b2lNVWznFgibO9yT8+tRcf5SCYDXkFm3Y/QV
qLq5kOqf2du2F8s1vzXcfKLKrM83JmmO/E17IUh1E1qm2pcMXA28iqtszoZOnRpq
pudmd7g6MYIctBUlNAea4u8oRIghbOcwe4Q0fRMFum4gYlXzx/Yz7b+pE1qZFd6a
qj7WdfqN3A8V/0fggF6L5zx4Xz0zQ+vBcyJffniT+MI3h6VyQ/WkywqRzDvUDFS5
LK27iTooVx30PWcR1Sgho7i/peB3xbptW6Q9GikcDDryFjwRkFX4I2dPkp7fMQw/
7jJ/iY5qGDpel1l9mPSDvtFZb/QGM2fq2yCevojHG7GCFEgggQEuewgHfYxb74yu
6AyrBzTcVtRkPUvu2yjeDGFQocalyjWqFinn08XlI7Tiirz6hui2PY5RJYnkW3g2
tR6B2cdiOXoEcYHvlfM/r6Js/bzewI1skhgPAw++O809OtvKl1vk8w5UQEu+tS/c
sI2ZGvyL5LfNWcpJRhSyGelw1SHWPCjoYSKRZjIs5vffQOrsmLZOMcRl6MCyqzvr
m1wkPskKWIk0BzCVFvPYgAV2JBmSU8P9ezyZ16S4b6RvQx5BenOy0Ff/YvX0JRg+
scr9YMRsugCHaE4aKNylHfCXXH8fotGNMLe4HVZWkWetXzwuaDF8sMQqaYzfnn6J
h97auyvf+5oVceGIqLtpLDShdWgQU2ckFeAcK2mNTZQwPXr12GPB2SXTGeFBNYq0
TE/myow7C22Zj/dLIL8+Ye6b/UxL9qFfQm8TN/TjnQyxfgRNvSsQjitCAzV+UcEk
0Ilno1TFcGyGg781ZDbN/d52zLvAgTS3XgibmBUpWqH1smC+cmgdpUKLwQNTEv/+
Q6sj7o84jrForZ922rpw/+m46dGoV9qGXWfCEZXUmClct1HXIGEuKmPtKV9jrwx3
UaS4pXcdiPG5Y0XGRcd0Me+NFwjxidSGl+2dvnyJft+CcRVcin3rx/pOS7ThiG7h
7oEBJNbRiHXQ/Cl04Utq1rdJCzsHbruG7gynWrqhvlyOg4CBkDCwqGTqZOa43AtY
pyt5Y2wk+YrbMYdZG9kCSUWy1g9aGFTa6kG0smung1GJ57jSCjCxybwxli5pJbXV
P7/H7afyX7ut5pptSk92nGl0mzXYe+WXLG6TcgNQhJo/T2LXKcBB2Mq9b8A9RwOj
LJGoKDh140vEy6J6plgqsR2fbzXDYDL83LMH+GMRSs+VKsUaP3vJKMTTJWrvCmvy
4Xswo7KWASua/O4twB6pEJ7lGKeQgsjHMfQ5aeH7QpvEkA3rUO9TI4U2EK2gvK2O
8rmfSoOyFqH2Da/1iyoHheR9ZNB+2OUY8dm2oYwdD8Ui0LoKk9CElYDKfdjE6mpU
Fm0xlqDtb/0mz/x4DIu83Ie9OBpzT0xvyh8y5Pkoiy+vOJquYhSgVVpSlUMF9xDP
Ti5XWnOZkkCk/ECZ4XrDYRhZ0zgy+KI+MWSTjoJjI2mUozolsKDnnRWUCoDEeYfg
Js5yPGhB8M5M14qYUL05ClE50U4WBKLAYenp+WCjfFn99LBWn6ih6HrcD5V73H4b
X8hICCWt6sQCc2VX6mzAzlNiuCbmcv6q2XjzV2wh9oWvCwd6kDl2SFIBe0qQoWBI
yClvLz0A4R9evPAUzaFA4iwo2XA+CT537L3H8zhKDNjEPqyUtthHLmeHWn1EfkCg
ub0XfTjjxcKna7bq9rtGtzgV0rcFtuCWDpMGJu9dAV4T6EpGXgOTKmjEtIT0pakA
aphEddlhGAGC2rSrSxLrCwbgGoq2SNF9K3NDnJn/ItB7lZth2yeIwTetI2Slldl3
qzyaE4Jk+hpe+UwAMO3T/0mgO5HU7MJd/csyTpwPPjavyqeCVJ57+DL39lNUZu6R
Szumx0eO1cq23B8+40aAidUhaKVVOQ7yCfIZfJMyX4e6VvgPLj90eQXxYAYzs2hg
oveRwz1LetySYMNYQGwZvdN8Pg0I7VShVW5XA/XJbKF5A/5wddUa+DQFoMrwgdHS
cys9FvPpMqVhR+DpvSfzvP65ZELYveTnFTJXxJAjeJurY1SkX4I6uE9ov0DxoL94
Cr/XxuxksuaPUzOKIRCJeKR+F+shyq9nn9TzE/mMUUr2FRhlM4XLCRwIfN0HWzBG
+aLThstv2j5dKoxLUaWQM4R4IUhvoIziHce/BY0d0HjDMMRn0B5EbqV7/TL8X2LO
ha6a/0f23Vj/SJGY1wruX7SHTZwwDeALxIuCYzy/Pvlzp0+1BUTq+pRUyDaDgbOX
2E0MgaB7DOecDcOBbPfY4ybqJDCvKXgVqgKz5/g9C/I6MYpY1E0Gv/XWfzHcGtJf
3skZNtaVmi98ZsEZ+Xo3LzCUnkFquxBqa7RuguDhtyzMwozYqAgBjdLeCSrHdu3T
NqEPUwYkCHrG4X7ivpc5NJJpl6a1c0vBVOum5ZaNoBQNO3DF95PdF5nLXKFdh/DS
N1BeZNTUV9GqOJ9SojvRJIYFm5hEYVjSVty2/+qppYeQuJUDFzqz9gQ2oJgzuh2F
bSRShzPtcgr3XmqFaywn/Nqfq1/citD/4IFri4jHKzbg2j4E0mf4iemLjtWv9UWx
xXgNAOvKFpFlYvQdkL84An+06CdTihJTe6mn7SC6A6AvBtnStpLdy9lwS/u6vn/Z
395izV/Y7lUWdgT9wUZRMMPpcjUt91H+6arCyHWK4HgDlkknZMH2TGJMYeSIPoZc
L1PHKKnEfGBo04QPLQANRK0wY9LLL7ayHLi38c4Tklj/QLRbWTk7pjiUdeFrBOGJ
UXctGhA+qGIxqu+oKvRwki0QSzUn8Hj5tWCleYqx8GFqhHo3ukEc4fyodG258C7G
vX6JTc17aXvcMKlZsde3DVnnsWMOigpkAtXet89zliZjQOJ+nYNfPQAeCs38fdiF
8CnGIg8OjPzhlCztB+5Jjn5BSXKhgM8XSPCTgVxg2RoSAh0M6/Yunn3eBOEbk7Qb
vPAr1uKXZZZvhBWlSk0cNFzjO89zvvQdVxpQe1yPcXutG1sabyttK+8/LiPme+Kb
+ShRDYQAV780LgzpFICDgXtXFfRJSZQrJDqw38aitPsX/yi0mWAs8hty2Rpx4r1O
ztffxx8xWOAsp9CdEt7zN7PIFWl1GZ9nDeLX/1RxXT3WMSNimgf3XRVZb7pQU/kH
mEsFGSSACTvA+kyuGx+kSxlTMTr2ElnPrO3quMxtM5XldHncP/zu1Vz1bk/rMD+z
yGeErAM1XXXyJbfICHnvC+Ia6rtDkOzo6k2vKT9h9+MOo7MTb1hXSNiIft29gOZE
U7g1CHNaRUzVp39VfE4W8nDRYhaz90iA6I5XNEdnXYBe2CATUFjJeZhkUQ7owTOs
gJz7EbkcFJdVyLD/3ZffMKwQauN1sXXg5Zkb3aMp1IBYmF6na0gotz/TXa/58f7p
OC3Z5fHPjIiNnc0OrEIXQ7yeEG/vVZoybOs4oHG3IgHdEO0x7D0bbQJfc3ZBKLZ9
xNn5WLs9nPS27+jJN8XJP9HL/Y/WlZTDagRiBFUrMKPQyxb1XiYw2SXDkbmxbDEG
tPgkgm+G8eMhMtzqENDtWUbYDAvtvamx/MLn29guaGNoD+dj/5APYQSdeoo+YTyb
s8MwReCfaPlzjPuP0uwTggkaN8sXBYmFXKMe0lqFrrlra8blZQ9OtnxPvmzcSv4Z
1/XFBs0IZ7X9B6jcVN/GycHAopIyIQeJtYNW87NR4uuBOSXlQvUe60vb65NMkDad
gASUx0RF+0+AD3yGFgP65eEFEnmirrNeh9os+0Y48y6dZ6zso1r+p/Ak+J15zt5I
uOhqkUiDEJqCj0YLT2Llsk7m/HRTehtMiwT24lQRiVT2aQN4sw0awVSq8qWyUocu
In4wm57YQEMlwRPtVyNwZeijIPnhm4Ubs/IYPm2ZvWNtbuyYjNSpKXxv1jN1FBuk
icVQFkvd2UPRu11vpS5SZTWf/9vlTq3SamgBRgj2wI2JcRgrJG9AH0FOGjnrRy99
iqjdP5L3ozoT7uYI/ejrABbNQI4KaDjxRJeK1vMAD3GRpg7oSkfZmg+9PEsla7QI
CMHuQqQeBnUaSGgO+SRgu/+OjFvZboCbCATGgU4nLJNFQYBTHXojWx57yxhd0KbH
NKSLrUAf0t8TSNng9N37JfAIDnrkZpA1le7koAFMjepoMqkBotl/yEnTFTOn1xnR
X9xJK+UGM7lLJCsJ09LcV3D2b3P4ZfNbkQZKsGLzV7VHPL283yE37D4VBu9hmgXE
6e6fo1hSWStmWsY9yT6BEyi/X74nf6oyPtIj2fW17qRA7UlR4lKmgc7hIJnEDbzK
3riUqf6Ozv8/7Q+VHoYc1IzJLASsHr+Q+rS8Ahjr6KkmlGEKQ7hp5+bjWVy28eOa
suNrkORwRRaorHZNe2fcLS0nZgrrEqD5s4Wsga8k7SxWBbVuajZMFFHBJopV81j9
zPkx9GB+lV6yF6Stp4qWA4muCQQ2rwrHuD7s/XzWA/Uu0HSs01mekjvVh4V9oywK
7BL6kHNA/QloKFsXJHQgw8QueU3mBoZWzP6KXsEAE84y41isTe0aEvV9R6GrIl6b
xQqLy80JD54Iniu66mMF9IiyFh17zTR1Ec4jxilyIvmbcgsMYBn+M5I7blbQuQUC
upyYR2X9f7PrehntSpR3xTyH9CciKf1GpwLAdPLmfBc3dLUHkgVHBJUrQxe39wjO
3Qu+tnO0p7hdIzvDoq9oVve8r+/tZ5h6XhVNiSYFj5+C7rRaxj2Ok6arTTmrzX5r
F50wCY1LFZFEIlRwAHFvffQMiXx3XAuw+RsOXAoTENBvt3qryN09PlgPMVQl0c/2
W35nSs26Zk3RLbZFmhvoMJEstLqgkuBBkIy+zjVqNquTcpdjyg4RsaYasrcFgy0L
Ox1lrJ2+wZ7LXzxzscXafbWcbSoiBB8ZUlTVsoOQGQ5MsfG4SeibHhXWVtLS9I6c
amV8K3dybV0vgkGW5/dGthq3F9NXeJfo0Z1Rw8mOIzZYeX8RlR0J5H4JDoCMVU/e
VOLwA1Sonn6NC9fACjQs7soSlp4amXjs1Cq7AiB6CLiyqEHzjcYPtCLW9IclOwnj
HiYUowg5VTVCWnifKVWPKuYuI74H94c+MvoES7VJupMM7eoUeuX0uCwkcibWhUn1
BMEbIAXVy1oCd5xtJ7AucTNV3Tjxld3nhS5kbn0oJbTVl6ToOASquXVEonGlzJb6
G+HvUYgKTvq7o3A3xyU9Jlc2PMYRqzxJ/N20KzLhuHQU0cE5PLlFFKgNrmo2VD+B
KypYWySXFldgSKbq/P+WJPNEN6GKrAnUDtaw04nUMIa32H0QsTWA+LZjfMnrHfxU
2ATqNiegU/wmA4e1rBL7uzuEkWM4E3yn3SFjFZGkbglrmCrRyEtlFgQdH8GmayhH
iNTc7U9KsXj72v8Q1CRyWH59NYZRgv4tzYkBj/CkKk73tt5NeCmIF4mjDV/DoVn0
9zRnSatP69M8sWbVsBuOg0+4fPFdxNhuME1HbHYBgEYZUTgXp7qejncLPCglMyQZ
0xvDKyYvbANc/JOzwcsY7S41wzGZ9YPcKl4yyHK5xOyFpub9bssdveoKQvxLvQCU
i2lla1oS92qyr1/oxClGMIg/dNbb1JWPP+yUPKlbYNcsBCuqaR+O5ibNY+TwbM8f
gcPY9AjhrkXNQOyy+twXqSF+0TmmOER+SBqtjxuNRvlizCWMYuL1MytcNoi8uSKg
d5sp2CtI48Ugfoi1x9r39OVCDE28wGS2xPfVE3MWU8EwFDvNd9ANBz61xRzco+su
HHmALvDDVMv5luqamentfWtwxGq32m97r7w9EYJvYADaDzOHmYQQjYqL+bRd4Wl/
EKYJDcQBIxdjjLhZSkZCmZ2AQp0v22vz5lMuy2s70odp3F2lWX7qVLbjJNKm3Gte
MjM150cqUo19YB79JRA3sgqRr34HPhoBw4eQHBTHxGVm7IcxaAadzsTGQGJ78MVv
qdTv8F1+p/tfwbngvk/9Q1KZ47rRiBKwp1JsXyHMb5mDDfSZehnFSH8nSDkY0Cg7
ZilUO/2AhnL48hU5xWvYJ1l7j/SxKbcEzUXuAFa0UpGnHteW5Y7RhyNag/YahW2L
9UoBTREbZBVGiTvFA1qY56vg6yaUsZbYD4abVC5xmvGhdoV2u8oIdX7r3FwUtf0K
1DKXlWPLRliOCLHDGEQbiebSr/T1DldaGqOdFcv82OAc/lxfssyEucAxEC2sJDTI
lhNRdSwzeEO3GVJnowWHATQG7uQUxH2b7wcWBDHhDFf2sgy4zErWVDYXBopCbuZq
Dc5pHGpZvsaVDu+3QltV2fZybTMOuaVz7mV91B7Pt8dk+l9sFAtq7emusTDLCeYi
+vwSy4wRe2TP3ejYMr2Y2EkCd5Bt02R4/Z/KFS3V8yWbAype8sdtr7SgXaIQxwxh
M+Kbon4KuZO0t0CYx/suWHTw0v5Jtkpb2nhYqOKiC3GgfNQCuSxhXa9sEvS4cW8L
4HHP8oRu1PH0e+6sdgdVjYr0LzzxmAJbhecDbhWitI6p+5KHxTg4DYBKZny3jFzj
RmEPK5t/xvqPf7eAK1xjz6/5JxlCgbW74HPsVcXgREFquq8fo1VFf4eCr2Vj5wXQ
IXvM9DFe9mGuz25TscfQxpcPjdZ3AINsMbqE/KnR6ikqhuiazP8vJ6eiV7TFbbwx
5ziPTlmhFLQxUNmsauLhOifNJvZpGbEHyrkSEV0FXnjdJFwjwkx76i40ApoOu2Lk
Nftwo7P1msGO8a8aykMFK6+pvuE5qs3HaZzmoJ+bj1wVR//jQKZpUqECRbVwpTH4
xsYo+SfqGfx/TA30p57tabEPWU5rykwqnXkhWe6EBVZMIsMxYeUbggQL7jouMfrK
NZbi3XNNx6FOCg3Oe/8f1QWoxc8Ioc3ptVFV4FFEmAW5d48wv8X8it5XvPrJ3cb6
7MUgUQNwt39lhpqDJ8flQxfrcRsNeeJ9u+1zWZqOJLu153Glqs08MjHdLipFYKxs
LRcNGqGnM3nASGqHeAXH3qYYqBxRluS2yD2s5ToMWW8BHc4EFYqJWzm91AbxxaY8
yvuSZJVtY0pz8e3vMLO0G9mPYEU0M7BO6nIIP1E69744+1WQVrB2QMuUcJ8hDSYa
HwXcR89oe+RV5SMK4YDwx/To1C7y47tsd23/THlodPmUkum6DR0FV/XF5PimP2mc
AXgOzxOfoKo5PpGzZZK3empoTtWtxSH6xfJzfl/wbZ1QD9hVKrOd6kJD0tU2lC+w
uStItqZfDDhsEKSgoGPT5rsbef2mfA43nXncnmLy9hRQEDkMntX/ZR2CHOKy6360
PTd3vwAmWKCyWZI5h/t9n3N+h5YK1hIBtbvl/Fkd67cggXUNOvKgWXmuY7R8GN9y
F4MseA7sJarYAOlbvOd2SHnRNN8X0kkOP2JG1JIMXIii8xzYeQwUgokXal5oz/WV
cWGC68IkHvCphD9UuwHxDWvycG7x+MYj3pgA4CJn21qWrUfFE8/6zVTmLuJdMG89
UYNvc/5SFnExygu9xFi6PUqBc4BMe4lzGFJZGrzTthXp7iF0bCLME+IiM7trszAV
AgePUVSMsJjgAQ+sRIOFs/9KVq+Tv9aeCKm0sBvZ1Cyh6VJaVi4I7hR697papXdl
erPQKY8ldFQ6sYjk2cOjJaYqaImL2dh2BCPP6LmL7SVxXdrOgjotbNMM5XVZ7JGK
njRYyD21mkUBhxn/vrjD41T5nG6js/hP39lX1ZSaNyBEYvN39Uc3az5dMpXeGgBn
uQsQUt2C1+I/Pk1A7d/3gHmWRAahwQYlJPZfgmaFuJiTsDMDOMnOMlWcJDLDPQWF
qjXghGkp+TSVuCjSluBT8RNdfSvdky0UvZcW/+hi9M/pNkEUPrZINPLvPza55YCx
4Wyl5RwnsXtMQf5KtbQsDcNwe+Pn1LT1oLnZq60uao+Pss4OPOVR5hTLBAqOkibp
0SVQYzVq01KGMYg7H/GJWkgkQcifUhGFAsB3uNp8RyHSsJrTiMLp+AH1qVHBa/Go
TXooGXfAc9s6UG/mswjZCDdnbrg3VQ2CvmqgxPq0mSUSJchryJYElYQtXQPr8x3R
ugQPV204VqIOUTmDRaNnbMGNmEAAxQUtALwReq0vGINX1qI8+b4z4RmLTFohZvG/
gQJJzu8ipMF+hSrBtx7U6fZJ2ZBvkTjMeU1AqW1ziOJ8qTmFnI6rITn2pexDQg0P
5ZsSWsiP/RKaC4NmU7iZE7NtKXIpwNIvIkcfR0fghVPEcCh0scFh+4DYwAEyoQYl
7vDwQdacZUW0rwGhuKKlrvM3VBcHP569KFOr8HXEdoaLz7Q7tJ7rqD//GGoA0Zqk
C9l68Mw76gmvIXaCcykBUk2G/WCnChsTACa3M6a/yz5C+RKxrCVxgLINUJcvNQ3R
YVXZHZZT/Nk7GT7ipGnGAPztMRknwFnp74qoA4C/i3bmRjjEc6UXLEKCPCb3SDHR
z1dUYuPDHAMZrFYDk6kjPGTxXxQHx6QCwNgQl0Hl+iBI5BXswXrQ/pTGooy7KBtz
HO+AlzDRazhi+qrKTVavW3i2/DmA4r9tH+/VPsdebNDGh+3+a4sLRmU47m/JIjdl
maYaHPOCcE+wcmKpmwDWz/JUtnO/XvLK9qFGDpUW3oSYGLTaWLE00UAA9ynsBulF
VRohg406w72h9bMAsUtA06DkAg3ONYmaW+yno9Uf4CtAojuTtoVlWE6uYEmi9nsf
wxcTyLh2ceHfQzDsXNC/mCdzY2+KithLWFyK5e1MAgU8GCcGdxPVceP1pHpVVi1H
62C4Qm3rM1eKLgR/EPh3+ObGW7HfuyH24/TNdENVzkF+fLlLTLmN7aK3f45SDXKU
irnpVz9Z2xIlyIz/OwC7DDWz0+L1c2LBAcjdhJW1VsQuxaQVQ8mqfjIXiYTwr7pu
8KUDjs10jtnqthXO6uMOcpYbcoI52yOIlySEQyDaEtA7Ylz0KuSDMppBmLFNxfyy
Y6OeIWiqSMKARj9EkLFV2JV/8FZunuKMLKWq1cJ/PdEI8cvMDzyUSvu+wq4o7Nzp
ZEghQGMPoNV2OBbWHf6TYpTqdrXIXQqjsQpmJnITDgUgN9ZmxK0eGjhZBQX1FPBA
bK0lcABP+TdqwQHt8Una2RNsh4AC7b4jhzQsHVIjMgAw01cppHlg7GueqZGVkhIA
skS2MHVA9Fhjf4GazJUBghHw3/RMl5e7Yx9iifUl/MrPp8EfE22vL6vf/yzqdREB
hNtO7JgFKUdqnbUX9VffLQ49KOG6HWoYThlDLpuRbj2uocKHVFk7N5v7wdpgtYg6
VwOQknMxOjz9ydEA+ensiIFLuHkqXhp1Jz71B4k0QG6gFYg6MMr1Mu4TzsvkmQIs
HzRkWbuy0AgZYYpcEJeHDeaJZrehBXKLtbaeNEtbGblzcv3FNEeyZHw7ZB0GdF1v
nttiXs6dRoo1GTlsfNqt86GjUz0AJHd1Vdlb/yUREzzJlIBIalnOryfw3YKH9NXD
BDRR+unUOCQ6bMqhYBgAyc2+YwF7RDuJ6tTmhWjcg13ss+USv17MvmF8eNqSzzU3
wW3jlUnapVGX1YgI+HsaKh4C8YR4T/oy6z4EvX0ntRYiHdUAm63Ag7cSDHNkHSig
r4IaFjxrpub7PI2zLBlns7biKySX5A7it4XZH+eTeDtmXSGpiTu+k65JSfRgUofR
zKwy0Au68UFlciM1zDPocRY2jwnroAiizkS62lqNx4lH0fmGsR7f29wKRdKeB7V0
Q0PkMPUO4y5Dd1TdWbKrlOMrj/7uoFYN+BV9X9NpAElew2STwHzoK7zaeD95j6VH
l9FFd8UT2vv57ZruLPMs338ZMHoymp12lDyO8wfdLfnchrLbYH7JX6OxiSi/jQmf
QHTSzxeu3YZrwDWwL0fP3znlaijDSUhYMNKr7BXQ16X+ouDMUaZa6NTeLOp7fEty
/EMXew2u5/o0kiCXfSEvYULX0yhpWQy2ezmWrAN4AO6kLyqn5G9uH0r29Gy/d28m
tg+bRf11HJMoaGeukc3qvUIuXI6EXrPA5ArYdRn05cc6CRuAaSta/eNsoMIyd7Nd
WrmwlAKWt3On9RSI7ZrQ6jGD02paiY1PucxTXD6nZHIRhZTvOGU6LqwgVo6dVZOc
mVTKnpj3+DNhRrwvd3itIeVxLURjq2v9aKJTyLKBUS28tqYD+DI2Xtz4ocgTOnzA
aZ9FnvNm2ncrBaoc36PlqdUeCTicTITWV0Wf5VJex732I3SPV2oDw/rWUMQ7GFK6
Xb4Cd669gUyRaBhGJ3eNYQE07yuqGxYE3/bPDaXSadH3PRsWDix/8V4SXujDVivS
B/PfqD75SeMAEXYYOJEcFeWQbM3XEHPXI7tGy8ZZ/3ZjsLxxBmobimlq4hQ/WQpE
a07FocqrHI1pZcoqks7oV9zFbmhrZJrwj9RtZBb0nzZvqByNx9pl/NQB+VV1l6ol
GGgAB2hjZ8oMPbWh+qeu/SmmcVp8PRJltyXyI9cvLa/gaOVUWDwKmq2BcBkDixpO
QrUNnxRhTWYLjxneUnFrfiU1IDFIuqYR08oaHVCdkcciiUclw5iw3zk+AOfL+cJL
QM6vcPsB7evYyM3eVp9ppbRIE5y9rewIkDt4yeklibcbhemrvsxg37678sQCN2Bf
EZu6+Aqn5bP4TeSUlQbNk647btFWpLQfvbFuWxoAv5WA2PaLkf8HWTNL+v7a/yXC
VaadKZQt+1rmG1HAxYUC35DTXt8CEw7MihWR8fISsxPUgnkZjB0lNlzdyMHAHV3j
Hy6dfnT5u6qRsR7/q1Ckp2dqmidt4e27KQM2NmfCnV0fT+wIAA7Wtvricu0yOS4s
XuDC9w/fFzUOaIHb+SNnUOgNvQivyyPvncMlxOxkfokbDJ3icUL/9GQvZ1e+JZTA
oRwDAlUTwlbrm7QNVqI8xExJsIUKSY7MNxASL81QM7dzPbdgTzzsNSC2PWfpEC5P
pbESPzhk+iaafhVHJHuU3uPHAnHNzKLslvM2Wf5tFEqqQsmpxgI4e295VVG2RhQ1
QhIk3Tg4libaSI+3VL+j+z7gxbjUO7v6igaZ1F9bpOvNZnBJlaopvUOAw478cYBU
jBbO0KgBycQQGR8CLc9Yqy+lEdn5IB0dCrlbWGBcS5/bT501S//Ji5u9+U9SRDvc
okEgipszdg2SfCN55QEMxTksZNm9PvwV0uKNcZ4nw4RupZLdxurduYZCMR0HeG65
cQppL4H7hmgjOMbfXAq/fMuO0uvOb4OA8dKpfjHQ5TF3GSe2MNjzRg/7Awi0kOJg
2hjWeI++Fvo4EzcEsNmgDo6Ast80MOApwBJafY62zCXCMz/vyAqQrncqxTu34NRz
Gg3bDqL5HlRJshj0vJolDDlIWYdJBSe6FtbcsrZOey7SrNN30zTQd79gLk1W2y3j
bpwB4MdWUvqNwIqc+kyMcTpRsRRcShGY235Ysi/2uaQZ/b3LIyrrQuVi2auF+eko
oJFQ+2Mts/iIEVP3HbwIW8YQgnrZ9g3T9KfFCkjufpsaMX/xhwGhMcGaDWCARy9K
6wQhkfqeK2erxbIUeakk547IYj7k6hRNDMJYWkvkOrBguPPTlDU01SCprQULBX0N
vNI/ZADsfNEkEgpn3Aq6I00CFGb6PMPzLmtDR+AKUfFAVS5c8290wnFv7tVzCjmn
m0XlNpN/H5CNEb3IVVpj+ixsnaWuK1+Q//rhXhxShYaj8vlple7seyL+Px1xpGe0
BJxQ9YTwHRPr50GBc0s0R6nbaYvagZRdBro+/QYJZ/8CtXSuJyhKkKfW/sehyeHP
bBCQAYPQXrnzhqBVzv0RiJxosUhQAzY1simIE66O6i0611iGXvUDP6UJ9wu6parp
ZcJQeyR8d8paUyPLw5zUy+GX9WnIF1ZXw/oeRJPh/38yV3KzgqppKMGmIdz8OTnJ
q9JB9QGQ0sKbs541rhj+6Dqqd083X1+fRnkEQt10nV+tpdS1sc60sCdxemfebSYp
PGReB3Jot/BV/QSg79aRWLdMVd4h49V9dLxnndh4lVCvQYx1KitOgNWrjXRu6dPU
5M37MzfeW4t4n8NUk+yKCWlchoZNMhEz38vdjBIcnBZTsmSqdQcP5Kd7vUsec4F+
/48leIykz+Y3mXLI74FnJsgO96WWJBjJHRoxc8WiW9hFMICdjgOy1plcQU44oxbC
WJMlZZNzPemrQMJot5wOsaVU4R7+MUb/lJVjHhQIis4z/BzIp85oISdBIEbQUHMW
bbTIOX+BkPu9JX8s3aP+HDs5SBvT0vs+j3HWQme37sXhk8MFh3Jk13h5y8ON11D6
eULUqa33e38ZXjb7OcdaFYIpMeB2+QDZ7gD1FAPD6oGxZUZOyaa6ocpuXdgbH903
kNqh/aSBxzQwSIbLPB9/MhZXrlnHZXXOKTZrbxFv+HWgz2Tjf6YwMCGB76xKOSLa
Mnv/Pbau5zkMy4Sl6D8LvrDDEiY5zaq//KIhnGJFvuYAZfCTIPo2nrXvi6e1xYcT
i/H57Hw+YjDYx+248AmhlIMnoNnpq00tf3zJ3b71l+gOHCqxbG8JtUuot4n+aZFi
ZEucG/C6YKNLRUBTKdQ+ibVjiUMf4S2NOlYnX5NnTHzXs0o4OrNl+X0g060ach/v
cGTMpCkDzcRbChb7ywyKT3T0ywFMGqN2XRyYkblhTmmLZdnZZlGTdYQeKwejP8cW
8CrRDJZRh/vO9g3VimEkAbun/chgjlgHZ7SI7dFgFJB6Gzl3IBGV8gATxRLep0Li
bXYKhRvsZH4GJbkM+gHvjAE6MynPFgBjd1RCvaNpD9HXyWRRDFCAkgjfHh/PidND
IGU2HFdCkKcdk/USBleeSRlBV9zEDTL6b19TnMPPony6+tDUibj4NKYi4hMJTQm7
TSmSNbGXH3w2kdCMo7mfTNT04rOXoQ5HwjAOT2uQp3LEhdgxSMycTndLtjyg9s3I
qY6gNcSWW/p4xFebStbDY5WXfa10SEjhzb6Sh28ebvCnex6owjBPzWSBeJ4bapzq
6HEZdDXOyqXzqMZUb50FUXCMMPw5fTAbXUcTiRjIaH2n5wWoy8ecoOSkGVZiXDTE
YDIrKYL3+x+QoJ9l8IUFdJ4kUK10ntVoZuoaBKdffdlAQGUxpziDHPO0R24pfgpF
HPxCjzHepotAsIo/RyFwdduGzsvPBnDfo0OGVmVD0/h3zHeJqoIIVtytMTYKMdId
KZYt4gbtbJUsbYWaHq22bft8dqxpaliwv9T7Veo9o/rJh9KkZ4bUnBlS7EjB1O0K
C0rtrI8ZHY/ACvDtwbNRiJZKC2hCADr9fWW1Kryx+pX0jfzfmrYWkUbGqEr7EACL
lB1XTvfg7iZynP1U0JW7AFPrKFRPR6uGRItCx4wPe3SBcYm36NvQw5KFnAuMtLg4
/BlMYR/IY0hZRbAIHzVTgDAaNNR5WCo3kG5VNWyP6XFqrWKpCBZpENxtOFwLUfSA
YAdmEnAwIGUKD8ZN+TgrbDdkfVlnupPVhpM2u0/SqU1qUrnV4qZ7pfRuNIBet+2k
8SWplTlG5z0HyfCI5u++93VatVfisM5Ep5j6SN5l5x4H1UFH/9pSTXEyDeF5Z6Bh
U5pyhwoy0Gd2gbLL5xc0SzvYgJHOgJaBJKKhfsnUurVL7niiUWJ8Kp/MlyedR3bO
p+nX4rgxYqBVg8Hin4JPDqAa9sCYh+TyAWX68CwOMzYXmRAM2HC2gHozM4eOvbkM
2XUhwVSX5X3hbb50vVnozfsGVX1b5BZyA0G6NHWz9Si8owni5p4Cbc+t3aNjvhAe
IV/8uDv92lEiSfUDKC7ngcDw0Ip6BLGYEMVUAyxxtzUCNjh3Z1pGZh2X5VrzjZhb
lBx3WUwZebEZfjDT+61nfYlXwLH68W8PpFK1DKBRIRNP7pkdgDoZsH1STMfemyTJ
fVKm1cF5/+IIsPnrh+i9bdV4u+EQUpQmEctkUv3wRlLkY2QxkqnWLBwE1EmJm0Y5
a+MwV2UnEaff3l9qAlXjyxFCxSJaSGqRqaf1hqShOxUxLibSOwDrlPhaDIarvUHh
JtrVGuGRhrHG9hldL+DF3nuXq7eO7qxdjPXXdmi3TSYFHhdUjAulOq7PrQg4XoGo
/vAO460wO3N0rNgw7cTilnkZeAxpC3E3KXtpIs0q2ZvoHlkLxhVGKnhsrq9a6WPN
uoaU+gGH70a1a7w3Jl63jcnmsWeRihPsFUwMquGkpX4mn2YJIcJCQXW4Gt3YC4g+
0p7yoir6clLwyD4erE8hv1gQHsCZ5i22Q5I+4kkXa0wHX8L2udd6tEbyy/9JWmSd
APNiL/2XKaI9gzNDqdnHh3x+wRTlcHuLgAI+0rlVzt7Uj/jCpBErQ6YNuDQQs+2W
HBato4SNkm633zApS360XuBixlbYQzZF2t4a5hzXOyX58gA6wG86DQXZqZXshbl8
2kxGZwK1zBsxzTe570f/lDij/FQCOj1i4DHHrZ5cPa4AKdxIkWoCAk5EeZi+JiFz
>>>>>>> main
`protect end_protected