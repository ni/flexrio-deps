`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
JqcB4Dlx24+2+JyzNOorx76iVrkJHr0zy87DhpJ1f4HJNhyIS05Ec92+FFDEBUov
3sFpGjvoBfdIhgvn7jdPyU2PpCv4fIThgVXg0+/pmt8MciJkEeHEFiF4ZklmCHyK
a3OslTX5Vfxo9ZU4rTo56I8eOrYC4Y4+lO9/aoZlS+CSKMJPV6Ce0WwR8Da1+kSh
IfA212+8/3EIvI4EiBKYfkDGd3OheRvVcuzkCylX/afcbKw0YFq3N2fvB8iPE5sq
/iLMlYu4soasJ9xgCQfmxbRbPIZ2MaGDMg4m5UE7UOZQrcRwDh5zH9ekYvpEyG78
zhy7q9ruoZ+cfBMljkDfZ5Ho/GIu7xvlR1pKrvBXNVaC6SPzLhuyZTlDarlH6PPH
zRn/UqIvorJzKtXPdOvajD79/QJf4DaI4nvguWM5BX5o5IkmaqgqFfwQWBSNLD+K
QloSKkINggxFvnMG87hmU9+mPEyw06qmGRpswpruOT/u80K4gU/AjaLUe2ZfJGJN
iIY+KyIc1MgM38gajXYoKYKOtJ4N7BocNBcRZOIRcMXkcz5iaIBnC4f3oe6VwYdj
UY3ZCMIKW/xSMUbUBtAc35I9nLKDAnTEVa7OM9GEJoJjZCwDEF3Vsq7cGBGz5fM3
GQCrRAIPZxcpKiDUODYFmDthEFmzZKvnSS2RgU4t8LGNoSiSHTWnEAi3Vx+DMyYQ
8ojvsN/sHvbg2BePyUBFBS6y8jWbVl793//kIcp1kp7Lms9/1Woq8u3c+IfTD+3g
ANokmrYKFxl3b7/67e8hg1ukdOaED44Imx7qzxtbetX0wKa6hS1eRZO+JOVrWOJo
TC2zmlgbYqNdBK0mA/IoyfbPsX6F/tu3xXTl5O5Up1OOwgORZdpZdRlPmroKulUO
0rh9tU1wg21HSCvH58rl9uNUyUDZ+mEMKSqcoRs0/3oiivwvyY2T3SCqrCAPXsnO
UIzg+SqSbMImscTPDJQ8rsxE1C3Q3kFpMwtlQuH/OJFlEVJ2tDNcax5SkLvy2MQX
mH5nA87BkB/TVlWMIfcdVX+wgXUTu+5vWMg8X0p4POY0hrvQZHvt3JW6IxQ0zTs5
eB85MZDa1P6yKT4kIOOHHIh5dOQWhAFVqszk3JMhIUurieIuUjwQbmheI4w0hmSV
KmCJcXEtwUxBhLfRsDZsGuA1mjnbGu4UX17L6/3CS3feIBle0GwWU/fHMXjS69Hp
OYCe38bX/xRbDmnC4FqVoQEvrPWSH+2z8GAdJDCXaaotx/4KyuCQK/wxlPxSnnJx
6ocTLTbxddvnir+ASGhfjcopfS4eWAAf38+hsDfENUi0qUFuhyRB5aeWGe2mJbsE
Dwnhq0VkTOPT9VE4BpccLQOBqErE/+z6PNkfBeh9qCHVrLXowHXVYtkMv0cOTWrF
77BTcKVWG+Nwt9htgQH/EZqVuWN3S8kutLY9cKAOPrT8bqUbp+ExWWLKzotXDlwl
T9ZAc14Zy48AbsSNZ7jSv5HPykKdCI8bh6mpptIlDsHf+H5TeuhDAmNmJd+gvVvr
kFUNtwV3SvUhpoOTZ7WttbzLqzMCJ3NsLGcaMsQ8gQosQ9FnuDnq++xn79qdlU+S
NSEDMI3GiEPNKzEJZG7V8wyLn4jcpetzQ4tSaoFVH5T8AxRyRvF+AcIEjZ8+e6gA
UcPKUqnICKYdwqpRd+UBEaMA/rd7mUF1wGuOfnt+VkhMSpJJHVgv/KWsRryxqRhm
Ij2jhOqVmjuqOSBUyBf2b/0mad7hkOaZ++0RPltlxg0I3AifjFpb+v4zJ4UarNcH
VRj5A6S9+BjscB9ohidAY/XBLazKnQ4t9CTMMvdpzw+/mxxVBdJVuFN+ykqPfGdt
v7lAkQi0N2EwWe96G3zLJJo+oN5KbgaM3mDtYEUaye4Ishu2RzqsSiKwMiU+gy8d
JcNg6scls710v1ymRgtPDD0gx6WKnlyEGScbO2DGwf1nEI8j2n8RqpdsmmX0ZAZg
1dl3G0oxj5dMcBXu3aIgQ9B41NcKWP+U9A6hNkcfEfhz+nS8Sq17+YDqq/i75xhQ
ZsGrpwlppyxxH2l34Shd+jGP8WmS1NFqD8JGpGFU2N5eZQQclvddpB3xpJmCcjrU
dz48ikBX08m+9njngevM09UpMzxobihD3TRzSyw19XDquyjTmYUawifq176+BZ3e
8d5XhLi4ej0IhyoQ0Fy2mVHJhwm/o8U2pPQ95duAU9mgrywitQ5egEeBgCDjla2Z
yNxZ+iYNgz5Ygmgu/t9kUHNOX9uxxHlmCk8iL5pvbtue5ZdoQzuGqqWL2QTqIun2
p5ABkfk1POWcd3bqo6XPwVFX55Y/GbiJbNRQizUP9gLGD1HHVmVLWvbwgrk75Xwc
pkiVcbkIoAPzk9mjuxKMKg4tHTuaoCLX9crk4Y7XHX5LRDHOS7XmHbtQ/h/IXJ3z
q1e87o74Jz1+iug3xvUxafRjoIR1YYab0sHx1z/YS0GD0NylQvaiDDY2x1KuK94o
kFdVC3s+U2frVG6NZcbBPXzCAGno8MfNOudLjOyXbIpfLFfofALFDQE7/0w1X7d6
2izwXPnAoOCaDpfNWSCS+HWYKMRWt3Vifg7ndtlpWvopFJx8NH+KOUJb4EJjXFI9
txHbVP6tOksYFp8OXeCs8kTAAnTb8mJmTaK376SsgBzYrVH512ycAbLa2xVmLapb
mWpowaNkyJpVy7oil/fz0w==
`protect end_protected