`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcB1qG1wsgtH1+m0gFKduqxYyKcCI9Dc05PsGZ4k87GOe
EF02LZm3cL64OQ//iyluItFHbUOmKzt9FNDX113dH6uT5cE7tGLmpYQ6r/mIkVDb
qBDzs1HwsY8KanYce798RF2R//8UfVrCXP43x1NEVwkk7rgBssc0WNfCk9pAmQN8
IAl/L9FgcxA07GRrrwtJj6zeGxMgMR+n44AeR41UC9K59yjHo0bx7fCuhsayPYSl
TUhhW0zR+SMDi3FoCLA7PDacEX34Ga77eBS4Lh29beeVVF3PdKgqTqCabSDkGmn7
kstjLl4WAREo6glYm/S6SG4FbedlLAw0dvML1YhTUH+9HVGGn1fo3/6D6aPYM0Qx
dVPHM9SHHbOxQnqvrLIwlUIVcijeRiqY0CwBm0ZgVu72fMRhzdkadiiXqWhkquDb
P5KNEE4XejYCWmc0YfXhrfUyzPHY/bV/q4wH+vVPn5gWRcWti5H9FPpjCLKPa+4o
ZZNt03/C2LXxQfl7dLD4L06G53wHZEMyf4jC94kGPzaWTx8KFxP3mKKKwGxTtJ15
k5GpwgEwN0jLRT0ChzL9IGj0B01+pixUIX1Ukr/HN424CD7akBIKaZ74PmtvG6Xb
/XLzwcrBkOBUHe+30RmxhcyhHzfRqZh2yKlgmJtb9t4743xmD9oa1dRWTOpKCYCj
DTIzq7/+M6dWqq5TVITUmgE8DZzAcXDgN/lTnVpg2dBSalk5sbLBHB95LrjTCxKn
cxBpfO4QmzrikXDb0ivnn38L+y6zBdLbsvD01exZGvBbC7XmjcXdW2P8AoNbTEd7
0g7KmnVm7R2soxJfQtxdbUoUEh8rxWt56uqi99M5E0UIkl6JkUmyCOEnVZBrMBfY
nyclBKFkAmeTS/TzJN1ydacs4w5KTThHQI5sM8T0wUm/KllgugqzOVOeYHIaacmN
ixjJAznKSny51+Of2Mjk44RVPnx+caAri7wPXj2AwXrhQDY8bWFrwt814Jo7yQcC
espNN3cxFPTFiXWFQi+PIyD0IbcSsxRVav37wHP1KKbDyr60AiUQJlY4GNhTSyH3
A/9ZA2Evi7/H4UTBq3Le1FqshLUuo7p8SOwiQLmOJORqB9FiVPgJz+HiOEEk0uyR
jP/cTR4/d4doyJZdJ63AW7rEUDv9TaPy7bp0hN1mzgGuYsXB8TVM3+9TBiHtoChV
cOWkWNVfaSMzPInqyBIp/BxojisCAEHWfJLM/0vv8WKqhq32mpL3fa3o4wWBk/x6
P/bB7dROwqPKOgXdJFgshGoWeajt0JNlpj3Wexek0pFT9rAcN3CJgwIzioxqn/OA
GCMOB33xZkmoO38YstVrr0sjNYhAqTex6kEmztbhjmYDEAaSX7ctgrs5BqKyilH3
XjNCr2OByJNahVUI3ebqB6ny+O3XIMQLj/dq/2Wf30wfCh4TZC9XeAb3pMy5EKAx
X5Q8DyD6dov2hYQ9hpEpbP9TyY1o+tWZG6hC+CTQd5XXy0qhAL2hSZQZf6g3F0h8
kqzTtrCy4nJvGimhyM4J1ET90LidhNcObTerBWAkD178CQCV0Lf10XxPQUNo+/hm
YoRvAgvpMH/WkNGV5PBCC0fO1ovBT4VybMWymKrouYD5kXM7czS34Q2vn+yMQpbj
g1drdstR/rFNqlNH6O4meQh2n4JTj70ruefupoA/AcDf0XzeQpQVZR5fJZj1zWa9
kLz/jk2QEIUl0ghIaVqhmJguRWbZAK8rk97B7vIGoD2Q19K2AyvJgxOFzij6k4Ps
JM6fdSCjE2hQzAkxmYA7V9fyYXdc6L6MWGF4EB0y0TaCuWIRalMQnNVhdSLJX/ak
nJOXel3KokDZajMUNJ5uFKIAE/Tnjm/VjwvQi4gtnpgeKSeKOd2rCQAGLzkye54H
DKP5Y60+1HmU9UxFaaJF7OtQ3zvMO8mCPiAIEv+o81KfRiajNEx5o8HStAJ7Jte8
YfwMGiwb+EMn96JRYftel3MVs0uNiJGIRYcaZ1Kkx+dWypj/hZLVvjbu75HCjLuS
dRHYABK4UnrcnJLCpVx9RfxTeh/3SguUWIHAx7dvoc0mOdnsUzmuNWpDHDD/8O5c
uEHSVlsumadh1YsWz77yPnxpCl6U2UTOZjy0XLQ4/0fRtebUBEuQAQfFfQGVqFZb
qDtv+nZXb5+9chwXBmqR1fB7i34dAHX9W+VLYnirFIiZx3onmL7eSL7YF1VZVf5S
aESvzfwX2HxcRW72gfiZJDvNN9kKAcu7DpffKgHRlA/zDFgBPRQ7gkkGhrncgH7n
pwhmt4GlLJYPFTLMa/QW6w99nqwKprf37A1kMK/FEXGG1a8tyV2AAOQ66aeOnVA3
ohFnDX6yna59s+Tl/g/DEEb/i8td2Io4ZecQybBhF/nxg6aTYC8+6qdH1/w3OQYq
q5g9r5p/n/rSwY3WOM9J8gtWUnQddTumZi44nPMYASSDonaO1JywZKDEOn6rvuay
D6wsYdey1EmffutZq1fmqgfJ8gZx7YCuHaLNdhftFjIt3eIpvZTw8OED4WqbsdM/
M+3sKmdkCbBan6jSuez/UkCaXud4cnd5aCHeulYBtXdeEPteBlZcHUhIcVJkq/tz
UXerrxDhAIy8kvciouJJy3OVPKQ4yEz9E7bfb5W6QBCxVVJLskzSXemMFHoaF7Bz
3kISOmedoRT+IuF8n8q1m2b5mDXYGR/ne5zJdS9rTYC6nYho+/9URyeEU6kly5dV
GX7tD4gGnNEtMMvvP1lX3ATZ9CRsw5cBKqJSsRUyvua176SNnD6lQadSh8fEr/na
8Woy3BixzvCSBauSs5boGgoPGSoRtZbdQeqB90w2piR8plNaFmDxJtiWGVm/4yut
DEL/gvG2tJhmZuwyEFkzh4RuZexJgvYOehzpTnreF/UP+Kosl6g5z1GAp8OhbZlJ
e6EJ20Odh+4IsdtH7v2rhp/X/Bb/y/ktGq8dNc/pq8fUaFHxPL14U0PtWHtD9cI5
sfcckRJr7XiaOG9IAVSHVEVexfK62YV9w/xxGwhvlkK20AQp7i1rI7xILnSmqzzU
dMCtRkUAdY4D427oxQkdRo8galsh4Kc51nXv6/JyIUO6077/Q0m4wVapdn1FyXoq
nE478v8KXy4Te63neB2ryPiuSM/n0NZRPPBcNXHrbp5NBc2y/NXuCGBebV+NFlDo
AqogCGFku0C5yFK0pquwlnDJHKKZ2P3Xuw4op/8PKMiPXJdnNVoIvSC9/GLxFswx
D8QByDI/XEMkFKcoQGHE3xB5rT5gDxdYzS03L7n1mrmZ4439dZzjK9xGKEMrVt3+
U98luQTC6Q/Qcl/Q+MD3dh7IMfi8zeaV7q1lzOCqB9uCuzFhKXW9RMnI/rPnqF2Y
lcHvG6m3IlyrxJj3JS8ibzFzWCGqtRQ/c2NCY6v/TOae2BAcbLn4zZEjog/aIVqY
4vhOPEIsbGkS3cKODgmMYJvlSxIoq8ZHMu+HmEPO07NJ+72Z7QBG/+X44ZdoO5te
/qwlttQ1qROIFi+cGnx9JlpMj76rH4B2CVmeno6RNrfEOGxJUrxdbp/Gt1gMLv4B
fhKGxd3wrg38L5svJBntRCoRl2AwjQ7+Vyt6FSIUcvJk1LJWHFxcS6dBZq370nzK
UrWo8hsE36z+6qRAuxsMRVfb0IvSSFzNmsfwHeDJCrOGLQ83y2E1Rusxii0onwZt
N9BEqiQlTEKWtN2Ks12QvNXrKObPbuesF/sLqwznRhUbeo8zUGftKe00mrLpBUf7
XlWO87tVrUbzQxH35fUJU6J5mc33uLE+lAwbWpxg+iD9OXOsgYJNfkq6db6zs2jc
uRCtED1kNsyKbNA0EG14CuB/k/Oyo4mXf+TzDAoTHnAAxan581E+/Nnjy2ifzgFz
pmLJEa4ElUqk/72yronLB3j7KMBzRKUIWVT+KMDnOuJaHw+wfFDsLwQ0gCsrfU6l
2Lyz8hF+n/4NQc8AsrO34kPJwaOCPrRFSnz7GfK+yUXge+xfWJ2IH+LIq98oUwc0
62TY087eqJAH9e4ebZspDbBTvTAKiCMH1Y6Ek1rdRUxwseALBnO/IcU2483u4zYu
tQU+Tr+PyA1UQ78hB+l1KUYdMSqXJm6svjvc9NjmUbzwxwHqmGwza4TKhAn4dPUs
GixdMkndaI8h6bxdvbihUJ2v6a428zInq+Cz2AbTvRrLgBF9ogfmYh5t63+ZaBI0
CcwzghWZON9FkwL05PiiWf/1YkPGyxwFEJSJy+6iqh0W5LBoJDWmarvuUwdeTllQ
Aqi7KICF1r1xvN8rC7OlwF4+LcSWjL9bfxrnuWRBvwv5WTwR6UbnxwmfwVrI9PSD
ow2ay0PBwP4O1w5XOpDmBhE0RX1KC5k7rfYHP7j1MOyTZ5eEwk2QjkpjUXn4KfQt
nR7Fgdg5YkP9+N7TESI+BFPd0p6Qh+bAmRlN0EWR4Zo2OGYZY+Kt9RXeAW/gj2lk
weejBBdWtrG18v1ngJX+N3wlVqF3Q7jh+1TtzB/2ojqV6q3sAxW6cJ4CzSBqkk2h
/WBqng50qSuxVbrNnnC861+XLJX7aBwyxufFPy2DGdrC8t6EBdizOqUkDWzPA60r
JLTlYQfJueS6wIW4oiBoBrE0ph9rQzfmFsrieoXMvk5vmQWszKqAKnme9olaSpJC
kdmtkm873TKNUaJCfJJ8WAPEPyNIoJIHzIBYAjI3QEgvopVmaJzWlzlCKsn1T3EW
Xi2z67l2S/sxPjckaSk4xxbKxCgX+v2mlhs0aV9jozzV+hzYz6vdORqsFTe1irW6
XyFFTAD3HiqnKj6RA9ob1ur8q5K4JDlXY3wUjgI5GIsVeafyagkj0R7Rc8l0dj+M
Mi2s7QQmHELyPcNs/mo+2uiMt/rQN21BNOsC0YEvBqz0EZZCUHEsEoy/jtJck2fx
x7D7kUIKfAZEdw3+7CPchHBfgPXR3jtLkTWDt3Sn44phzbaVpbV7/clMZteysXnM
ferIJs+wtpqER6tkfd2f7EajtudILSQpCHalSeZwBgfFOd2tuPaxYbM+ilTTGKnc
2qPcWNM3xeeWcqiKFyoy773XvddzAleyXNXAfjQ9IN6HMCt6804V7myR9r6FCwN3
ea3O9SA+qV/SDGwofDeSV/Elm8+vZGa86zaO6tr6aVD+q+7OZZFMmTvAm9YpHSkd
z+jLX7RP84jc8qD/sjjdXVYvT6p7XvOQAlq9KiI/bU2aUK45gfhPsRBnP4KaHd3E
qWGj1uFvQ+AIjQK6D4z/AdwFXnPoAtqSZarzB0Gf673jAMhS0AdBVV4mcui+NGi1
7UZFG2oRfH1ZG/uNaiiKd+S5xmuaKe1f457zgtk35koNLuo+MBEh2amtXHogbmlK
gQVvUCej1/HEJCfCQ6FQAx+uyl1unH9Ul4aivru8X0lcrz/xOQU0jkWRgXSMdrWe
YTJceJBdWjCjnZD4YsHPEfK2F7L9eYf1Ep+nsagRS7BDmPrh86BH21K/hedmHaBF
Npi3pybBxXP3ZbSqn4S8D91o4OWMtELfa+y/f43Ri3RB4B5CB+EIPzfiCU4i5riA
ToCCtwE/+QwpfE25p4aSkSafVERCyMEVzf43e3fau4fnxcmVo4Y8qyV7H2KefW3x
mb/P4OuHFokHvnaPYnXyfVmQimi5JF+zu5dSCzjx/iec+iLw0nHK04h8znCbB86X
YGeYddzJDnuTD/IHAk/xTG4r241qYIes+nhvXZPX782yAJE1wbdzGbhx2gYsSvJH
dkQKJddVTZMpquc/8+RPp5sj57wT3WqsOXfRpSdpEnKGrVVpTgC3BnCHGe9stzw3
A8Lg80p6LHVZdvsBeCx2shxHpk2VFRxlsdlRs3QsAD7oARZg97z9uPDberYwZAnx
TppROClSFahgap5ckmUhGEmYaWOnE05DWBFYiZlgBy7hYkaQN0sZgSnjP9jCj005
FC2S+x/Pwil8+j0hmhacwN/EbXmFoHolSd/+HtFtk2qNH4b2nml/s7Yh6MNRBy75
snT1PYBu3xjWczN2kmlhMu/J3BviPRTsCRrF1n3o9bJlgiypUlL5u2NNz3FbnUof
vI2KZG5AbpM7Cyi/KEZ9/f+XsxtsXL4haXNGWmp8NQ++/FeAVyWr/O2brwpbBMEX
fA4w60+DqGrOk/xFW7FAv9xpo4+qGaFriQZPkLOuiJ4reZoqFrbafkgNh8Bsf2Wb
AL9lllyy4bxEC2nu4LZrewBbaYqTnzY1e/bWCSNFquYTe6TXxZw+NiR8lmh1rCjq
CYeymilNzFq3v8DcHW1t8fKqe/KnWcP28lnx7sNwln0hUh8CyYmEn1YhqQKQpAlZ
H2ewLRd5mL85RLProiHuZJqXGdvJZDCjbtvXW4f2L/3YuSmekblWQEyhWZZuXik1
kCPFNiHu04hEzLDNw2iQexe4CrMdTfhNPcqKQI75+H8NskFjoDN6pXlDUM3X3ZMb
56qAK6RpxDTZ6e3QGJwCYJa4zhenefKmDo9/aPZhH5a5Oj4RbCFHpeohlQV64YoE
wNdponDbjkx++78k0/5UaHq5rTlcAP+H+U3//uADTVij3P/AD2sF4DCza5/oAo3r
qJMY/I1IGSdioo3JPA+GNK1Y2J3UJxwDMtbJCPuaPEQFzaVF+HOyiiKVXedKX4vN
CSAnwCoQ+c/UolahX4uYjaa+z/xX+CsaK/U7lz9cKLWfOcXfBOD61xVKmTHw5Vet
Fo3sfuA8L/2vclvJOj7iuUsibGMBdeQF3k6bw9TmYDYNTwlmC5iSKye02tsUxiFe
uZ15NW+Z+hI4UXzGKYBn+YXa+o+1O21uAUsZlTRP6Fmw4hee0oXRQinYjuSa3cIc
Dllh2wSVHtsRz05ERJWiEYrJ0RAemD7ApBXjnilY0ApF4htzxtPDmQVgVZLHshGU
d5cOxmWNin9s4AhSFxE8v/5GOAHK/L+uwPiiUjUH7Dcil/WnoZUskgH5rU9D4/vc
zmZqHURRW9FvPdNjGVI5Ytbs6SB64slbjvbsNa6hpIT6eqwvnheT5nP94HSr4OpW
7DslLyZBx95AASdSqjnOJsnJ9K/7hw04OxfrVkRAZFnDg4F5u6H9F9vSz526b+oe
Emfc6XK15BFlc0oGDbITnM53hUAl2eBEIU5yj8LlLYZhfQgz1pRkc8bUWAasQhRL
F/72lmfGoFrusMwk6u8JQpVbaxzk+ruQL07ER4tdYBDsCe1yfkrXtbnAAoBx4B89
l1mWVr54pt3vkg3Yophp7kRtMI9vN7r4BoXPPg84MJyJNot0vrESiWB1U7xvbb1a
EXH2TQLu9LJHZVlZg445DLh7MLswggU2niyGCNsk2iUhj9wPXYVzv0WcoT6xoRHv
5j1OGHVEGMqu/CVMpQTFwbQWq5bCen3w5UqBz47h9I7ljXZwYuWXxZYpkSUWOa8C
oVtTrwvq4D9XH7/ItBz35xsnJrfFqooIHY7LBh1GjSf3Wn+bW3oT2QHHTO9aAs00
AEuRd71iMv96vng7WS2iMQTWJLVa3gfnka9jYWBcXiagNDVaeVE+SszS8kNw4uw4
Pr/6lD0POq68quytvf2vPbs7nLuIypasEJ7lQi8hfiqjXPAsP9/02zQ4oy3ApM5E
2ZO48DAOf0SZaM5ZwtDCixNCgP1k+HixPFUbfoBi1AVZDLp+dUnSRfL25A6ZlgsQ
4vYOeflHUy4pDF614Y5zW5cbrbAehlYZB6G2lT3hw/YoeRvR4coDvJMc9mlrORuZ
CQ9uJThC+2Qdibe9x3gzTrc3crk6gEZWfUL0ygq0q2xl0cBPTCXmhM/n7BqpqMvh
WrVgAfa/9hlwWdQzUzObbzOSm9cjqRyNCSwi3EzbFDlZdFkCPE03AJSQ/Md0wneA
IQDB8Rh0fZOqVg6hX9O/3PBzWb5B3VFrJ/E0QXx9y1ph/IXc9wgxLnRgbGwNg8X4
PJu5tdh9bgrDVSyLzyi6IPFaudH+nClG+Gh47q5AhjsM4sUzgzxao2a2HpesewrL
hKFpQnt9vrIyfMxDvoTm4l3k2BiI+HUhkxjjVXfJBfiQ9BZ/T0xaYi0VIqXqzxZ/
dAdZPMw0W/F4jAeitNYeYpvZGBYjRQXQYomELIgOOlWHMg/gENVl1/bqmmn1BLD5
hH7//J+pvHKZv+7yqk5VzbvGacQ6OYIxBiJjP/Sb9ZhdrI6Sk/49xxWjIvrBBBkc
G5n2G3sKNUMdUdTOGOQSxm9sp1OhGVDFIyYvrMAN8Q2OTaVeT77YIx/29EuqzXM8
tRNaKUuccfhMEMg7UWecKLi/Fn4dgwydZmdZh9HTUHznRePbTxCHor6Wz3PG07Op
hN6DbzCbidHhbv0gOEjkM0seNxLIXMc3v9URGVxzQR1WlfMYQ31h0w3+JES8w2R+
t0ddtHNUP1iG0AORbwR/lTB4VmARYk9qmoec9sOXD8IKOJ7R9qi2FmwE/soX8BZ7
kn+mDWWlTXyjV8POc5VX4QCXuOcUL0Sf/PpK9h0jPLAuovGdqzszP4WevB34iwa9
VINgV8BkvSIStYW0LZUVKpLw/VVSbBZ0baXJbqv9Owd99hXSEBoUGhM2gwIi2Pg1
v4oiyUPy9X8uWoYfMUB0kminfCqffkdN77Y+P0HXdk9+u+yrvJR9UTGbn4NGx3o6
9mrfMFOvr0p2SZNqIGoUsu/AHkE3eUczajYMR9MpYNKHYQol+wmtJb1nAtBWeCiW
bnmxRwmwjxfU185Vu4/M+vU6YS2/nf+4Shv9SFYCEy1YniIbOlZA/AnwxJaz6G1a
FsWBvpa02h+KyCf04dEZhNEDuzFEQqWz8/xrTvYzEkGD0U3oF0O2xYEbja+JSHkj
8600NGrO907aGwdaQ7VXxmudxsXncdRPhVqb9MJa45Ra9wI3mvlevAY3TtRu3czf
EKQxJa8lsim6MXUCjVdJMWwk3eIq3l2ariGibf2jFMMXjjqBRpnxp5q4IVW6ZuNS
ZeJJJqc6+RsTM6dFTX8AC6OjNTxQHie3Up1/Dor8Hx/QPDgceW8PEhuPh883mh84
86MWKCaAXX31SV+6leb51p3YV9/0v1PwH9p2uQoFv6qVlC3YpRdjhiFOFjvByt8q
kx494OaL1gLbr0ImVHfmmDmCEjdD9TxAM/d0OFekowYKrGrljgGYdSx5ZQjc52ha
Kod26GGD4lPRqnDQrBCLFYV/PaSpiMARkcwBDrKQr1pL5fHW+TZTiQhtDHW6t81K
e5K/aIaG62p/FAGgpd6Qy9ZxYYOY3FoVVIAD4Ik4vu7fwe3QUbhFnKxzt+Crj4bp
ZH5o/Q27lwoHuaASYh4rUR79qHLE4+4XGROgf1UN81uNMoSAWnBwfS3vQ8F92S5c
cYsJxclrVcLDimZXbqlcKr0ocPxxbsvEp5UDFfrkdD6B/Ng92irRyOKHvVBMkM+g
cPWTP6hJWm4m0jg4Eon2Nav4NwmGlNVCzddnKkzwKwhQVDAf4reZKVaYcwqfgxj9
7w+06zGrBp8mgPTA9L1OreDU+2qcStB+9mmHTMUjR1lgLF1Uw3uZhqQ1duRigDnK
JSMICg9CqQ+JACWgWhhDoHmwXkQyeA+L7asvFx8sF2jZ6ObxvuVaI++icq9LqjFg
IyhiH1I4NyzxMea5+TPYUZv5UQI7kMj4ri+nWIYzmnGz3g382Ipe2ioepuY3/FX8
gCiCmFgP9o//a2GuGoDvWrePOVF9jSWhG6GZoGczXgDqJT08BrtXzRjO8U03ugAY
/5zKfgGhHMwyTPA5Stu91qB3ls3QN5ZmaLDZadIw+U+HEGkwSDSwEuGtpBvbPa2m
O/60FO+BdXB8GdHCV7FzNpuZfe+LUBUJujcJS9qSe4hPZ0UQfQrG1jLEZ1QYLgAw
cmVWNfCjlWYHQhBiku7YL+Fc4MIDxkInB6VbTTuKnI06/ai55/oHbY+Vaorx4IEo
UD2G/03vf0LNQLy674S+g4+OJ+8cHI68JSUjF3mM/M3Ij0QPZBeUqhtSB2ovL3pL
uyGRq1jT8iBDFvDbhFJXQpqBOvE78fd/NOkzUnXCwXtQDZjvkdHjlMhBqV7I298R
jg0rzfpTARym/sqd2qeEGNr7L2+kRDRCor7OtQQw0zM9xXikxm4YoPkcCK8MjDws
g399bVBSPfQ1rDFv2+ZGNckI316ZY6VjEtRx4hXAvhHDXp7g5GGQeRhnqoRlNLnw
4upoa/sDErBhjFRMJ8BnIk+symJLkwnoskY/jyUsZIE+OqXX+PmD7TAYbSNmvbIW
EpvtkjMRl+nYNIy4PxP7RcGLi2sezMNB/sa6qandxamM/QpstJYJJHcwgbRU7o0u
iPlZxMuuoGIHM8DY7XAYDm+JhJ6VEwZcYArnobFdQ7XmD1U90QGQD5vNilTKfx0V
4jCWpnvSCus/1KTUL/K7v4vNn2dfgV9shfjW1+vk4t1AC/3k13tCehDHy/SoiMZq
EJH/wcwee1SgT+sENHkFhogUikPCDeOj1J7ZBcnVynzh5aXIoPv8PP3XC5i7emkU
1ynUWX3z809JuwHNK8QZof7nsjpTrkibguG/nmxN11AIayH33BriwBZb5eXBWtkv
Ab0I3WgEKIZSkLAkOB/0Ekq3Q4NrLQTSX5I3uzXI56MUQ1kC5Bgx1yhmd2rlKAip
xTnVUf8+RLvE98iMsFCgxgOvHmP9oBSwsObd688Jer1BKoMLGy9YZ+A1JNW1VP6N
oTCrBeReaTBpg9tm368SBgTP12ljMUr+biUFtLRoS3KAU14Xjf3UOdHV7UFT1dxz
ni2lybbRoROfTs1EPutUtnrUXFnN2jBbP9SGH5/YV3HT1WsVUcCzgxT6nyIf0J1c
aPijEYb0c/kCt9vPDaKbh5xsswZt7OBpSPGLbX/huJKxa0IoNc232m8dXpC/mp3X
+qNybtIbpZcqfjowk5sul80mu3WZQYk/lqIfdGgidxyBnN4cwmeHjW9FQc/fSBUK
H5xYWvc2nty4IEjlZ0MDxNDhnkmEJKpfAovBq+8ZyhmeWVSXkwYKkIWVQnivp7aV
bF6iOc+I/uzAWIXcckW47dCJNpe3iUvPAW3VfWx8jxuRh7O4aDiUs7jQrO3lfJ1K
J5HwX9KTfaOzh+eh0OwD92S3v7oq2ZriN8tcpTVxiAZKsq42DiIhXBCzqe1N4y27
UTA+FsNAkAZQ5fX5Jg1H/M80M6n13H/P0ASSTvdaDfY62uUvT+DmMx+7kXo8XGFy
xrdQ2gwC9Pbjuw2175aU5R5weBDSSPoHh0vEfmCmNyawQ9KaCx1Ci7HUP1O2maKi
cNcVNwAFkTelNoipqZ/Bu9uymd3Xw4tYdiQfG8whtVh2SqtwfN6rhx8U81r+VFXC
3XYQhVZy7jvyMSZKyZNQek1PTRw6wgEw5jg0338R92Ih9hd261hrCaCztrH3DTYB
SWHaL/9/B/0CgYbtRprurcmmJChUDcnPU7hM5u3GoNuBSdw0w74z9WABL4FbYMMJ
aSgNZbETnj/bO6nM2SmRBZpZcp9chCRv9LLxuEnEtCI4DJrhJXIS5IRR0N2iw6Ku
L8GlihqUJEJHhs6ypZnn9HxP2JxbENqWklrzbzDBfuzUoj0DxQRpGCAFbLcr0CGc
ez0XDUF5TJL4IBN2EZoB2sjCMlOuWEiE7X+hkgAW+VW1xGrCq1a0da0oayyyjp3G
MOEIWciy9P22m48Ec48izhbQowgzW+IPNuyDd2/PpYZvAF6VQDsWkFzXsuOn6zV0
dMcl569+xJED8QLf/MTLn1sb9CqoYOHLTP9ZPifJZLYLIsBjrxSnx12xVFPKZGgB
XFRpd60dc+2MOa9mhoVdC9bP7xbm/SdPtBSx6zCB540C57JUlHw898K32KUCWa9V
+fUJo+sQKmBXm5U6tuapCqJ/0m5kAQoxWggRhkfi9FWjMotBFwHmwbP7RJHMJRMV
VSDjpcMgUPu8/IlLQE3roY00osjYe71HnFHCCF2KCGB7WIBdNxxdeN6h3UazGMvJ
H9PYnlR66L0IkOzulE6sw1duW2F72hn5Erc4BSpRmvbuUKVK8SwbyqSWCvgoDcNX
gggCUg1E5SvWlpsYbBrDVrILUYOTRvTFlJgevLzes99f2vgXA3V5g5I1vv9YOIIi
8m4FadgSvEhd5vEATxHlLM5YkVLaw67hBD/YcBH8nqcUtCLuQwZdi5fDP4hY/Uwf
B7uSvQ9VUpKDJXDkCHFyTtRLbwBZynZ8ZksdXOhF0ZDpQNBJ88rZ1Sabidx+5ORj
89cL6ktx0fNmCOOMbw1M/EFa0Y/CdwA5XN0C6C6NvZsu83Ycgyym2tzBHlbTKA7h
hHEgNsNfUN8a2Fi9Lw8CPPlf4vZTImr+1WRbBEyZBpyBHVY1CCb5L9f0f2BiZsK3
N3qU15EdCvt5OZnUD9jtPnCITd3Xp2upZawxwE7DN9mLCDUEH0eAMWLiB+5rElTO
dImV9SGEykDh3cNGug1Qa+0UATbQTsKCLA7cJlxSDd6lDb3srybIQFeb789XeQ3o
rW6pMc9xz8+xGrm7jOWOwafe/EMvrL0Oe3GYXuKlMnsZTOMVHEtaerrsIgdI+TPD
oXTvw1sxZshdZQLZAwo1rW1yqTmt8cKLuTonbpi6RiV/omlhzkHPeNw1orjXShpJ
6hL1R6rHYMTbv84tOjzFn/Avk2GcbZPt9Pf0/TUJUKJNMtBGD6W2lOPcOZko9eXg
m+yW+DflmZWIgso6/5U0m2VL5TXJObuzu1eBwgWRvFqRseGBDaNlfSVLgzEELjo1
VRW3iz0GR/wrdKDu3iPmNwD+ysh2vwwTgd1VPvMw3WRKyCo/t+CKBdsUxil9poct
lGLV9rLBv4xvpUVGsL3tFbdrvVvlwpPSs+OpEuEPqmUeOx0uvE6OkmYsCBFjjNim
pF03UmPeSBBKSzRNwhn4xfbd6/2iLGei4+pwarS/5JwMJBYlaCC3F1XuJ9p8EbwG
WEOPBb1VyVdhkqE02y6UxLk9EVqgqt8EtPT7zpviRx9zTcpUhSDSvpX1SzZIpLo7
zVQ0iMgL6QQ5MU+QrhspaqPDvjXg7Sb9qcH3GJDDzIbRdYjCUANNSIx57MsmCaIW
CxouEjJIAhl3DbMg5IUocazQ2foJL9dkhekUA9wxzVY9MBISAoT1EhIAO6GID0uP
34I3W0JZyeo67wLyLb0131UsPC8RShOr6VW3VDU5mOLMJr6/QSr8sonxuGplPsSV
si9yFkwTrNsnOA8sIOjCeRU3/H1Cki22cXcCdFxtsPfw4z5NGmOQjKifGEj9bJNM
vIfoiL8rlZlIc2mK7VkfKAj5KKsuPLV8CAInzdQg1bOguV4ZW7rU8h6xn+GfUcfF
EIQ/TxgURStRHbu+eAt91V+sJ78BZSOVxyOzt13F8NuwoAXds5YdTevPo69+MXhC
PNS9gQ5Q4wQUa7wzRWx8J32IM51qR4ozqu6womKHMHO3xGGGgwpddBVfymxiCZ7M
n3XBI1cpu9ywub/KvSUb3CcuEJMfN85BHdo4t3kpoHhMTG9NFCdKB1wy83W+jAGR
VDeevkHtyTjSsGVqqStrY0svF6nA7Mvo3GnvaToQZ4NtqHjHFf/hxKX03xvvNkga
Vj05Igr31qpItHbUdQSFN3iiN9W3ChwoTopSfds8Jf+NtqI/UJZ2ivWTtx71Cgvj
MRozwpm6Nd7p9qrtVye424U4WIoN6elzbvETA59piEw3MUPvSQiTKnEbvNJbMBSj
i5+KLAmDZ/SUB/axlpqC8DZyejuobs0zQIRCDHW9Fvj2UxcI8gUs7aZf98k7dKrV
NcUP6fBPGpzT82S6d0MY2HdgfWcng1eIkxh5ry6ITNFwRiJKI/2MrK+Bq1XRot7k
LWPtPZyo7XdbN9DLkqgqjsN7N8o68i6TTa3Vl8DPzqF/daAPHqM4T1rQJMZ7N85f
6gXZ2JTKLQS4AEsH/yZXrn371Hxr+F8ND/wZo5XPYkGqvkLGj36AQF0CUqV8k7Xo
BUEGB/RHCdWz0OZP9UOwwVIfryR+Hbf/pdzPpNlmERH51xyRpH0hf3lC+RI/cWzI
Aj4J8VtvFFLV6Qgadx2mdUZIkqCsRXeAA9IwehXtGfsPyZRX+r9821noRiveC8BI
NzgqBeNBM1kpPsMyq6YleJuRDFOCEllro4hzAF1jny5CCKz/XKlPEwFAUodXRprF
4MoHy2nrERNpmZVqe7qWmFlm6yOROeNv5342Ttyzl4OKAzyiraTb8qYhsT+RFYGB
ySbAvbkh01vgOjUKRYKCbSonZhvk+7YIlO03O0BK1pdvTKP6hShxLfIhEXFeiSSP
d0BSUzlK60WWvJ4eJlOUSbHPrMFEvfpDtkPzCnKX+Ng1vhTGMhY9L4R1rM8J4Hed
axUKJo+JbyU6WyFIy7lYOgwFV4i8OgL+gMlYYc9tdzZxToRnJsMktnDLisq+3D2a
xY65f6qVCYvWV9tdKq6MeWhAQw9m66kwEUOhkMCmELU/3CvM14vpLlm+uL534SBq
u3BpJWmI/pHSWHYFS6760L5Fwb5ZVFWx8/N1UG0Yysq5kjgG6OuTQR+wZDnAj0AL
pjMwWG36KB/T8GxFUKdJMAcTsQ0U2ikSOy/w2TApSBqKuegbpdgOH/GPBodDOvXY
WAcRdxjIXWIuVqygDtBGIjIdAP41VA0QM6xpj026W5DdsFFdQleL7ROpRdyY0QwF
RWYzuuCEUbdyoyp3awA/xRtmMRUlfM8kEMHWuyIPM6o/LA05hIstcNA+nWKRiBTq
3kv/aw4/9qcIOBAri1J3pSkYaZqHXacckpLwxMbpvp8kr4Udz9y+akz9IS1jOX0B
JlYXqXp65BjjNl9cY7/OhceFOlvjWdq9+tqtj03VSYiCQoJ+MogSBRjDFIiJH9/r
BernCTRm0HPH6Voo3CVdC6fZi/683RRkdNF6jcRx61KJxG+u/muN7M+5EBqEwR26
XAjs0DycSgJ+dDDhStsA3hPc9a0eG1fHazOo/2QSBOexw/LXnty0n3I65cEPJ2Ld
7HY3MZktZitID3tE2fV0NOnRb/vUabiXA11fmmN671B6qcXmdoEPlZ/0TtA8xyga
rWy35l261LrD0tEWzS6au/2kUpyCK1may03ujXJ3t+g9X4YjH0l2s/J/KabXbpG3
vZzlmdB+/AvEN/VGatEkhn+DtbKhEwWv3AOIpbjKgsSlikNDDM9Rp1zCX2HQbd97
Qa5wdRVDwwbaT09Ifmchvni8+sFjM3O2hLkDNCKlsOCeYvXBjxNgAlR/Rb3218LT
mnLxDL4pr7hLn5f7egv/MEKv4kyngqMwpSmOSvVv9VLXRFCpFcNm27R7kLo0oGF4
CPWEErjHyAu49xQ4ff3a1kAULq9tlMYelZE8ahyzHLrYijiT7euqN33wCaHLFCo2
ZysKvqQ5k/6oIhEGHyf9R9dKeBvjyYPx+NiPBNPk3PVIYezrdeX3eYAhcA++Tj5c
fGahYLJMFipWc8Saml+hARlKR4lfLhpYSmrveOKqw6t2B4KSrxIVIGFcLL1Qyykf
s28eEAEM82teW45QPceTwBLqfrKd+Klh1+mSvO+fu9JQcnsZWZH9WarDT9EwBbWa
3uzv8Awr0BSKdHwD4bYq4YtWRB387FeA5om/JT08vgdf3gq2r6vVWn+Fvz4f3aUJ
wiT501gE9D5c0NjWNG56yEn5NRhlNRJ/uanlUPjZpy71YQo01UHhC1WmftusBmw2
oGxLpUYNjfYPKnUUAp2HjUS6PrOd7urF5ud7pslN7oqeUX+1zjcYYG5xs4yHCjx+
1OBEodQ6UaburSF66pxIHp35uTeooQACqZhJO1xxis80PvoFdvYzlyt/00rGN6OT
Rggy6LXiD/B73i4P/j3NygREgzhHNx2EubL0PVrhYZ6rfvCDxbteLK5uuug+AHSX
qomJPdqMe2QBHWe9G5eJEAPS40I8ZATxRA24eEHjDRqYPKwNscsRLPD2M5PVHPta
VaTzxdHzUPaoG0E1JavOeBZMhRyv9cNX9+mb4hYTiTjrCxS8oe5Kpk4Kk3Vw3Trc
MeBwBhWsCegH2ijzBpAL96pJwsZd450IUeZh52PXsDEQ7Cs9MqwGPIDUQZinZ19D
RooVq71rv5s0+kzNvGcE2HiZGsbXTelOVXvBEOKr7YwnBM82dPFgZjmA42quYq23
nd6icRZ6eeKN0B+wke064rk0OarRb5nzKK/WsvmC7Zl139DQn5aCq7ILrJgY8cuU
/6oA6e6dmRNasvY88dtz4V/l9CB5dTlEyAz4n8+1HvuKuswqri0Yoc36zpkkOXcm
fKsDlWfY3lKK33NVbCnOB7Cx09miB0bDZ6827hApyMRe8whC4mpMgRQ7t4nzhPuF
I4BEPXelB/hydPUsKqLrv85y/tB86w33JTPZxTNS8ZUm7D+kVzZ4GYCGDMkeUoLx
8sVYs9WRaQbPysh8ybMDsgI1nGL6svLDyRL6IkDNHzmyWFKvNkD5HbxpjU8pl1HA
5Ff/QNaZ5sQzaRTpdFGC9b7vnypgDMx8wt/lxm2FSpYebCHHdgik0r742spXCIeu
IO7/QAiB93zpM/4CnuuBhVn+kvWTDgDeN0Y+oi7e3WpPjoYpg1ovUHxqJZjCloOg
18IVdrpWHZoRvGs14OMS8cs8IEcmZvtqBV9hmJEubTfLKxq+zAcXcNxPvAGrYlDt
JIVBZagJ3E6m59gE+zC0Mw7LwaxBx82xBQ6QQIP7HlqBcbuVEBG/UrxsfntbeMkk
YrdWxHugvm4gVhQZQfeqnarg/jzK7DI39POJGadKxc6KdsGvn/1YjRStWidBGc65
A13fdyj7/4rYabGXHLY0T9jJDqWRboanGWH+HmV91Vws6NFGLihhYfLlYVz6wnIs
bXIoWFfMIDeCanZfeiIYyFvJ7K+NcwmUn1PRw15kCGqE9ctbnABk8Tn7MHTsYH+/
/LTvjzw4IlKUBcODEdT30nkHYJdUwNIrjX9YS9kulKLEKboHSPdYJhWWDf3NxIRb
PAf5pYNfz1ByMCB/uWOVTNOYkUSTFeRHqZAm490oXyvW8UnHGzYIc3bIrXRN2SJS
E/PANSyetdToGzZmHr+q9Dzv5C7JgmzsrxZZy6kP7PbeDVTVufch+y2DvMCE2mJ9
HGcFBPbx8WWWZsUpCTlWLNa/+sG+sPJDDXUVdkOvui9nww1AbGL4b5cWNq8/Jz1C
q+a912SRAsLWv0Fe3m4MCC34NaJ5jAL7s5/RpVMWixmOgXP2cyDZSdTp5vjIiY/u
7yq/IDiqSKk9eSmQYpeVHWl1vX9z4lEAH2xbFMmij8qwbwb+WewgMLG/TWyAghFD
VhN+u9eLcqF2DmBqPWhC/5QqCH/Sbjy/5zwo/Jm0KYY9QheosiAD4bP8JmjCAwnL
wW0hOoO/KrOP2DmG0XnYgZZzeIKFLhVAg3VKkba16bAZtY2Wd0ykWa/BHHBBAVZM
D2IY5fN/uEl5pT147pAnKhB8rLCD2nE7mT7ir1a0ybrQzTSCbjEGw3ngnfXZQlf6
1uQAw9K1slJyYhTxh+L639YZngWZdzOizAxTIOyij0ohmAl6z5wSR/IHzs7miRFL
TB+da3VGJX1ZD0a6MIz20WLmOKXN0y+YBP8zcF8xcChCX+Ssv+nz1BnK4hHIpIJp
u2oGJKhpcmnt16YXFNIXTXmuJYdusRUIy2c5F/86hVLhzoYKKiNsn2m9ugQYhG0N
PEzqDKY/xlSzDqCdXGZiPOgETRnlzEKvq5WM6G/KOIB3PlrWFlcsANiqCZAfHcwm
zAFAzF3htEJTZhK39467yyEjNaPWwjAH0LGH2bGwDEHuDE+IwdzZKGWKDEGExXd/
fXSqtetUGW1tFi32nMbPzrzWSOaFfx+hYJMuS1FoNsiBPWr+06E756aiBCFrZHQG
qtNLXnCU97PsSBJbIaGDsengb1iKOnG5OhxLoeptJnCh3mfyI+gdWEUmhxcwnm87
LbhTZpJtd7GuQ0Apl7yo3o1oSsiVxO3jfKb9gwslotriw43aTuZZI1cODZRGZQ94
IhlsDK7C9PGqZRiOqEgKDYK/cV2/wQttjEwEahpCkTtca3NlyB5x4bpTF5JMW2LC
bVI9EQuEfnfKRf+6S2qmQI9coPsqTk3c8SF5eHHDoEWt+tL5zAByHAe0tBkzpzQg
InIXDA4B57PDTNs9hx518Ath67IJT6/2nphuCyrjc2K4Z6wFkeC5/mPFf95vYgkN
7de/QGN1Kifrhttdz23aG3xZ9xLA4uJVHGvKeWm3XUx60vMtT6CjtS/uIcHoe7Cm
6PzPrFZsu2bKQL9Pf/3eYhXi/2UrfKOXEC9wc9mN22HzIFMcdxFblnpt5eYo7ZFg
LWBG87w9GpHhsMXeCGluS2kLj+Cb/kI3pPvnXck2ngXbBQlodoJ9a92esinzqP+4
Va1b3I1sUF2xjVLWf2UUwjHFoR6Egrs7jwvOwEktdf868nH/jjfEe7fddwd+eUL5
25sz4HIdl+9UyNknouOO6jei7Ix1DMdTTHGkAZrXT3KaqtKV3HEMjJ5DVHdFLYEG
kFfg1Kj2Nbvv8UbwRyfNgEJHrlCqrtyEwgpTfLf+FARIkRFxKZ4H7FwXyp3KGWYa
Ne2lro2WyxJlI82gDJuOF6S9e3svpMTu1RtfJUWW7dPzuXhTxtnndj1wGnonDEgs
NyxtSv1JnGVKzY2L6vr6zDqsdv9PPaLpjjn6mo4VgehyoH1riC2sTmenDNkl5BEk
/hKebTW/YpeKEcbiE1mebwTle0ApEAC1v8mnnuxSKv62mD4BdWOG8YoixkasXHom
7Ce0fDGd6MLvO2z304fLeSLMOS22J4wC2JUt85c3MBYL0PEtY5WECgad3LXX3Y8l
XC8tEJjrEuuPwf6ekhWCoz/pShhq0N8e579owJMhV1UGmiClaUwQR+/7ZhIj8/PU
atIsphn5BrYMoGQul3+BH/x8TBmC24Yv0jKrf90bA9l1btkrj3FEqIsoQhwcyP4F
YpKEuCvnBUSnfvC14DpcWKKOMvuP1aTXucMZmLdwe5mCVqajSv7MW80y8Q532V0k
UogvWZ4eTqqKo4MC/vG5A5nbaTCx/tL4FNYArlwVKlTaX+CRRYBK9I+dbheXhiji
Zqd9uQDph3IZhcZ0sqMFUecbtylRNd2BbfZePxTqKBMW78A9eEGx2r8XayNwCI66
X8XHqXXC4lY7WjOnpQ/jD7fUVTOxzKjjeoF7mVEexiZg6aQcEyKmS3JOx0cD0adJ
ez8wroRYTjsc80SZxeeGVuun736se30+7lhifZ6Gapiszu40ZHdftvx0wX04nfWO
lsIXFthFXL2N3djDXY79qlc7LvPy+sNEl26oVTAgsBU4y2nxPth+At2WsLc37gWk
BxZE3z647ltWihOczQsjVhfz/RM/GfxyeKu68c9IYjWNMDBywt7ZXIaV0avrHpu0
s04KpxR5z58Ytvlk8nLNigoYh/hCtXKom3uzP5tsTZTRyiuH3k/9D4Wg5KOpzV3l
TuncxGEfNDPm3xCchnB8JZUOvIJIDOTWM9Dwtb9qEttM7IwW0BaAiKjtitBKyteL
yhIPwceW+Y8BXMsQz8DmbP9ZP7kksNAwC3LdFA0J3g0zDXOTyNnqUjYPAd3YTOql
8wQxmWMoGiwI4s9ftVX/Vvb4csj+wJbC8f+uBLesdOM93qF+azi8Scig0EM6YmYb
KrsThVnZ2XUGMU1RDk3/eEOl/qtzXvUdHPZMCnRWwmmzVM8flo/9heF3BKtTlHlD
V1TG6L7VFEJ8QeZwi3H1jdjAmO+HAQZe0DN7MLVII96Pa+k0NBpubwvpyii1e26Q
HbnCMKFgkSmBZr32TarfBwqDH0kycFFWUR92ceLK2AodbjPpx+hTanXX/3oNvdbn
AKWzibm6vyx+Sm+4eMrGr/5LN+Moo60TXTpdBhXxSRjEm5skZVRbM7Yc3s+zXD7t
tTBGtg3ca7PQ8KVd0HK40ZoAZF1Q3mIQwNOTRqhb/MCYbVptMsvfiaKBB+WLiDj0
cNyoxSOHwTf1S0T6FIFuO8J4uw8nPDZg5e4Y40puTcVUd+MNpz7zJLzBNtixfV5U
leU1umHW6ntlQDKhEkmzJGnQQR1g/xzw7bv0oqkjHL0hD2pIxoN+uQT0PRWnWuvn
3lwaIeFZt+6bvNjW9BGKX1ZmOx0cTRdGAMNr95m4qMipoaUhWJTJEuOMG9lxOyDR
XrKY7PZKV5Xk+KI6B7aiiGmvE6CPb6h8FWAL6gLwJggnrgGv1cBEAjQp/esocCa2
rlr6ItQF9l5n2WFWjLG8CVgd2lpjcBz1MjACO2Ttt3joINiHOoXqjz5uRvWiVqHW
PziZCO6SPzAIxqDb+j+o75W4ZhngHUdOmc8TOAMok5ayxM1gQJW3iktRKV6QJ3SL
saEiygoLaLmdStjCL/1HLVh2HexC/jNL1exb4VymNBvrbAjSbx8BeN/VdzSK9If+
y1/gQtfy1H8G+rzwbTDIgwI1ufbjX7opL6aGWix4f1lpbwA6XZX8yz0/fhxlPpZ8
zuSx+r/IpUF2vJno6oZtnSkvwOqCoj4nf3VSxldmmzB/zop4f8aPUk66zDw4TeWC
znkawkXqgLXokuaQoebhZJq1oc3zyPAD2glRqKBNytIVwDH1/wpVDm8QT3GZ1WF/
yysDl/SDFWAo6O8ydRLQiFupMyuRGJmk8vhviGKJz/m8ivNBB7nOSsSN6S5Ef/Ls
006G0jLV4qQHHgL5yvC7FS8vOCxzkhxZi7VCWbf6AP9aNJRiPa/DtrU4e2zt3I+N
0paSxkQufbtOvsXr7MK3NQh1JgjjtMfq7pf6Kw936WB7xdrjoWL7g3n0T60gC79e
qpXkt2+lUEjgDQit7ngvyfdQU8EIhmbIhbJHDaWEPp4SrYYqec9iN4x5BsEUHnWd
HRC+FmNTKbi6MnUH90px+EeHA4NBFIwg6SWgU4fKK/IofwyFwRKNCOmVEaHXRmDY
d7ua0/HjReJqm1+mHgA0PFwJWxbeE4K3/PUErl0KHpquc2vK3VXf9hdkhIcp7Rca
0rQwfV7NNP7thqB7qqrlfDygQ4fan73VXqLtD0GE1+WDqX7yCgFs1LAFMhVIHhRn
n7p9cH3Mt/ZwpxYZLIYrfozLf2OWCxDxM8Oc7XiTRpMyZKUvbSPJMSelLRz2cb8T
ELbtUwfmTKGn55R/mpf212cC3b964enPfIZfQ3S0ALrUO/w9BqF441DrzKADnFUk
SOwC8jUEnxaTMnBIOOphdXnxFCd2Iu2vvNahUTrA6njXeGsvUE8HSHN9M7Evf2pC
nmwsl57JRJVma/PtIUNrbx6Tu+VxlTdRwUCQkpUHDEs88QEZAO25/ycmbylYIhJ/
slY4xaxpzKHGilJ5zcaBMKRpYGJLejGIG7cBkyBn6R2JbFqxurTcqh5kaGN5QU3e
zVCn/0ECRt75dL1NA39YkC3q571cRyXx4nLcG+c3egZbDZJWJC609YyfMhVYl1/3
ntQvRr+cLvBL67AfEooiz/9OcVQl+Yxs7ni1OvFkvXik5cNyEYZpYX4jmYE5h4Fb
BD/vGETfduBFFl+HXskLmWFu3XZnaDPwKzhHoD7/5K9Z3Ce5ICsQaIhlfja+yaPT
OKnWAf07xPrPaQK6rS6wXIrZM/4QWTsvo8cl3r/25uUXEWjtrWobJ89wl6WwvMpv
StLLVFkf+6jlUbfQXQCWxUqYRzp0q8qFNR+BmKn3dnuZvzVqQQtF9s3aVBBBFe4r
iIFqA51AEQU+yIq3bXqNoKffut/qZLWMl6m/HQkcKFYzTBXSuoYfagFRYq0PNpLi
u9v1VjbAtymBrW6MkHg5RhN4QKEv1765E+wyIJsGcpWnY92EwcgtDoQ+E8fMx9s4
+neBNFzi43NAMj25nFe1SwveCNug6RrCMW9kV6uaB5Vv6EA+6YH5qvDEZV6sPfcE
tCjrT+zHsVveCTWxi50TXCM+CRPff6uOak1T1O0Wp4Ll75ufYc1kuOapn2FPnW9G
n3iYn2u5+BcqKkTQAncazA4JN0PZcaFyhbFXzbc8eKlmeSrC127iB5Au7b3Z5W2/
htH97XErBG1F6m5Hq1EcshagvfH4iTmQEbQlYPtqdf35A6znANPSM1495KGbc92s
ntOBE4Lgd9g5DSiTGI/kg5/drmdi0a4odpsGFm1iLipBiNDyLPlR2ZSST/eyoWNJ
ajeEYjlMN1g/0tTR98jMMstLKUONkvpnWbn5tmLFvuU8ZMXz+E+P/dhw7PLmrKyr
ETbk1a4Gyfug3x5/2hMJnwKuQDJnmWHP1hzRQe0IZzpdFSgAn1Wh36Lu8nk3c/uS
LJhGhsh/EaBDZk3vYkyddM+hD5cGdimWoQ76/Q1B12UVksD6+RidqzzlNjZdhSSb
i/mDEN42EceMnqgVRG30Tovs7sIzhnjE+D04OA4bJ8WRgKbCcP2KwTegIcoPGmO2
VAGZm/RvSObxkEU9esNmxWEbC7QGw9mXXj045pxSm9HGlkRTXBdB/gNcrJ9cBfRZ
sxwugu4EDOIRIFz6bOdwwaZWo0zoNPDtttH1lWnqI0aHZQJ1SXKzWQIGKyy259At
1Hp2GyJQtDqdUxWX8Y/ckDgmwyr5YhZVAK0MxvuHtbQdvLHHanWlwvkTh/GXKJ94
7ZsDGC2goHbIQWy5jeoh6YHGeyD+IynBqS7ko4ycDEHLOwMS0DLutfZrh5LSWcNh
5xe1HIhvpPCNvJYNc18piXfPUCmSxjA8gLBcErJnzuhXJ9fS83umiAiKpACH1AdN
KqBUb6tqizUt29FaVOEhS01nyMnFeDkW7pNi8WEMfyBjUzX5mA5zER4HDdyZdsW4
e8qsJC7rytuLj8IYrCk3GQQDSasUV/gJzP8ZLxZrPLitj053NuumnhgHtlzvD+xq
rW76X1DOdLyFTv3StSWAoG9y06x7feD890fuipFpAz5q1VI/S//SdFmuJyYhaPaE
HDcjY3Ceg96wSkxB46rK56G3DN9ieKyPP7ejTl9q+gmXXwQLf/uDOYDJ1AUbXDUj
GLo4OjZPnELVduO/YQNu3CtwcVtiJIASqB3Ju1W+esaJPT3YZz2pilBky25iTLMH
D+qcsEyDmGJ9WBYdvtidw719uh5aJdEbH0r2r3Gavzauyv4Gy1U5P+7ywspVLmcc
W3nwNzfNzuTvxGTwNSaTTjCGtZAR1RRzkKYr8e0Tf7f45wL3c81RnSXUMst00v9I
WJeuB+rMoNtW+WhCTCWqImzC6561Oy/tmNQoD6U4yQjtwRb90+OTjsxBCNbNRdO9
ZkHOwvQ8dXKt1D8rIsxGRuu1LvQTliTl64VmRiNZDvPFhFjpcpAbT3fjazJJX83m
alEq9JC8/6UKrRDFm4wiaq9byQJkWP7LFvtq01e28YYWfcUgqlj5FIyISaesg8WT
Lz0J/XXlP0/NnqmEbwIzxc27A/NwqHqFtHqptuT92ReJ32OC738my9h4KYZ9RfbL
mPgrHLWzjAU2ilndaCkGcTkuoexvY4Gz755MVUoga9Hx5RTUpaQznID+bC1ak8P5
C4sjw0OifR5RD/9UYim/p7JFGjLGGomHRVpXUtmbEC11LjRx66rDdl+KdODSBdaL
/r6UlXYq5Xca3YHzwXkZuI/rzqE/mn6avKQJQliVGKSkvw0S68ngNzjeDsd5pztk
Mn6yz5BitC9RlBPN0cDoKg7waHnERQW06q1V0KIZUxlkQO6dfj/ouKS+DqMBlBYe
GyflHrSlAduXCbisdx3F+sPcfyP/aIBpACzOMIE0jwoxFJx80vn+rmNv7s22QkRj
95GOI2gtL2wG1RjU2tWM/nhNEwH5wP+AtA4SSs4urLUJavY6sT62t4zfcXUqarD5
PWvFgeM0dOhv3GojXOP4YLlkW24IzkV1qYR7YcaTybeQyWQApFG0Y2cL19rPP2C5
aDQsU9q7WVjEj3yQFbOGkK4eODJMhneaNYhPrlBs5R6U3H+ATZSkvrr59+9QZ4G/
j0n2co4ps5ppufTIOsCXGTl5S4O2vDGX6D+sLfOJi1GZgqg+xIIqi/MzEUWql7U0
cxUER8cHmC8qbHQ0gGsPFfi33Un2uGbqgZbRmN1e+W/zOb3P41p9y0zxX/wLTMnx
XPM3Tx6NRwO3HPBp3iBYj6Tik2qOUdeRlmZ9OcQVr37+JOJzzcRAYM+8c32IBR+r
kCnrUckH1LYPvDBvblvBT8TetlsKw6pk3pw0yZ5o3ZPTMOZghqDOGfGKN6ODkKeo
uzd+pAGPMn/8suebACo+uJaYyneBX86q2pwmczVljd3qqGfjRjq8MjveaanIDhoy
9+rKf3drTUapr2/mNkTLktzkZT0DZ2+cHdtF08yPobrAHn9u0/SXwOpgVlLT9cIn
pg9Ua9LuQ0nbucOIyBTtG4bKiz/pAQ0pMe5W4WQPJ/AEPT9lt2nFydeoCmpvCT3q
pwW5uH972Cr8LaY35zfOveofqxoX582eJRFoDYUhox4ip2FkwnPRyvYSvkjXL0vY
fC2EZBhiJEbQ8ojkJ43KevDHnm1PQC8yomV3OfE3pkxlqd+cBv16TA2uOKmLNlO8
o0WkyKHmNRKBG357v5GAG430FioMgy70tO1vjwUS68ZfXPz8qZm4jkP5rBqRBKMk
zyA1a4AFuyofWcP2fE4XulAEH5p+MvSfa7VglxQTTdMhdvkrtd95r1YDF0hUzqem
ScrMmU8VuA4ldj5s0irAccyYEuHmb/JYMdjAqiWl7jPuCSHXL6GbttePrMe+w/nf
TcArBlPfdsEr8HuRGY06tsuBzCaep2Cb2Mj6RmJGRNDjTfSYvNNzokZACkLX/+hF
CKCrk+AdPvgBsHyvMKjW82RPiUQJxvIeH5eDqVhuoAR6n0N9krOovb2OFG5/dJge
GkVbXXTZ3AQ3JW9KO7jEeZzisldOpxdbG++Cqk+xsA5POQRxWPqfmunwJ1dFskax
DY9J1eL77E6gJyS+Fj6UNqfhh2UMHtQesdh9xs+hfr0iZHJ8hbLEegoq6/mdcg9c
oRIk3y/6gYa/VA9FPCTtaFqJn+dQ5qcZBqcXmOoMn24zb9dLe5KP1RAP/zvc9OTF
l0qp6j17pEKc0vS1UyD1cXll0eLFgwGPwdv3Ag7fjF9bnxf+uJR9APD/JE6kmNrn
kAL5V+iDBA3mjj5lujIp8dvda/ewjVMY+EiU/btK6ntzPB0KWd4sVa5QixNwTUzv
nSe4dGV3xTA+KuV0rx9FIWQ02H5RxIuT+JR0oVr1MXEWd2hnqcxGQ3W8fFS+T78f
YSoKmsDG3+FwGjnH+VyiOm2rRTdSJ7Ia5YGM3W1RrqP7uMUHDjA7z8gEfzDuYTSi
T7OEYPA5WJA6dQ1S7zxkB6Qe6yP9519fPXqzYVqsBQw5imDMT5R9Vp8N2CmqRhU7
Se/axHQmR4w/d7kp3/xKz9BXbs9k88nnrORsZns8xOnemLtVeYWzQki8D+ccoIhO
a+EBL0KaCJNZTCD3W1G+hf96n56Zh+xSUqMZ/mwp0PEt2tFl/Cr2BMv/a+JWwqlm
pkL/FlkT/Zo/ep0kH8r07Ei9gx42NqcD5riC5NineNzZBDcn0guDsLPh2vrbKtVX
d4J0Ifdf/1Gl8dtqRfzhMWyFGFCEe1ztAUnevCzEoHbGhrLHRKS0+wEktHzSgf/2
5JpcmAldOh7CFHGVIdzCwspSO0NIP0rDqoNMFtBCdlBczufm2ScJXZYxMtEQZGvQ
hL/+xhkjPDSJkTLBdVJ5vzn5zHdvRuHKNj+scZCTSMcDmIAgUjwM5mdxkTtDNYXk
pgdUMsN3geggv9Ebeu30REzMJZt33CdYBqGKZSTBH2ne8byvK1ISOJ4y0qmmVIgF
d/SrKZTdouiCHZpFXdgpUBJZFLFN1abb8ARtYpoYVLHeHqhdDbAgb8Mzj34RXScM
OWLBulEnTege+DArloXNtfOMTB4/8dSq8HZiyFWk6x0IwafQVGu22cwT96XoaXcW
54sYARVeJXv4Um+BARNSphy9qVrlB/UuHm+Ow9ESsSKXs1p+BGvVJtKN6DHwK76w
82kjQmrnSbnzSQK4DpIFdrUaeC5mJF94DAnECAFgDXd3CSn7OePyLehuxeHHYiw2
164HpwujorfEFFGFadgLr597j0M4TNNU63jgTH/V54sMqrduENZDmZVhFKq7XxWJ
CQtw5hBUrVpwiqJOwvpAMwYlRFNd6m9VbiJqJKUDqsUiZsuWFy+q1pwmaV3HEGVa
66cmisH+E8fzXab8pB9roMsMUjjeHMcriC0ymRo3PlR1y/pNtVMiDFhaFkuVVvZP
oSQGnrGh6Ft2XQ3gwiGqux4S5wqVCzLBasF1YQ1BKS9RWbjw7d0qrkNxOfiSxoSK
f7ySSDzKQ+X5scpgkRerf53JZAYGsBzS1TBJM5VL+oNbbDwKT5dOsOK7XsGs7Ieu
4GZYD5MTdHX38QzKWG/CvtRJWbuT2oAGmb3PbATUXMIhMg6W7eM67aepGJcHdYsh
gxa8ukT2bUmSBh1ddx/4J8cJoFQ7DBGhPBmKr+NHJuYZzx1mJ0zuYQ5BWGnfTCmX
WFghZUiMo6WcHLKWpJ31dF75JgUJmst+h9qHXZdhgfoE9P+9+BTzATJBUIBpbl57
LdpEh1aQJwpiMpc2ISXyFUBXwFZ0a7qf2rWmmGvN7Y/MiNBcMwyF32GE4IIl5BGW
wE8k1jaNCBsju1Ji5s4i68QxD2VmyWlHsW7aD9gY9jKMsK9/5+SI6Ty4DbH19cOR
WGhnG24lczyi4B/OYIWEeXSmhMHEUYLygknvMCoTBE188NGLMb61NT5IflodI63P
Kiy+8S0o2eKpPLBjMCGcKChqI9+rpwjtleGkjZJYHsAuKYukafqFDTPW4jxNwIuj
ZPzvX/WIpbfxQiiNcKtvuNznGThSEQt/NvPCXxO/Cu3B/n6iXlZkEfnAA45Isv6l
Tfg88xyDQ/Hahd2zZSfbzbotqiX9RAv8MyjlpWiibfibCvlkIiChj+/BR3/5yVJJ
dm0R3qrCTp7aiYuRotJFC3AAQal8vn0jisNEZVeX7IhNw5S/RcHvxbty3Zo4rqZA
VPZv+51mNuE9iGFtTsFEogUQ1vADnvg7g/f9nR+rUgvwHQvI4MjAT81qQzGe9krY
HOve9HI/THlm2YXDZXlZuvcjUq9GQRy7EZBiwPkKvXE1CAK3DUvW32RLfGjnLBAc
B5rkPvixQiTOc5Nx9Gi7iYzknaK0edlnPDyl9go1Ymmfa2PI0qjlIugfsoLaVTD4
huIoWFYBrj30nrdvaDLN0Tsaj5R1R9CwKAgZ/mnQ96rqRerBlFrms6wzlWtKWlGA
z+NzKdlOfiYybvDUceABD/EODKeTJougzaZbiZH+qgorKZRybgXNUDbw73gcr6KH
kwqEkeGvZETxJXq6oyhQjohK/u9feZBWB3/95laz4FJI/W+3/hu31b9GXW/WwPTH
bnXllQhr1PeyjS5PP2U4+kUDusAObMaHiE5qxWSGVylgvMroZpT4Gw4Tj1fEdOu0
7FSfY1KPwJtcnIL6fqKd5VHwkTZ3c81/DydF5Rq2MWgCNbWNsUx+kCemK+0jwyOR
BFHI7hW1lKH8vb2ahunk0WpK+ti+FsKG9rw3r5s/W1YYCSeUFtgamfXe3NxVruKm
PLz1kYBPotavEzg6Zpr8IMCVb9YBRfgSnbxY24ktPMwOdxFNxOniy2z6XFn98xTY
zy+UxUo6HsOliAgY5sWQVi52ezochbUhfv0Uoycqe5uq7W1VIMo26g+v2YJDn3JO
ZhJYyvGU0ydVNLq5zK2dHAvxno+P8xZRvdnN1An9BiRuqiQEBSCB2DCCNOeb1YRA
0zUBplSspoxGJirKhimcCoEdaKtJDAWUVZ1k7HCA3v+xb3lRro4ua5nxlCIMAx/+
ITIHzpOORiWrvUMyKZeXdVrRO/eUgPk+Hi/eyVxBUi9CYahO/xRo41UCywm6LhUV
JvhsfVWuHqP/nWXI/J6EZ/q8anN2fw2LxpQnxzUkhi/bJVOT/7si7l1dFyhPiIME
xxzKcNsyhYFC3VSCYZTXLmc8E+IYPYPXmDk+yZzMlEuBe+IXzPqzCeEjnFzBA/wM
vEyMgCX+XvhBWUAu8bLDY1WHOKOqcfkegeWmeyxUT+ehRI08yTUJIFvsspFydAL/
xR65TDX+YXnQCQKSS6DIVMiJKL9SMQgxPPby7DSjyqbWzQwqLfBY802g40EMCSFg
Z6BCskY4KhKuR2vX4v/91IvNEeFw4WNUSM3tkYu0mPLGnCKZR0uJrwpq2lH3NKMV
RlfmzElLOf5Clae7oBeYOeXItIvRSBFb2fIubdWRSz4p4ECJhZE74JPNmCjImnJw
fxLUpkmfc1lqANoOesvlQFvlyxysfpPwk2lMcihA4PyLJ715yhmm4DaOjyY+VKCh
a7pWya2xvWdBi1NwQjGyGzcmSfySbXfgMiLj2SOtDHNH/xl9g8/bkJR3hJUpyYCC
QW+/kCzMqYP09zfN1J4tzHd8fvk3Vskctvf6JfDw6j+BSPJ8BsF3QERnE0lZCic8
bwXsvT5DysDAiq2UPG9McxYyNXBblZMkc76FXYlYk3aSmV6DiymzbJNM6GbH+Vwg
ysG/GlJVmbOKxYZdz+VK8r/FvgyrMfrDhjOzmD2M80wCckpJkwGzo2YLdfESoWcp
xFMZZpv7+sBrlcGoOdhQjfORC7Of2WI/dr+qeG1oNHi5wKFd/FPxnQqNpyCvhxiC
fMnqKSrzsf/hER02ddtJBxBYnS9ypWSE9aOsFZODhlggqW/voMBXJ9y5FN0tqkOY
TTmZ3a75A5RqBPygjis6uhYQh83o7wYPqSeWOTkkDcfxsyK+xmeLD70sry19nBx0
rwu0WHbFLtUQUe4f3KPkJ3xlqhFY7KEbOIc+FKRhf1OpuykP9KPXFbKRG1Jp5FOD
AmIbNeQNs2akSwL50Z26bGpR6HnGPEDurd4kj8NJ66TOLEIt/1QmwSPi0eRRnFQL
X/7gGatxRw9u3UwbiV5EZ8jzo4w6EENaRJm6FXIidk5yRs9JJuofEkfxLpENxn9J
oxTavPZHLX3f2xp014MLihZnq1nyrodSYqTiiBpsWpIwtANqwUoodB6TRFYk2kGQ
1yTvZhCAv6kJSskPTVoVGsiV99oIDlHAZahpvblj6rkqS6m6KLRBN5UvK/Ky+AtR
U/nbGgsYBu/eDhfZuLO56MJRRC0jxzjHH9V1tR+bOrHP7WYayK/yaROUEEBPN572
sNUT+uP3XUz29hLjaUtOw6AjDOAczBXifWRp2ZdU5NXPKcNFmT71PsCWczl4GdKz
Ldj6PD/ZR7wlkHty93jj8o6dxNTWvrKx2TW0KTd+yejE4APt69KecRx9qEql0O7f
SoowOP0dajYRqxuGZlGO0meOAENXA0uY54E1RQ1Lvcd/DFc6e7/2J4I8dKRuMVmB
UI9CKKQmnddlsynJWbQjhSY9BUSj5wY26cFOtPldVi8c9xkXz2GEvSu04pe89srC
cO8QRqkZjIu4omlLRCDD6soGLAINuuiJoUOEzR2nlbtUa/kkQF8GuUN1KY9tZnNz
Kk8FtrM4nckHPHRjy/kgWw4pq2GYOf45JMg4U0I8dbPaIQTNdO4FkJtVdRuDKhzC
9eLXb/HhLl6zh9ec8IkU0DNRx5hvpTSxVQOYT1M5V1FMt5ecpc6rhRGt9S9jQWJL
ASqI01XA+G/PxN1WBYKx+yKJwXgIrg7nFcFgMLZFn7tLHT7cRC3068cFvcf2g0bE
t5qs2hX5z8sRTIjcfh5Jegg/fjEfTDIfmlkgc3kw1YgXQrpilokHM0TSALdp5wbG
/Gx4n1yRZrFDXzj8QHOUifqABUrRaser18gJhRvYrf0eTK3VGXeeosZo7x509Z3i
BB8v0vc0zbbVCx2ixNOKwSlcMyBciSjFqtYkigEGzRebyMuZh8Lz/2YtGzlPPZB+
kCxFCjPxxOBJPPZZkfqVHdbo00CHfzvMmZWaM638qYxg53DRREYz5UPryaXI8xvt
2gpMENL/wuT184QAy5i1+OiMzBjY352xHYUFPP+9HIMizWyYkwfOyEqkhIYzAvWQ
4LuX464oJzMaQViNiHUoEBq3ee4XmDvpiiF2sJ5WfpO8AuQZMV/vjyjJWQREnpzO
CY8bPQOcWi2VkrTenYBwdWpqhwPpCcAKc02tqv2Ih03IuHyYwBIuyOYwpcQxrqOL
/QTUsJyiXW/pUxhWHvAGM33T4zgeQr0DOCcYuoE0tUFzQ4kFjZIo7a98HBiNyvTp
ddFN1Rb8f3UhfQhJAtvK9lTNe6B1ERE9HwwwC2Q+vuIteofeSAq0jSQvjrYbQ+pf
pwQ0pqDH695yAmFvAdAgb9V9zWR1op/HPmFlNIHb61k8t3/rApKM3TAwc1p3fL+F
2lZ6O/dXJg+ssIwNnXDkbun6qEXzCszjDud8lg3dirEjW3qf+3cCx3lhpce8Ru6r
El7A4Ft1TFrKApRuVfFgN4ryU5bU0nqVbMMm/ceuFRKRAzARqMHf0z9l0WJLLmbl
2SYrS+nf+BGx3A583kl6h8UZgRJVvwCGEAa9PlWTsiBY9GNYcXEtPLDuwzn4T3jw
aC6bwJnqOL6t6zlr8OujyHvWLrGwwpPkPw51Jyl7xlrfOYmqs4Qc6LrbbbWYPv9p
yChTLh9pWCNbT7HxaEfgV+h8vavBQiNz+91JwfxWqkx3oKNz6BwcLZUNXk+ApnRh
dHJ7tyOLnzVXsHQ90zc6S0R+pwdgCYrX8n2hmNHWs6wtgFEoB8ibhjMzeLoXU9vR
eJb3AzVwCcgsZPBZ1IbzeCMuMibT2FjxNrgr1toDR/PMvJ5C8XIfpkvtZeqpNYOv
zQmEwAogYGg1YJWSzVTcObOV+F2MkehrbC1EKla2h+S7dU7IOiNptywnwCn7deV/
cA6ZebGK4oeDbgF+M3iAoXf/quSHNjQmn/0gKEgoF67iT9u3t/sLoxlSlfwRDSvz
NLv8Xj5YUe3YbJZ9XnUSRWpLl/bl9jnoS0CrxlsngHsYMKJYAYL2CHoEkaXHbO9V
PtPtUVqAbD2HSgqk/xdjh1a8j7YGRLgATxiVYsejwscQ+7vrAJi6gs2Wr/Bilg8j
jvICcCtf+AcOBM9iYRPs8zih0brtHNTgHnTKLbVW05uwKtAbRKsPR7SpArTtaLZM
lbQaichqmRSbATWtKe3M5rG6/hYhGi1GtQHlBwBqsAr2F8MNqlD1X1ttvtBnhZbE
kReSZyRcwrMYcWAAZOZPyd4qvpYW0ygs+HUnppBvCpYvVIrHhEGHp+BVF4/Bkw/a
l22JS8BvmBuAUOUaDKgrTpNje8za6mCWn/b+i4sJrrKo5sLOh+9DavutLJJMnNjO
6KgRvUZJfDF9LocKFGi0H+EN49YFqVrneUq62mnaL966/PN/S9eX8iXGArLQlN9J
CpEMvRe/CJmkUIyemP5iBt7kyClogsGRsptNdY7SZ2iDBtT1hZDdcUjSUDakTCiK
O4iCavUzcBzMVif5kkYIp35C7iIdGAWMDfueU83SQexOZgTXl7FM12pLF5WrDDDQ
3PudIpjxEAgH6jIDv4XgZ2lmRustY9SXwkSOirqaC6Ohoc/88gJZ6elXEeg56pEe
jZHBvNYWv53EalDT8Q4HBuZmM0tUC+nE0VtY+GZDXxy+/VTi+2Aws/KxSyyHhCoM
B2q36Z6KrjhxexVlapP2qjBN1RbKohZ+XHseTdsKX1k1xnTIg0JoCYjlck0iQZa4
8UIARI0ZfjT8YNUicgEXpHrfAHohcYSa/DCRDW8wqNWFjV5vCtSCeOHVnKz/vdBa
t2wMCM2s0lYL2szazYNPh8dJzYMs1kyXv8MWHDWwoSESXrccRF9mA9xhRZo9zbwy
eTA97cOeBri5mesPETjwKUK9W8fQY3714ZWk1pRacjpiNxen8EqYSnEqd9IwC1hc
vV4SLPm1L6Bvle+t0dvuBSCIX4RUUZQARDCRH2Li1Q0Lbez0ju1GSOcvnXGOjfq/
orOs67OrZOh6VEdrChmoKEOhgL5HYCYAe0J37ORxCTdQ9GssvegrswrcOWOnMCcr
09uYpobMcbV1Us5xVVs7txt6zZGCFWbAXn6nA2zKLR9/rJ7eeZFMFiofDiKAI0DB
p3/nEDUc5lHz3ntMuElVazsxTh4+eYyXawtyEa1hD4FOIw+ZtuoigLPU4faJxOjp
QOi95vtgDvw6z1sV5MH4vc6WcZw8gN87FEL8l5//30jKMCcqCwNBBrYoGAqF7CAj
WKThqDt3dMaao39k1+f1XFpUPLTQDktfAvdK9+K06O76YRBhaoj7Nl0j5RrAY4gS
W2CFZbz6HWaNSjp+/Q4ORE3mWhj1PE3hK431tkb7xQWucXObCBzrwCLZ6SD8LGUj
eaaiVpuFzSax3FXsTLcV8CYLlI0b3XvUEnswhaXuM7nfGnXxxm7Dy7AWypKbEQGq
iIeibtC7yijPYLo5oCdYErDiBB2jRgGycQg6vwONpQq/w8CmVBRanDBN83L9jyyJ
CFbn6qP7l3YQfrZOUW06qpNNXmKXs/0380b8hu4SOxfatBnSL9cOh982JUtNk9/w
x4NtV+ByGOwJ5M+grpHyRQvQIz/VjyHiN+CcopG4YdgoRW9y5b4Y+mM4xkRwN7Tc
7uSkfr6HdZlio2VQ704t6ZrWr1G9/dQbh0cnH69bMNJaLTkqcgOJ67Z2P4IVQeDr
D0zOdLClESM1oU9vGCOkx8a0n5KKBYgLXJrYZi85BpfcLcu8WJWnuqR/QsUqdFKc
cZm0nx3yn2SkDhPkhEvf9jE7Ynziramx7EC+TXBuV3An29WvtcGPyxDd9M9sWQqw
I6RRYoRtS1OuI4tdKUMttl6OA+66Y/ilCAkHHtiQcfryCQp4ZRcF8+ewoP7X0Pjm
LmTxa5jyveiK0DTYjMHb2jlwI+oQ8Ueg9MugZp6NF7vR1BEJwMhzGtl0/RvBnndX
Ghsk1YhvaLa44epwYQpL4ycMgEk3FxWzwpGw3v/mhL20VpGBvcc+bybpndnJjcRr
xrwSiYPDVqyV9V2q5HEMYFta47AmXZJkf1jTY5nggy5R+Np6i2brVU6DPom6lv3N
MeCNPVmSjsNBhqzQwBxqzmCplk1p0DJpBkZRRe8DU+JLy2EVxQ88sQYn2xCU/qrC
+65qcajQHoUzRzofyBKYxJXhqkgWbhKyYZTdQo/xmBV8LRzznF5miRZ4fsaUZNXX
J4wt0OH/sEu8Pw8D3t220UzxRMbOzKsTU19XZaxEc+FEX8w7qXBh2R7/Z8M1Zn4Q
WzZPE2Fsgifxh+JRZHMMd6R+UnDQ8BgCOqACODcj5sbzqHdYUbzNFf2jQFXVzZkH
HwHLH3QXsVuE/skamzdCYzR9K3F0j4laQGTvmhe+p8nyM37ivNVqCXl/CX5xl3sD
XDGMOGPLhzQa3y9fvTV7YJDkYH5vf7ShRIGl+KQNyddhNRZL/jAiPvirUNNCE/4u
4KZwdzZGy2eewHcFmp4WG2Z416N8siATB08bFbtfla8kDSznMiaYjgL1lYxEJ86A
OjahXrhFaCwlLxjX8RqxJuyYAQtBIIA/c8Hs81UdO2CvoElvF/S1j+NiVAqS5GTm
RGT9iAV3ZEG+6ZSrZJT+QqJqMPqMjPImk8Dv8p8uyRSmrPZhC3f32Odl0n7xjahB
ckiWZ+T4LZnppBqrerDN4bs8QtkGfiUk1nyCtwZTL31C3blHyxhN3HwR4jHKIvGU
VG4+u55REEdI6XU4XH/2LqCfr//Dvv+xMge62Dq/AT4XDAXeayEGIHKH2dG+aT4z
vCRHMWmVjHZ8WiyhE/Vl1FJROQrfSAxmO/UXIJxNpB/5sLaEfDiTte8pfmal1kPa
d5eOG07z9sygjDmYnrFtlAPL2qct2EoS4Dhw2i1j0iTVp9L7VVXP5oFx5uTJnFyj
mgGfTSn2ndwJRTmzN8chtJhxCRb/VgDbJHCW/eIjNJ5WMEo/yHIsfin0C2Trz+eM
hsaw/k+VBaXATlEr3JFQW3A43DwwwZNsKXFPVuTDRLlmxLB33Oh7htN2r0ozm2L9
rrovkuWw5UEY2sogSoR2nCYaBKFM3i146ZhDykRU5ZX2dxeDtz7HdMiLlmNQI5bs
7QFshkm1ngzK+8NxpqqwCRKTZg+/ZA6DHI0Q04xmBS72nlOcrqKBIV72n9CbXvmM
r2O5KOQv0GPMe6HI+DEleVKzjRYuD0PyBqDtlw8Uqn+xsqWgdOebdmYoX5xeJ4Bq
uYFjqGMGxZUGiaZ2av64kr2m/FQpebP4Tvv+/Yza8hLgOVWQtfXigHjy01ZVjNrn
jTZxtNEnCCLkkIf8FGz0wM/xi2s7dL47FxXmlACVSvHgKzsDGijKr3uuuAD0gT9b
h2T21nXNbElIMam7LaJ0R8NmTHhaAGTLrqGlj66ZU0S8fIT7DuvgzF9A/pOOI91z
pEf9jCF0BM09TTQrcRDYZV0LhyVgHaCOaZ5huQxPNDpQ5OHS0xo/MCQf7K2lNlkq
9FaFusYHEYjHuaF8QAmfhk7NwohMxo0upTs1/hM1fRG+E9ItzjOJvQ8Wpjp5LR53
wC24aKxf+jXY5GgcQDHFl60KVr7x4OD2iK5Omcqc4VobRXAl5L/nmuz6zt8JOayB
583IS0XNhXi3bqW1DNxCTww9fgaGXmLJtBuIvJhSBmZAIWI/+LmILw7eeki9bpir
oXJGw3kzz2v/4Z1xjDB8IA9PUDvi4x1BXHVgrCOuIcJxFeMxhh5AZxgK2oGq4/xv
WW34IBlsoj2xz493Jk2UvXKyDco7yv0U8L3Y2HPTlPVYkPy09JQDPvC7PiltWc4U
8+T3z/zgpQVFDQ7MfDYBx7j3N7hIXrmIbU5PQAlnPZfL6lsZX38eXeK42C48zNsw
uu/Oj/7ck4ThfaiXgF9fwJvVs3AdkOBoDcb9yRm4rhdQLWlk7voWMiyauKh334OO
Xe2rOciWd6GGJwPS/Edo0GhCWorwIL2QflGfqg9AZWFckyCfAJcVdifRTUQYU84a
xWaj5cLf1hEqRI8zyOnbyePikGengesVK8i2drzSPeWKI2tyUm9Ya3hRvRuFboSB
7i7a22FA7lHq7jBGFwzwVabVAHGaZmur1p47wHCWnCqrZ6vR7vSZ5DX4VmSsEuXb
sa15jEfVEpTrVCX3YYDaadpHC6Amt58ixstix8+Rpt0wOV9JgmeBirPIkF4qDUkU
VYpM3xaAvhtd4Fl8YnV4nw6dhuCWgXbHxVKRzChNwOPqtV5lcFrPMqgqluiq89pZ
xbhYllECcts+atv/hYUhRGnTFGDK0X3yUO4AzKwfascTBydRt435c2iKK8xafISK
1BU0qujmoDuzYtX0V9k1pObGefhBodFyuEjvA6S039kWOEHzbNZ5KcUe2pAgxtbg
rJ/jswUzV/dKAD9XLezl02Qw7EpF5KrSB2C0suNHTBZqvlSwIIj1BBkla+OYgR6E
De+NknpC3Q7IoIEMI909Qo0MDWnp0EiCjaGCrgx+zYl0xfATxSeTEObHNnqxaYoN
98oeWoSvoYY2JGdueHK7krIT9JMozkIT8Qytw2Jw7WoFg043dDK41Q6rM0XG7an7
+ptXkIZr7DvX3R7IxpVRaJbMgOEPMBtMpQEPbpEaIhlp1nQbOGWGoLXwjDOR4JDH
Hy2kQgZYhKvYZD5Od4CpdXHvZ5/EywxWFJx1w/s3AFRGaSJN1flKtrM9KyrjJIDs
8IW4sOfo2AbRvyWKtQsT3OSmh7UVnRYa4WNSbIj5N7+/v0QG6oZ5jTD7lZK6wXFN
5yay2w61UA4h+dGSBj6xUhf5EPzFIzZqNXxc0EhnmRs4frU8X4GEVhjErmsTRd3I
kaOuBrUIwYXXDMV4TblF3qTxHM38E/7260OiwYJ+qgJJVToOi3YQI8cZI2zjSzGz
CIs2RAM/pcPnCFjjSYuIp72mPmZNqtQWunBZACSSU+FSEwCl1de3oTTtw0H1BaN/
tyMm/MF7var8DQYHKaCfLik2UPdDtNqGI/M46sP6Zs/VVqJw/xv1Ggu3u0PAqXW5
02/g0fGsqBLqmyKlp7zAcA5LyVoUe+m1V4f3WxYJdMWlDsWaAYgcAgl9esGZT6by
dzketexUC7P6oPrYbVMZzzZMi7jVfkYhsYaeS4Hxhchzh6rhPHyBudjcEvqw1fVe
tePdoWwq96JU2DzVKsDim7b1OaU12XlITDKdaSgkMFfv0ZM8L07s7KIm2wzpEbcj
bnSR04Lkr+01YL5/Y2chtCKE1HuPCledJslHTMyQjX++aKXHRug10nGvOTiPU7oA
DwrZWxdYxXVtvM9nZQ/d9DWR+GvzcqZlaJ44I/xZJH8mOLoqArYpnAw7FZzzOtQx
auXNDzBb+dcPhmHzhbrsvh4yZQdzEAq9X85tEHUIJDsH0IBj6NXmWWnMIK1IfuSM
aB+MxGKXoT6zvSJ+dw590WHpfNuFIqkaaF5BHBVAP754x0TayYzNhevGD7WLrSCi
Di8rXCVj06aZPlP6+44GVFRjaoBohkGMA77NjYH2SoOB8cXM7Vo6OjFryeo6mIPg
fslXqy1gRSV+nQskmxWD9ubXJJtPcqvOQ4OTW/vO7F4Xrcq3OUIfhIMRsntp3+9N
xc//2Ly5ZJX4ehVH4vgcB7UxCkHBTxC09TrjIGLYi2aKtJLOMfrAondId2gmxuK1
6WzaqfIvO3CB8FkmBpXytpiom23Hk1UUH7I9TTdytkEe3NNSekdy02T+GeD728/l
10YW0f/MXEOjfxm7KErjygZOlODgmtnpOqkrIOxR41zjYiRiNsRay+HDimB062xE
D4LRafjcBhKbaaHK1YesrR3RkjJ6D09zeJuRDoa5TqUZ9O7kor6uWFZ5FgBQDP1s
w8kVbs5LGiJUnILSF68kRxHJJHQ+iqgqon1Cj0EUjTmejGNd2Oq9IkLsrZ3wnRO1
Vgy3dzXIxhZK+5lFC7WKn68bsWZ8JHSFmLZCx6LvU/4NSejUYFIXXN2kZPivPDno
gJDGAQO+qonNR8GXSkSib4UqplqM3GSUKwxOkwldiVruFg6O54YjE1G1zXvz7qn/
VT2mD0TeUfv1UtrlTRgzTAgnsJnV068ClnAgcu4qtj7MLiLWvj4myYRx79eQYg0W
jUpkdBRZYgjLgIhirQA8Vz+fRbORC5604haRtpz6PNQQxANnFq/9HQ7eS3y9BRkh
hs6kpLTRE30SP0uBpPY9mCyCjNnL0pOMc9IKO84zbntXFDIb7EqYczrfcr5srqh3
qzPifHx+pUWSIRWQEeCs3+PgqGJkL5JFEGI1zMuEIP6H45+WVNc2TRySYTQIs5bp
zM58sgnWA5OelRpnpu4ty94IzMRiVBx+A1HYsA87kyupS1PaOwz0GSY7GCKH0KAJ
hGElA42qJsDgBkaggu7JhgIOgA0O1wrg7R0Ls+HaVGSGY/KzGpzhGcZ4hfTOkr81
tTAjpFa3GA+W4MdQWLmAEuhhLt2d/dmkXvIILGSBsgCujYKIXXLDgZ3OUrtCmglY
9tE2GjY4E5TJ6zmzuoFHn+7lNvg2iJwSOnK463+p0KIRAPCoRodkcQ+MhzIJ5ij6
aI/ffAVrQoI5uMLu5C/NUQ5MBxEqSEVCbV0Xjey9k7B1tqVb/u6Bhvu5t0IPE6tE
Ie4sGG2iCMnREOOuy3guLz+Rlgp+uPQ97MmXU86gFPzkSCWYaj3yImLeUturo6bo
Tz7F88bKumCAcmcciHJO8OAKPyaBhXl5f2ZB/Li/KpqNfQ3nbMBfSNTe1Pz+wMT3
lpWnwnwVgVGG3xiAwEXRq7xePu+X8vpEHa+Th5esy5QkEJTXB/qrNRzQ4VJy1vl/
gungMOSpLuy4PgKYk3f7T3LB8JpXlsTbZDdE0xrPQXLr+f1o4kNZfUoS7HyLzBKA
lUrHiLvcmFpA0qUH8WfUw4rS9ZAxyNZ4aFHjIVaq3Hf0B9HfrxnUuUqOn2MdIZYZ
7cpVeg2wBRQ4TA1qRlcW42x9hAvNuDg+dE7wKQsH9VmltLl74QY1kBizmqqM7zcu
ZJRjqUkJHAcqAl5lRnGRz2qLeT+Ef/b0dezPuwkfek7sukufg20RcQUuH6KYjr+x
dG3tXyLWOdhXHt5kS7r6/VmlqOm+FxSaIQ3qc5hM8cyoWbUitLanAnG1AnHjr7tN
BJo48Rl79xJ9RrG3iBXhVYbw5x4OhXNgTVuRj3hF3YDX2SEDyUd7yc5vC4+auJVA
wDVBxjbEBl+wxLbm7vqjf7YWJi73mkTatW37UwzwEwxbXAT8wCwJlTobNwjCWVa3
HQ/+dipb1S3o+a1kWPSl1nJZs+2NtawwzI94a9mQmbuxmw/1sPaSao9grYEcMJRL
DxINyQ9pJJZHlwSnQtYyqEr4M6jygazsZ/sE6CeEou18x8yyBM1bV6Uhq9o96czd
NCbtRp68GvIvFNYEmxBUp4eRf9P+U4Lr3iwqEe5U/+Prcsk0Jjo+4d6dLOnAV1dt
+gIiSxqJJHjqaFW56HYivEwqxNsOxZWWDBdj49/CPGW1/qBZZvQ35CU+q6ovrlU7
bGFs7t4BTQF2WtBMpBRT5kXiHojn93WECe4qsOLG8JlzGmiQDWPIlOVh3RqdBZRf
zUNVsr+yehbnmH/wCnnKu1BPJBB2OwcbTc6+KoKOLaK5bgtjjhcSdBzCZmJ6N8LK
Oi65A3F5uQQooegHzrMJyynaICyyBFhdFONJrwPvsjeOlm+3QMYKTWHXZKZo2qxR
LVoAjQ1U+jyWTcaILpbZTXNn+5QcNX6T6iKhyGZeUoM5opa+G3vVqc1Cpuwh/xfO
103UlNlcvZntT4HP7NX9dHec7slZjiUleblH+aTaqTfN410HnoFvtOgkFRz94ILq
MceV/+ymqlF5SQ9v00Y6u1617xSjZ6pjC0OzsFfzSW6BFk6oxN7d3F51nKrwjWwg
M5HF8XW54GmuDykDTsQ8Mjv/dn4BbYaaKeptgcg5Du2pnEKbjNgho8WTPSLzgu9k
bUlRgYyCEbvnBmj9lbhPajC7EqK5016oHAV6C69yJ35ZbVNXT00z49sGM7tQC4BZ
QI4gg22lF38TFHi+GRxj2v6PXVTlgAi4Qv9kb6Ja7tQcsSyRfZCUNMGhiejPIvl3
Up37wp7ft74Jx5F+Q5yo6+8Rs/qfLQk9UhwJ4iH2bWMO2ekRJ0O0v7dKlb4uIOLD
vfD4Vwx3kXHMGOd9e3MGEZhsHPNiYSMm6pvYJJ/1v5gZusPRkuzxKFpEKN79f6h5
ZkQc2g5Ihoooo3f+pttGyykDlZrlh+EFprWz0cUoyMSV0YKwvi1Fa3uc34YOenyq
M9lqnOGirPTkC1znwy13VBZ6yV0tcGxurme0stBjqhtoWuLP1o+mlT5Tvb+Kvtmg
QLZDKohJ17Ze3WbKR6zoTJRdJYIBC7dcpeFgVaTPb11r8g/KMZJEplwfloqz7dYp
4M5A/XmNMugR/vyt28/5qKXDdhBYJcSG+o+h5fIFUkF3ihdJmV5ZRBVOk+mC9ZZi
QJ+c3+aBmZRujppEnvlOb3AOFDuUeUqRBBO9WKTlzUa5ZOid5w+ldqJrliq2sQLd
awxTqe2KFQSQTF/106Vi8k2SK8N/ViwSk0HxqnQBudplVpJqd5GoGFkCSLqlcLRR
o1MW2xWcfOnCgcis9HTM1hAtPUEf65ZjfAbZUvMBHVT+WuuJ+2Z259nk/0f4n/rD
rH6smMSsv61zefMoDacfZhHf9gulmSE3EYiqHn83ziUbYMwg5A/L76ZjT4XdxC0y
tysVU2E0g5Ohfx9KcvdZnqJEy7iVR6RtWwtT4FcOrDedkWNo0Yeyb9P17RR27oCE
ELDPRvnnkqdw48ib1U7hDsbeFstTHxdJDqChkhXVEywTdvdhfnsN9IJ+p4Z9Cgb+
Vr1dDxPgY3IizdWxdmbv37nJCSuswXNWjez3zyIRnz+WKzyRbWE9v46QwpQ0H9b9
J6aM1Sw+NiJ7Xnq37lIdjtTEKrkuJPuItJzANqxnH+kv1i3YNRjgiigYQb9oGY2v
JhIuOmDNEzQuw7Wve3fTQx7vAghXI7aTqc1LZHl9tiqcz+vt/wBCzYQgUbw1QXBh
5nNprRXwa/mFUCMwMlvDo+FuhO04pbv/etkJOpc05BfifYcrQ7gx6m7uP3YCtiYt
nifSE3KwKiPHvgCqFfIWrdsHFoVXPjefBhIQyua9jy0wAe4rLGGirHEooBfhde7d
Bjleeku+ZwfmgzD72DJPd4NeR6LWX/Ir9agtmLn8LJ7nNejPU/TCAj5Tt6XoPKbD
ZSb4MZ+RWZ87zDm9bIdkI4mgXcJfBRqK/ifOuP5oZ82Nr2m5E1uAo54Aq1QowwXn
yq+wyj+FeYnzZOfFx5RQ3mzFMx4BqM5ODyhZ3PbsH+7POhEeMcotWxzihIWGGGhf
mP+lUSBW/vpX0NJcKDP7nRdjHcIhFaHkf31wlGDcgKOOxNlmtBeLXh1YBQI0Nf4Q
Uo9dXl1876ttfqSlKTTDmto/S8P1sf1aYQh9Q/vYy0EkBEA+rgA3XP06rN7ttcLm
0TBA/PIKGKXEkVd/j7SiUd2+zv1U9EgPIom2AK7B4Qju4QjAcu+qIfn0OIzKq/Qi
pRSM1EAmxLbMVGOibGVQT0FHSxeQJ6z5MQWlR33aY3MlXI0W/y1+2EHyDn6I9Udw
Od2eCIv1XhV/m7joGOcBFu/Db5HL5mTYKO2/Ez/IBvMYRI2Pf50DmZIdK75CtJOd
mXUW5nsqXUAh1jkHajwzMzO+QXHfCVf/lkigQy0jlA0RfhbCre9a0WqWVs2PweVJ
/V330tCGO5Zpa1L0k3EQAyKNdgLILfPAPNdXXPS0/4LhVpl/MBgP7CbOIdWrawHY
lTppllHfqf8UlRlOZfSoTGHQwCYz8dCk49gGr/wP/JA/3Gl2bYykRT0GH49+ODm5
18uBh5HjFvFtkwDtYjG4jFCDoJrils0cytZcOJMbvLh3WZUiSF5wqp8ZomWlaIWI
gZN9sOt0MLnuI5hSoNPtowC3eJCNgt5yibrTQ0gH6wSqa94bB4hnW8iLLN8/9cee
t1D7UAJwaRnsTvTKAFcxdXFZ7ERX8Faw0EGH2ZV/lOAabDx3zkt23LH+K+nDyGeY
iitRp9Um0Z5vPpvAzv9hJxTNQb2GOjTbDitbAhuO5lREmsO0ybDOvlWZxychjqEs
dMlfLM6vkaKDHqjYI/IcK94scK+k48bF39tsJi2Tia2hhkOp2mAbGzuD0xrY7ynF
qIm9Imm7klQhfT/G6OHbJIo7sQaz1LuE/ImEkTuBn0dPMa0kKCoOa38ryPQlZ4+F
Lu7DOMay16e62kFMvO0SgzjWWm+Nlu+PqHU4z86QpDIi+ADLQ0xWK6xblSymayF/
pSQM/NQezPkKjwdHGmS/yqdB7ZEVDt6022Oia3itR31TtvFjZ1AJ3nzFlf2deNbh
NGjhAnYg4wLUMO7t3pGpbTVEli9V4p4Rl+n2uBXruYrd+X8ecj7qDMNUuwupjQRm
NOPpvxvRfX5giF7keFKDQimxkj1BGiRVDNXtgKewVeQjbscbFU1EG1SylOclYTXR
64Dr+TWA5LuavzpuTJXKf7SxNHMchAdTHFL3R7G4rhJywg9zMbczcXOvbIt47FIu
l33sNzqjCKKvtJUQnitMWpJA+2yLx3ifR0WtarBK2UCRE8GVfqTYWetBjVLKZsQD
0M3kiXPBttrSvP6Fn7e9Zw6Nd5+qaVddSt+zgLI4Uz2ZUQmsmcAkzoL4VNosz1BQ
P6RGTiPf8aznGAMubUlhPJ0/girHMFS3+I9uDMU9EVn45Cqe6INw2jUYVYZzjIOn
a6jRRlxlNPQqQvBCoVGki31L7sjXW1nJZrGfK11jZK3rdckjFlQxDRnZ90DotqhO
JHjU0IZi32O46cGnNTwxXnN4GC5qwgkMYGcD8Uciwv0L7iZhzm9veXKLLBa26ino
C8t/Drz61nhy69oqkdzCsKe5s7TWc8ZjnzbZcgUusc/KfJQfCz4e7usMg96bpDiX
NckH32H3+db+Kcex2A/BaUppu+NB4G0bdXVD7pf8Ff9PkaLewhzn4lpfDJIlxL2Q
wq9IfIgmRaNVr5Gi5GWnXK5yaiYZyFkvAj49f44VUW67DlYb6+L7JyPes95IrQm8
MA/Sppoa0AJ0nke21pnV2ihOhAbOaHzQzxB31imBNUbk1NGuy4DsXtaqm73ZQFRS
z5wK5oQYhi2cTRajbkfkJljay0zJHu2Ozzdk5Fi5cNClOjFE2mFulBwjfDVApM0n
lMMeKwL7NdbCeo1+8GJxn2PFo1fs9M5WLrDSQHoRemHwcbiNUXqOm6WneA8FrGx9
RIhyxmXG1abUWzMxUrvp/5mJEZvpaLGqDJOf6WKJexwKqvYo8wnu+KJf6WYUXq8s
vd4Zt8lCXUo34swC6HSjNIaVFMv/LQ8tndo3+lbImqLHzrz/hg9HWvTNt5nOH6kh
MiU7nX29L5ZASoXo7rAweQ807BVRYzQnHLcNNm/BEng/AN7Nwqe0hyfmT+8W0daY
+xJccAOw9SdLG0Y8iXEFnPbjLOzY3wjluyGRqcW25csj3bqVyNs9UOFs/Lycf3hV
0A+1Ve8EsyeT3pim0lS2sXlaxLk/rjJbKJnHBABfB2Kzj+2jqY4wdezKMuvriy7i
EiBMVXumfYGRUp8hh0cI+Ue5DRwZxaKxsxaqi0fcVvH87OLo32dy015M4yyAAhe6
QOTSOiT/+5WfC7+/YD0DDkVNaRfkpvuroNjydBTCSDrBurI8JSIOZUQzXn2ZgEK9
U20ATNCtuZKnra2MGepuxtWlN7amgT9qyB4E5s/4A13L8VADatpBMsgntLmfDNl5
/669Kdju1PvhyUZTvy1530Kh7YvGic6lSv49WwScVT8zi2D2rPjC6JB4bz25xqFP
WzGwzG1myG90nAaN/ovi1z+UNHiKDHXref1ABZmnRDs8lqIfVvmWso7AgtrsEum0
Mr9stfijPGpo/Syf0km13qcI9aQmFbWJBUsv596WoatNa962QEyRIHSXoLWqU0El
evjlEmmHlth56jqc29jx9rIcpjlOWEZipfJYYV7eo8e9H6aQc82puOMdGUd5TX5A
rmmrgjYcVQ7h3BB6/VcNUZNB5mRBjACCMFk+tRQYsYg10xNuHT5FwIioweO4pXVJ
bNU+nvnIy2n6WlJMSVCrfW+yl1w/PXMk6SIv9/RoUzp/Etn6ZuXxyK8o2FMTXYin
bKJz5QbmrLGSKxxAmK56UK5AR0cO4kLZCn4WOggnrktQT2eIFLunHrv4hdtRo7Xi
9+nR2YfnWt6y3lx0fotgIRuxEIev7dRv69/OoU+a8GtHOPWHfxLX2auQ3Z/2qvKI
RuffJaeO8Vlv941WiOXXlw+dof7qP5NI0bcQ59/wvxUKWZp5WAgr4OxuixzE5sRz
GtOqMD8X29ao4a2kQ9n19z1VG8kNCND8al/U4KnCLOt6r3QiNKy3nTTb/hLlcIjg
2owIZH0jCq6OYot1f9f70X5WevVBKb3ZWLhgQrnLccYhNQuLOPosg67CRKcCw0D9
blqofjaJUzK1XKoe9fW5qMUtvmhS89e/vrpbMc/izyyWBe7GbVLiw84zKUC3YtBd
BWjwiQRWrFR6AG+BCkQkFzdbsE8J/+kcYpj99AoAilU92o1zw+QA3cs2RWhYxmsQ
+nZrTOWjLdbsBJKir2dcvYndNumXzty/EMizwCfjNU1FaWy3Gqls/MCi/raYfL5z
R/yelRQ8AD4nn+b+m9dzhGAwjhagdSUz09H7oB9bJMpTemWQlmLPWHvdjMbCEj/j
f9Q9hS29ogseRkrZ+F06p9OziPxpo5rlTjo+d2PCxV3u04T8B7gA5LALXL5sXZD6
/8+ZK2tJiO6PQ0ksG5oR2Y5XbQPDJBQTozcaHw3KByJG+x+4VD67IPKK5LIZvP+3
I+y6l95Mtf4WDRm7UD+ZbLcAH/Hx45DUL9ECyJ+T3IB4yqda8XB2hob3xKKe8STC
IHB0vdWaeHUJtuhSVkCgB4gir9YcmKBS5GXTORzmVYOBXdCxue2l/Z5V7a6mq/T1
VDVIxdwpInujiy3CsX4k58spWxWR8KRfe72kXigHufR0AL0t6sI9Upd9mGcuohBq
snnSkD1Bdq8eqXr6QSLuV5R2uq8hkC8Z9fd1nxR5xpq5nsING/DFqfIYHVLCC2Z0
w1MotMo+e6Unk7GbbZE5K36XdJFeb4rxP5tXfBZpYwMITW0jP6g6Zpm8aINgZEoU
IZGwQe12ubAqYGKnlwDIvTnP1/j4jCjHlLDvsnFxl5jfc+gUpD6jo9X4bLepsPcG
ChjKfKNB57G0PHHgQbYLM4Smo9IWwSuR8Ii2C+BNZ3dsSnh3vASOqaYsoX818yBS
Or1hLZLayglXtIO2EyJ/mwmMku/fE0EeoxYVAJNtkNmYZAtt0eq8Q7gHvbUyAc5Q
QUOQwKR78JGn32eiRk6HTl/5FVq2TzbhRmjQ455oHM9vMjxeV3sBGHvS44zJilKu
2BKLfAzxmg06dW0LAjEFAcQMsPnUXNFOY4iRLDeODbx9qPY8POoVGRh4bE9x1Tin
DYrnrrwZqU/1HTbSSyFzU2SbuxqZTfxKEJ3qU4qk9KDBNSGUnFp+jywpbJCH9aN7
7s5+0bQOPkdQTcGNr/2ABINB9C3I1PfRl0xnofUIkMK0kOCa9YJYwvy3vkMflFXm
2PFkkkq8xLyuZI2+ogohr7mx2Bj3R5LlCRI5L8FrWFP6JuW9mMSbo362/XilfXj7
ZZvYyudnFPnr5gTETnouW99LQ2eO346xxOH7POlooJtvhZqXUtd69TApIKFijjMB
oQQdPCOgmKUPnETkcS959pMoWU/8rAhafvwu4pQ3l4oQTkH5da9LS+WOoMCdJWv+
h0oamO0LxF6m+s+gTrP+uFSo7I3GKoveKNsCyT+q5btyDq2NKKWnhr8aU+PFVpjo
xquSw8QQBg1lg14+fy+pkl5B8Gof28q2bjCu9r7hk/qOFcGyDUJrnsXGdnHRkXIP
5mnL0aMqVYUae9nMjUt3yTxPWYy6paQ8uH+wRVZXR+6SP3l5iiyiTty6WxUhi8e/
OSvoScSNm4PQaIOv6/BHFFDlap9A1cyrJRccBoE2KcdQleh8j/Ln/FceeJJ7bNYP
bp9WhrLaUBnCZlkYfcMgZbqwajwmKbusC8cYUJwHsJ39k1JfTD3054bSiOTqwB5z
a8CkF8qKGKhz5GRTpZuwLttdmtgVPjMYL2ynlqXu3b5uJ1UgvOEsWmBqguk66szY
dx2/IsU2An+ACqXWovqRh8+y0iN5CJ5AkBVhxEjyl7DZJ6EGS9yzsr8H51WcuW21
QRdUm1qRA+7O/frN5FWRFOb3UMxge1Gtrlgm/7dmhmuAu0jYtgKCYv45cbpMhAuX
4BTQKhgB2coDbzgY9/bhIW9mnoZBXbSRwFe50QbAIu/2AqnpY42CMvpNsmDaOCHg
yiWKZink73MDUKciV1wfTbPoS0x0LftOXs4PqKycfStrVJqtLuH1/ZaDWAzeY2EZ
E07XvrB3O1S1d2D21t7xQDTYYXSHTXTj0MzDUl3vmwFYoBS1veI2ZkyduZx7m4cO
N67dtb8f/sZAGf8ZnfXZ/mGVIUHDH0YpnASp6sVsHBfPF8eCHUBDB+FD1K0zWCda
inmkXFSiLwysjh4i/Ezh/cQXJyg4uc3U4+z6rvxwc5BjUvKnd+KoOowPBf9PvAYc
ifUqwFOWhvgeoyWSKQWvkMDAqcBOHFu9p8TX/WGJEWourQ0m8Jm7vaUHiqdJP8l4
vgR4ookkDXcmEmWDBy5exqELkD33R4gTdqLn0knMCDBh8Gb2+j2apBN4lxpdSLxr
adKraZ4ad3cTcrt3GGZ0mjdAzT17LW6ldBhdtaI9iWL7/+pGQihjEVNkcrbZmYkK
Q9yAh4fJeDQyxXPttqJOxPH21kdelo3OFQoMTizMjdJrmyGmMXY367z5bHIJZIf2
BEC/wN20U2Uy2PwsEz9+dOKmRDGDsoZxdxEM3bEzTJW4GNkKWhGH49Qa7La7X63C
GctJcgqSg7HMyx704OXqs/vd1L+oO5eJDEE900k1tMlEdPqvZ0LQPjcDkJ93J3WO
YQv/5fLW0K57AjStaKiXNfQp2HiG/keMMWDuig5BwG/XKEBgUuQ5ysK6L8e/kdJx
MnCucRmh3IXZucKmYe1Im05pLfyRh0BT1wRZLNOGLgHPsJ3Wydi4ffa80NMs6OyX
6RwwbOMZhL7xuZd7jVqO6sCYf9SpA3Me1qXuAVJ8y2Ix8vkN6x7lUgCzfGvibaMf
4EaHX2eTS1KblmEY3aY0Ri340ZsOAJSgW1avbhzblcOh0ly5XbIAl06AD0oad0KP
f205huNxFoVZR1QNmiUzZu4xtpPfPCF4UDWoR8llCHL92YM5L3UpZF9xgW2sP6Q7
ndkUqzpimhg9Ars0qmitBCKntm2O1/CkdkvftKQ8q9boR1b7AzGlcFwx5xGu0Vq5
DfwK356OuqG90iqQi2Kvqd843v6xge3R93I5QDdGezFn7mwFUiKBiIl8nx3VAUqo
pHgtDkdRz5RzKlKWZ36wDvYxNmMrbZ8s3/eobFX9hmRDaH7XbqYvmKcgZHONodDQ
PD4lY+3yz8TnuQPDHiv8+2FiScqq/PD3Cy9gc5Dmi57Vz6LUnbEjNWc7KOG8ZKjC
OUivg6Jx0rf1nOvhCcAGjvtuknz9wFXbyD23F8CKzyXjsSzDxxBGJEMrWBTwZdLg
SCMFzVmLef59Gntwq+UUY0WsHmMLARVdIGHN26EYJLc7TeIr6OwMibLUEegK51Cs
UBL64fB+9gRqVUWAkpde5Eh3U1BzBBhUten0XPyIkxXcpudNmPhSdqu470wdIGtR
9L8QmsXrqdayISt4CGPI7ip+9Bp0pvMhLrj4VpUWenNXcZ/rkFjJcXd3mDYP7dyl
HhBS+WjjwmF5gPICMoC6tD2WOt0MrWgG3MuEv2zgu3hWf3M+OlNQc/08nGuXmwdO
Wo1rPQ72VCXxlvn9MkPrAiJaodbnw/Rso5Cwjjm+h9XiKwsW46UEvBSqxHyDJvPw
mWqBZ15ku9+V92h+KaZw2+zSxuLRgPSoMUscWE6AojEWW2idNjf8nG12H7pDScog
e4ZhTlWJoz3zfbwRn/QdAKxJ4sbki2xJzrD43VsHh/AxLsf+az5uwK7RCof/q3nx
dH7t5G1Q0I+uWOc9qre83RtmqXQF5uA0BYwc1w89qZimLjQBml3Hqj52FMau24uy
xTCTuELOC2aw+nMe+D+eEQ8RWR1HBfLczoC/+GQ1G1t2IDeCb0UImcekcfsITdTY
JuTrTqSHh7KmQT7FHqIvAYOlSbHMkgd/0oR7ihLQjope8qFFpnuB6+rC5idEQOp/
KT/FjLVioIu92deTzp80lGQi/5juyBKtWhHJj1hNZ1tOaY++8X1e0QXcJ74Dz/06
B/pyvrt2tAc/iNR1i6jz2zi9VtfJpvAPrqEIXRXRgeH2mKKUp1d3U+YotI9xH6Dq
WaAxGJl1j/UtwxlEUpkv15hHwHZwfjADm5/C5hMV3RA4veprBe6vu/R7LgUlben2
KhJm3oXxtJ+N/23ePk02dJQJou0T2J85TsePnTcKqMy5I/CpbmZ5f1KQnIhS/UAd
2+fLZRp6Ur0JSbCsW4mut/9EV7YOFRMXBjD88bofVwShrrhp4viE0+2dJgQuAAb2
5j/wfv5xZk+0YQn+AwmRfEc6BE1bvu1O5ml7Jb8KjIWGRiIBB3h+i7iDFcQ2lzjL
SvDlnNtk52rYb/VTlKhr5nsXQ9SjQcn7w2tlftADO6ldODX/LzB5sD4xZX2vLU/X
uOAVlr7vah0DNHDH/54odEBnw+GBK68Vy/rn/PbmjEZV2uz34BM1Jaf8S7FycFY3
7HPR26ba6V+Q15RUDOQrpYLprwWbDhtyLcpzX17W/FORSgXPb3jdo6KUAdH4Nd08
ok2wyx2QghbRvakriSjNRh1L6p/dsoZthtGykKoT6HDhzLSi2/F2t+z9xPXG/G0T
427miSTqi/UmoGw68kH3mtOQcsjprvpUUI3DZSK4kz7AaS1keeGkEpij18aMEJJf
KgsC1Qc6/mBeHiY2Dfxr4NZd05kXQ+NBBjfZkGkEVrAJ74Rd0PVLMASQho0F0ULI
tAmFMHTH8RE2Ollr+AFXkS4bdRyGMLrrch/HaPmP9vxy9l+r1t/bKgw0LACMxZRi
9SdjJjZdAdzCDF8QtpWqMzAjvqI0B6iDvKnGj3JpDKQy/hGNAQKeGOW2UCcecHx+
v/WaMONMDobRp34gACaJSoj8IGj3d4X82/YBez5pf8mCuEiWhQ+O941uwIYck+eI
KwMkHrcBBnbiQkS7lmEmPEyGYANZK6ZEdRTrnStNUr6OQVIYitKPtTDPV6dsEv6A
be9dx1F9V0MXlMs3o7fYpov8entJG4CtWNSUdevJIGwPTSYvN61DfLIJ+hIeVm07
VIqgI00YKE1CQViEwm3rUOvOWnWg7jKo3mJ1/xSTQC/2pNQ0aIgmHPup1wigCKUZ
I2p6Z3cyI52WJvxygUSp5v68O2D3gQ3+69ubSTegXDMFSC9l5PSNofkdX00wnesM
rJF2AgAB9xHBj5g9vFMZkjFwqxLku3Yts/nppsJWn7DWwamNdUfkzIOOmWR5lR1X
3FvR3xBghy03cLCilMLeAJuLaw6xug7z9LqTm/W8r012auzaEo/ooa2EP86urQC7
msZMNoUb/APXhI/0EYscy06Fn4xSYPud+6D62Ef1yJDNPiKp6HilXhj0pZ5kIIr3
rW3sSlC+Be/1ljSWxxdCuJIERebOhdDCkFk5dyS5UZLjkUcMuCI61Db+ucnOOUzG
+joXJwOzwt3l+8a14NNYvTv/kNVO1PtLJgKltQM0DoVOyJlTyg30LvOofcUGjdHD
Gn7v3UBcqVSZChVEoTT5cYlNnlt8fl29FvjsS7xVEVlDjl3fX5Nawur9uthL5orE
3NHB8tVtZAQyMP5mmMVLiRWkJqlHfGJ1VdBZJ56W5YaZLnVHFoRQiE9l7ZfMH3+f
nzkf0dlNql2rIzF4J/O812GxmxaHrDNYyHUYouAYEFqWOAX/nTbgfVM748r9rBBM
A/iYxDTJf0Ow2gbEIc4R2xbtEHgBUJnVoFUv+7CSxXJb/PiKJ1PY+h0uTabZyhEE
WD4vl7GoRqq4vck+ZTj7d4A5IzfIPaOe4/KNYLN80pqv75GgGvkXfQuT+OlTFN8d
C0IG/MMN4KS6sbAoZOSKzogpayFXa/sf3YECp+RZ9pP/jNxVtlUh+wTyVHSZiaux
4uNvwya7stKBP6MK63NZMFLK9+w1hE6G/ZKHQl86jFO/mGGrtifodOK1diDEp0+z
nTaN9Q5U+Fdr/FLSX7I6pfF4uXUojUII6mKUrv/RydABsqcEPpueLMmvFf2YyFFm
UClWbTpLP+DCQ/ngK5vQiaGUD60kY/i9J66rD7AWxul3B8SURCL4V8+rO1SOSNXZ
mLZv9pRbZVF+IXyYBlAQdc/hClUI3sqFNLGj+pTBPmz9cRNV3lel8dxNm/0RyPQL
tCqY+Ct03X/XJ3T8kCMgIGiXxhDzNnKol71KrnvFJM1URnsRZS10nJdnLg7fmT1Z
NjF8RvSFwLAVviYybzbuD7JTEXQ3zO/jfDosyxNhYHC8uw8rUFa8LBjXUAmd2fnH
DxxT+4fpdwmZoJwGTUsTHeAmr/7WmWRuCgK1HtAeFoKVatjDXEiN0WzmY06QJFWP
la8fj7Wku1eKs8jhjnaVjW6BUaDdCjUZWKsmjconLQLtimNQHZtR6rIFOvIfC/55
dJrm3gCZrI8EitadoFl3pbHOkv83Lg+2b3WeRJXggR/Hulj741+Q7pnZbf+zmclN
MjocTx3wPmWLdUx3S2NEAtZKJSeeP+x9RHmE6+h3YQVh/H62Y9VLW6GUw0PB/Uz+
3wg967BX/UWWvpH3RCqBeq+3bd6myUsyAqEb3q9E7McCJEzjRHN3y51xhn9n9Nr4
1HLOezu+wLiFwcl6ejDWyVuHbO4UTN7CEH6mGpI++KjhEtSIrbFORCPws+wALwk6
OSGL9Cwz4U4uQjoMza+8yLBUD/eh+JsxKpJrs8oGL5/FSm2uxrsvn31JWOEgEYq1
FN+S+0BlqkhkWVYWE062z2YYfmKIs9m9zOg+6x0lMMLW0sNJg3IcNMgRq2/ynwWP
TfHqIvmGcHlvOcX/kXrHevFyrCy6F6qgg53dWU2nPtLFcZJFowgeUpay6vul3kVl
6tGU4KGzLp1aqtWafFAuR3l66FNflIvgqli/jNsqmJG8+2RDTSlm4x0WeELOOxpU
gIMIr/I5M9tme8PMcrVWk3eGRzASJSse2Oi16BTbY3qT8Q30e2P1iSYIgX5UoBYn
myIfbtH6512HtFe2122FCAUimjuFQuVGzFqcuLVJd11kQ2Z7jubQOlIMahh5kNnr
zjwvTA2/7a0O6Pq1WUYHlEaIfNdKdguNqDGtMIB8MMHzoayrcKZlWvZ/4wRPT7+q
UU1CDyT9fMGrBnc4K4C4x8pzWYs7cX6uRNRmkxdChLpYlNk8tl8QXXW/s4VpfNU3
8eABwSuZEFMks+/lVk9BeX5W+jPv1gECKbW4dHuL/zFKiPMuEgnzgGC0mmSyp8iJ
7o/8lUjq6QtH7oeD8GOlz9BE2jNr+SCXCDB/I+ZByDdCu6rZnWAQgK9stEUADUSD
jz9dbtUM4He89SpxmmGZa8YXj0hEapZHURQeixkr6EkaH7OOlhSSsz0nCGfkfJQ/
PQ9BYDMX4X99enswNzp6iXaBK4yPsdAUbUo02D23hw7A68ME3hpWUAKl92udqU2J
eNsYI64fkRKpNam3ZYu1HmWEDE+Nekl0JNcwhtAt2AFvYOKb/p5jZCtw1aBpf4LI
4bmeaeee0AEIFO69EzcJkGmK+qysn47nXB9gDWpEurmI4jhcn/hq0QlnM2ZiNsFa
zuLY27cgk1ol18zux6TpN+sSx7l8SlX2NiOBenHLEP7sVX5w39SmxJwSTX9tt6Hq
F+DEnweggwB5/Hc6otkS/rzZG8Lq5qDhc23EyFcZE78dBSkBe5ZSnXBXmvYqnDAZ
PAyliaWvHWAl0Dr0EmqU/fnWjEkW1jWADy8Gfi2S5FpV34abeiquSMj9PDKQ/hze
2FJ3D8RGTZf047LeRmuiHRUN41w2TiAjX7cBHN1NfQ8tM58GTICEg6hPALAUD8ky
JmFMomhWFw9zU0zMNlvvEqaXPFKMUHv/bGSvf4Tp7ZP1Zt1sRvl/onQUIBB8Uq/M
wO4ktMMm307Pg7aF7Cw4LpufX8hP1hYAdGB8TkLeYBKgelEBxFTXBdP/Zmq/eDmu
IOncyII0vZy9AcwLIVRpps5mBpPCkFFNCdIP+2Q4fTTBwHmrljIDoNv6hK4F1y+K
5EqQTrs4bJkQrwXgbwAIhdRuusPwvvlxL11AbCXLEN+kPuoMfePOzPIKlb32pqy0
P27JJ0Nrgukl+OiUlFoBxxClkc0BHlcd/xssKJezWhbIoO+tdTwpFIdyGni4Ugca
CsslEPw9J1Q8mrGwzQjEf42dmqgsWh0IhQc3EW4SHF3qvgIt2C2305r3Rt3R5fBI
S2HQS+1LLpqC25vUZ139SKbgkagR3mjl2uiZp3jcIr0T+7ApwZtufNsAKc7JdAlB
/RJ2PgQ/UTb8YNyY7/stXlhZIL+BZALCHbhfEMLes72AWGUbYVd4fdpbNehMSALa
3oqKXjtcW1VGSuXjFA8RaRe6ys5QcMETzxCpxxn0DKGNnA5u+cJW+ZDYJv8DD5TG
+nSCZU2RhiiyhDpikmnJz4aVaVSjy4M3pcMWyT1QXpeehDY1BZeCmQjv5JgyR/Zr
YMsNfZxgb4XneQcshPDxES56g7t/KbcCOtY3taQuAZBgac3Ow0i9a2zv/QFCWNGU
ZQcVOI7mXu53WDVoP70lXQhhZ6mzgifYqKY5BjVF2cgjjlFRnppboGX0kQXCdpv1
QYbbqouZafwdQovonWOrt/rG2lYU2T6cx8ovGzNS8322UriJXidSjlrX532XESPX
pMrd/c3PCNBefiMvP5RzKcY/klCWQlEtaXxTEKWuOz1H8Zztb5nVnTRQf1orc8Oj
XAg/AT1Xk89mpTQwcmNh7G60VhVSpAScMQC0EZPgO1q9eowlxsS6ic/gDsgxB4W3
Iz2+IgByZsKlUJx0Ldw8Hq1qETOlF+5Uy6Vg1Hz1+KNGcmykbbePJs8tMo7/3Otz
NcOT0F1mIMcFOxTIwkupY2eCmBg+/uFq0UYhFQ6OpAjJkl/3oi3nkqnV9zY79hdm
WBVd7Cg/f7ztv0GlOdB2Z+j7K2qKs6h75W7nDT8FqbdWMnMUanYxQptROgyrvebn
UQZrOnYi62261+YlTEHfZpf32VJx+3VEaw7DGy86L0iGOidJI3yPdcui78TPXGT2
aEr9ppS1eCokGQtnCRXsPejCXngrQvxQIzg0SMUyYXqSHkj+Dp4PaPpn6LPeSY9M
Zxn71lj+wFTtWg12aqhQe9W4Sg2gp0YdVCKHaVDA9biNzz90FpPZoC50/OywqSq0
9EA558hULxYebBvZe3SL3CPJZGO6iNgRXumm3kVU7ydu/lUUrUaA7N5eCrhbgJTb
vAQahS7Eq08bY/v8oUPjAaIBzuOBhEOQTvbpqlAJUQV0jsY72jfnPImBBbHprvVl
QiJgAff8lCUuHrGK4C5TFUOdIa2IMIbZl9LgC25xY4cLi/gkUm8Hjp+d2xyp13KS
v2+9OlE4dnRFeSesAxCyXZT6Ih8PpUGPornWtDFsQA6OyQ8FEAQamVGxDFTvlT/A
kWO7EvByP4YTFN0npt89z2TzV2E7ygQGH0stskFHaF/Px/s+7YoZssQw3kdkP/pa
2oykL8ZuBTJ39HThzxzbUma4arjzUYDliv0bEEbirD3fIdKTV0VLoBUcDYnnLAFv
ZGgtKO75L+PwidUyRaez15xzXzz8qE+FpBdr9xzeowjECI6hUQeBO2FihJxcyo79
a8aPzUze5lYrxQLr708PRCtdUcV0ckKlj+n33WYvQFeJVgrUSKXpLun2UUU94qEN
/HBHZaFYPVb3RtMGCXWRH/wYDWZ1oD1xSGdYinqrdKnQAL4BzNZ3JXvbkmgFmEJg
8r/UIo6Rk8bOraUMSYczT5epXC2z9FOWkeTTMygLJU9vGwaGvgvh+JQoLGW2+w+d
fqqVTQEOQxuxQ7e6BR1wHm9XhuF9SA3owTcqknAObMfBW7L/8o7LUfYQj2Aa4eZu
jqoNTfuId2gXo+hpEnuMadX4+nJNEUcWqL1huClU+MT5wbsEkt0nczogNYFRoxOR
7A9QZDeEQ1fkvcZ3i+o66NIes3hB+iwTI9rWfYBZk4e82GIbfs4zZUjAGNnmuO9h
8QLKnQj10CZtZecGK3CD2YAHIAALMzZQSMGnvDp/yqkRFootCa9ihf7Q+Ed2NHZ6
1oBTJVEBH+1t1WVvFOA0HtFV1Ow+c+aGnczsNzYqAxHGAJVcEBYDfV/+athbaK61
+5Hk3Z/9ZYu4B6lUyHkeqjt8y39j86GgF8Wap1WpuwblDaqyhWRGkS8BXa4HQ3hh
4ErrcL3cgxVIZWQ+F7kTAWX/VJqQ2YdqAbSNN73TBIu5p7GGou687BdBl6QxTUWG
tCZEH1v84W6UpQOeuLa+lwNaWEJ0PqVEYZymtdP+a5x13OQEYCvTLw0gTzDHhWdT
1PwjmX4eyMgguvxJRk8V5E5UIiuMUvU0Og8Z24p2ItoVl7JzUfOkbCFyzbI7sI2q
qC8r8q2vduomgDQHKwoybvCjZ7CEYStG0zTQ7QIoBBGI9LniZ+rDpirb30vdn/gQ
x5c9V1Tg47thu+3Piz4Cpwol7nh1XW6AtlR44LovC2Pj8os/iX5VIkBk/vV+WmDj
E8/2oUQqKC8zhXOo1w4VsEb6T5RQc43hJazhTeO9VTRPSKyjEw5K/Nfh+VSYtl8q
4KrcPh5bL7joWxqLTJ+h9sAXrt5oH5CyUgrC9CCshaO45aZkcKVDSgl0dZY4Qeam
kA51g7VvTZVyG4dyBuPnq7IaBLKF3/ZsanwOEYx70oqpkhY6yaqgABWvJUZoTuVq
qiDHDfIBA67vrkF36baF7ksARHfowhHuPChcuF4o3iMNPUDF6nQ+WWR2Qo4AxoOn
6u8vAavfx/CXerVrILQb6WGzMUbQhBTf7ICxWL9SukeZLqEglgG5kYcqa/nkQ9GU
PzmUgCuskLfZdY9LTBY59Lhk8hoZ+EyeCTzdqiga0OO2gL9PP5LnJGO6HwXMKN4p
/oaFuEig2ym2eUDRc6ufFfGmAmYqx1KWBDBs1IOPn1w8KTsVxMYsHwsT2bmApRDk
1IIfI+48WbumHwOqGb0vf8nXBHGP9QxWPzonRV1iaam1n9Vq8z9PwWZfWp1o784N
2MCE5lY02ss/W+ZA55wUga0dS1WViZqig/uhqqWZ3fdS5hJy2aE7SY4ykN1AOGLa
x7RlNFcvi4UfpXx093fEZYQwHn4eaiwClViR7/BPXIhMaavbdu6BgBXr68BAv6sY
OaDYBLe+qkvIV4ZxPc67aoSYJzzJ3cBcN5fF0UhrwogqXh4wNhHJ4HADR2Unnvms
lB9l8YU5YVmEFZTX7jDgVUgcBnp9+GXh9WzBipLDUl5sBNUoSYTtpKq5t/8XbSGh
6KpoV7wlIDVLJ7bnvArptONkRB/FcVfZV7ir8EjDlF+xY5y3RzUqiB49xJgJsX3g
bMRniKn/lt1QDvKReiv9xXYGHZ+0SpQdFQZ4QrF1Xth933c4EvC6McH+B7IzUbgC
aAfhEBB27cSZ3whqcHFO4AkM5B49Rd3WXnORZcWgaTsVTjBT6/dCduktrqkKfZtv
pmod2pkAcgGn7VOFyiYch5hBIxm3I0S8BgV61B3AlnDJC4oeIpIjTd1a8iytGiM1
2KuP3cbtsvf0RCdV1RW29T9i0HauWuHoBDWxYIVUdcR4f/zC+pwLi8++vYYvNnYm
hOtozuUhG1yzVq13lbyZcNDlllQxsdpEwWYyLhx99N/HQXrHuGztc4ySbp90BjsW
DKvLW+Wu/0F4W77dgo8+SH/TaTZUEKJx0sYVUd3aYbXDkMXwho6inIBiDs7H0jaL
QLhACdTxwpLAyoevF3G4KPk1TW+2CBS3y7yPdtOYMqf1SCb+Qvm7vumgMWa3G7TF
OO+nl06Bcv7Pjvx4HTNMiV8i5kRui++eo/mACXX2nlG4MFr02sTgrUzuxrxkHtrp
kuTza9pvFarpyfMfYDWKjN/r59xkmj10pVmU0fp/906ZCsDwNEtOqRydswhX4+h2
7gIfTIdHrqy7zZapHTJDcF9Hy68pmMl/+h8qOgFvBbeuJ3Rn3T7CT+39m8QQMCBj
WwZCys4SbTMauNX73m+muGpeVy2PIJrTIgDKYKt1BQPcQ6WjR1LPafqcrsqbSliY
pH0SDdC7J0Po9Gli302ADVlZH3aLkLIUfBdU1WO4kuoiYU56PEdb9b2pkALAwped
c51V46IgsuZSn+b+YBYB5DEzTVXwCmRw1O5hry+LKWv9UuL7dgPThA5U5Tp1Lr8Z
tJuR4Ew2vztWeqtqkhAs0d/104ToWodQAHm2evsIM8dyfEjK0wcw48HUARYPPOrw
yCXV4/D00PXKC8zUnfb11HkM3UmjzvRJmw7sSyhpXfsPNxj2YcXzsgEb19drBzYP
UxH5lIvDDaPfPsTZ0Kljx7oSaZCSHS/IHh3G002lhSciWA3UcnvvX+Hsxv4fWVhA
QmfWp1yOWGFNQsSc/N4NSZpMFmag7AKvAo82eh/XRAJqVzbyY3wNzcwhG580S8kV
IEvafHUqK5AQTuE3M56J6y4H04JGmumCosLngKVKibvURu+BHHuCHDwMR0aPXQl8
s2ry2NjAGUKsN6h+pJnmN70UWJxZWin6m7t+H4TliMMzfVtGX43xpmxImFJ0L+Fr
/jp2vCSL4mv6fYTXEYKEm9rsH68L6mkXTg5XxTKGz5UdJ/kpDTRAe4g/wHQqxOxK
EGrBamW+q9G7iAnffP0uU9vBMyGsSxtnw5emeHGNJOAwVyp83hNvH45OHq2kFYR0
TzlEGd0xa1Ms4jst2g2HpbAL2rV02dtxaiw4l4AzznNP/EJE1VcpktUJ7UFs7WXI
InoQ6A+BKrypGFGS3ILEuU9+vpz51Y/Gl8nZeHr44/47Pm37JUiDi47Z7XWkyQln
Am4FaWtYdjCACk8seG2D06aKTaFverCONb6aF7KC0Mi+TdGv4wL6rQbowv0MN6Pt
3x55+mLgZig22HuRLHjEB4uSGPvTB4l4JNbLdcOvR4ckrKd+XBEhj6AMzRvLyO89
w/Z9H0cq8nLv6P5wCeYBN1bvKF+0cn4DZzgTVdDWdBlxw2o6HGqDhyZNCvZ2W5Qf
MSBZzY7X4vbobPnY49EohpS5+d5wClfgiJldr/AWgffueyFdv+mbbAC+GSEN6C1Z
kuegdnfLqOcIQRZCRtXRzdq0VjVNu60Tf0ZoubVPuzVZIvVXPMTgumgT6mtcHBh5
QTA7EnYBDpUuFGc+1gIgtGIMoS7egsc7Avo7LdHJ1h7BdCXq0ahIK6/7bw6SN3dd
E5w8YVHvjOI9+G0WH4hW9ZXy4Ae6OkXKLePKnKqds7N4SPzMYEoRcfKhUZ1qX6rv
OlKPTlZNsh/VmmR+sphJmlFZRc1WwYqW1RSx6WdJoZ6ytHj3l9/6Auh/FIGNJrBv
0N+1rHH0KrQov7unAGkkBQzn4beDoHFVYk95UQ00T7mkzDv3rFG5X5arzdL5QDuz
rLStVcN8o6j9TQI9uzHhoJg4+RW0/dRuV/dAtJ2EWJYNcd5qn4MioG/cbAUdYBUi
gcbsusGSuVFzQDz50U1qTdOWsdJb6AxtRwgFIeSAPL1OAZa1TFN3L3xjS3HeA/8J
bqelnL8YuMvDyhhiwE9iq0/AB7Ju89WJsj5XNSFBgzXUryCJEd3SsEzY0GI4IPdJ
irL8yLRvJPDwERoswIhz5QoWHrr4Od0+jave/KYFvPlWIy02+Qbz2X/VnLw1mJXN
YQb+50URgw5oQT/JgRmMa0XEe4yHDlUkRDkGEEZJWrFLOfiA9Suyqjmig1ZalADc
8zYIKP2sLdQvwsDE5umeQPYLxz6jrzoDiiyEsIcnxJv3JeSc2En4nbUH73afkwKL
rug30foNuqc8iwDvzOqXmqh2zTe98wuMGCRnrBQuEs9Ier+WK9DI01tQU9qFjyQ7
CYb7ONfSQ6A6eLJl0b9gK7h2dgBUWSWBR0uBJU4BRgbRScNehKYS+Xyk2phiG4n7
4GpmYLtmwQKk/UU0Slh3HnH+VRMcfUQ7wqjUtKT2lHb04CMhMaDbVjLvk1TYr5s/
50COvZIfpWfpmORDuN1KLSKueXj+QzQlzCTp9YulN5CGjJzblno4XIKFJ/gLROWt
poYDyC74XK+GPr/yjMiCBQYOnJ15cYoIPFoafhJdZJAY0KvOT+zifm4ZgGllXphN
pZtCjSe5EetAwh6OfD1h2JuvlX7t4GGSgEgjzBqnSW77DZkEapgmOW9rCxRlHd8i
mLeV07ZMfCNenbTgYsoaHaziZxW68lIJZlck89Kg/Sv4LCuGqsl6tS9cJAbeZ3Sn
qxNJnu2AWIBMuued4y4vu5ZAnO4kKBBYc/TfL+JuzmFSsTuX9mVK54ypYPBj2srA
LAX9xCAAxOFb5sT7kDzSMXVHKuHT2Os4kQJ4+5o1HajS9weKU9bo6tMMaTB1GLPI
CuDWKKaIi/SuCXzmf+U6CYOqjKoMTGhho26qW40f5NjQ/DwfYd+AiGNtJ9Mhrhw3
KZb+qEvs2mMEoqy1xFEUjTIevtGtwFr0JkRGQERwQxvP9d/PxePElPCgYXz30bgV
hXTt7ZBJ7T7X+SLdkZW5Ao4FMqqr6iJO5ljkevQzZqZeCJLJdka+71MNpusZx7eN
JddFhVQ2eskt7bZldYwjzrrCs8+BEKYIqz7fbzkQWx88E5l6uySn7UvSEeQgGZwV
7tsRTGREgTL3ZcBum4gGO7E5wVIlzVqRlXGDyl/bMpRFeOJQligGAmr9zOhCRcvl
Bo7MOgfki563H2hh+VSLn3PXiHxZHeEbJGR/1uotJ245kqQCQ4paHAI66fXzjXSn
HsPz62z3PG/+s5RJFdhHaAqPcTzxnJfkN3E+SsVW7j8Ylk9I1UX45T3kJ6GsRpLn
u5ueBLePqk1ybaMv4gFPCxvpfkTvF8/OOLVhXQnba29wP1uX0U904WuW2RDAJ8gy
wukbTIhFsvKy5MQGW4LrNgNNe7MI9aYbmiOU1bZ5QTBN4O0gt+9zWMBbk9YfLnNY
BGpdr80hci0tUcSI9w+o0GL43Z5JjM4Z5myuvcK1ElbRSBazCAqOMb49wUykt0ej
HdQo3S2LKNbqCcPfGPHiF0SvjVKdr1fNPb6nPQOGaBgJ5+oWbXdc8m0WMgVrWXz1
BScoIsJ4Bye2T42RqOnMUoiaUwVuDGGWXfD+5+0GNuBekvDrCdKHW2ElIqLd2jhP
LaI99Fdn+N0gYoncwP4tzhDGGiFh/Cy+VE/TLN8uu5wrAv96GhV6UfBelM8tGVVq
9UkaJTXkO4e/UhBX8wNJpFK2cMbU4o5qKu3MRU1wR7lerafg275QqPydQU1yI+zj
8KjWjwWfPik4yKkYdZUdPDnK4o7ejGtadxcbNaubzwykLuABvVBdtyK2HDsdnJzA
x8n2U0VQJANpWHSLax0OYVP12poPFNzhHyfydRDu0OQt6r2WxYybfN7bYrRYurDO
2KdEiouN3K6hy5UGO4i7F0midCnVg72ZK4zC3NSHhDnX1DdYyTzOchQ7NjzsA5JP
kTIVJXOMtlfF9Wvb1VxlHcJLS7P3iA4VwP3h7zWEqjyj1nJVvM4OWej5lfZKzOh2
dSbMtVLad+SYjPqPJaKUyLFuj9QIrYWhQewmx771asHOsBQ0LouzWnpCEVPZfFqV
waO6LLGzIN4rh+HXXt02L47qeazvdKnT444tcWbArfjyuJFPuZyiIJaR9KUxYCQp
+K9RY4PgDFeiYpaRHMGDKwjwhKqO+In4GuRbRxOvTRDatzMIm3jujjwUPUSbQOTk
+5WxOl1AhIQNRngxJGC/9N9eiWmo4Gf8MIRwp3FdUJsfhVkliA/kffsFUe9v0WDW
sFobgU+1AyC+/iy7/FD9z8VcI6EO/JXM6sIUhCLu+caMAPL9R6e7L1P0qmb0sl6C
AT4G+y5Fl9KqDwOofCgkWLhr+7nIltnyFW0ha+D8aIEzJ3ZX3m2VD5f7zBluRYTV
sLCOsk9+Tq5WJKTeIiyf4kb6FTCrmbB1mPH3CrqcLuO/Ov+m/bvui5WGS//tTbuV
CWwswYtgu3atmMlNGn5I/2velAUlesjUjsaSKe6Gx89Scl13Ynh8tMrR3q7dgGen
If3AdQ1ocDAfiehVGBynnJPmOBLrDqNDot4SO8m2P7ulSjnlru6WTnEs7jQm/kOW
41M6vBZPmSTAkMfIaFQQq3brd/R9XAHIw6RGRO2rFyr0XjxtgznieYyhVHOvnZwI
9OYt47zt1UT1SbOed1Y4EJtAl9VFfty0MbMmxU8d5HArOEu/iIJ2VmZgXkxYRkIx
d/+II19RcFuHdZ0TVShNUWAi+ifcceYNYsUNj6z6zjU+pfI/K8dkFk8J5sj0gWeA
vP5Cz4izImisa8vEkLNO4hsvFnW2LmoEDioXxbu/A6DSK/ZpHqculmFY8kN15uIl
O93m1yynqzyAw44MnfrW9qOVSrp16FS+r2TJWO9+7KPCjtixp+/NC/X6RFEF2i96
FOH1bNhhBaXI5IVRY0+gL2wRume/UlBeaifoQrHJ9UuTXLhlgChHeAu1/SMlkAHT
N0nAG4+43Yo9wX4arqhDeqME3ocOiwRfUjle0tFLSo48HlNmbdLV3xviFg6j1d3b
CmZn4ZFWw/zSf2JO5gU5DmGAkK1JApX5ShcthuPN4gQv5S/uULx2bZ4WgBPOOQ0b
gKZabtkmtYfbKjaQCifrj6QABhZOya2Eb5s0lHJK/ENf+00tvfwRSyeSz8wxVPZa
IDxmppMGQDP3eGpNhB+Q2wABTPl0UrmCV1gIT5kfqrHH8lxZwv3dq/AviqMCJyVz
2NaTu1qQLN2drzvHj5lUaRj+nGk+HhmmwimmWPYTR5fSfBx6dwL1g2dk0y52+Rkz
GMpM780kKcYGp9pGW3LxwkkeXnil4FmkK132XTP2zzIm4M24Z+445nkcv9r9Uvco
/FPA4shVLFs7g0bPypcnF11ha6S1fn0HnHrDtAFRKsvudL3L2IW8OpyN8qiq248S
TG34TnWZwXCb7J6AJ85uH/Qm9AOmgL22qP0kGSiQlAQpYiE6tpl6D+VqjFr6Zulv
HqFb280rQKb38OX25WNSi08vWsugDsL3V94mjZ3bdu+mYmJXZ4YJGO8gz7ramxaE
o8MeFRjJobqG4gl5Ik0xroz/a0X9OYUr7tEYuvMRSVgdjpm/9E6i/veVJAhgX6/d
22EEn0c/PYKrHyGRNrlNjgHScY2bWp95Ybs4XtIiH5ZP9e3ZH+hiZJHRMlVTYU+a
UCqWaokGqG189Xg6tDKI1SsfAoieBTUqvAnjH4UBjdieI4uFDQ3/+GRc9O0Ehh6l
SGGdxxBTkXbTdq9eGdXjDd/QJlL4XjjvCDeBFaxi2u/DBz4rLVnno6IwSmFey6jU
WLdWAVb92lHYFmHfQ55xhytXYD4ckpGouo8s6OPIlMeP6Ntc2CrHg3qnvQnQ8tQR
pJiKtDnv44fTvSAjGewV7SByoCem0uadBnX5I3qgXxnDb927I7j8/G9e13F4RbCh
O0YjIXZUIP67hUdk2uMND1FiRPVFi3Vfvb4LPbqKzFnIW2xvGfFcAW9NMWOWpxSP
EkmT5/VX9WlqIVI815+axPbUClw4BbZQiGXo4X1pFDEtM0lJHF1h4hnfBBTvg5v9
ciHDjihalJ41wXJRsD9NVRRFykKAyN8q0XOBJ0TaJso+6ovdsFO+HDDq8s7y+w7E
9Zf/GXwOiWXhtpaH5KJPsalGLkzEweq07efmYTHtZbjwCGroWJCCIXuynL2cAU+W
R/Fo/qsMBtyeFSOIExq74Fy+kGclk6KSdPIl4tipJkAS9p2bi1aZZLPJkW1J8NDY
085XRjgiaAmDmmoa6MPNmcfYzK/oPRNJAHIXlhZaz7Q0mtG4bLSuwuieaDYVVGrr
3xgbHR4JHVX7xhcBXr5HB1zIYKsyZASK4+lkauIwYfVo0juXVOk7nqhpYltwmjjk
HfCqZfTBOTnOC5MyIueGVR0tQ5YWnCB34iTNOuukdpeeW1MyO3UT7Ta1t8CY/3cB
vm/e27SOry0JbV6ZEnduLXNhFzypXRAJwqdbAQl+c8mJrjkVGbkzzysSYBEKzfwy
aaKkquwB4yH6Au+e/TUTG6UPA/0iY3CejKxtEHshrYZ0ow5yZ02jEBM3CvfCK3yw
5yHVwlzmpKqCmOpOI2rhPmT4znsZX+QnA3wjUXhfH7AxMViiPBXC6d8Bl6imRvsL
4uYarnqbykou8fbAfDUg31iOkkJwnVDy7YJDt3aMQ2NL6MqD1KKloJoVA9MVIjHC
bILYgbDhrpB/+lwjPCK0nY/2JJvhK3ygBMsjQlBh6LzTyxhS5dGLsOINBtLvd6hY
HJGAqfRD3OvkFfAzsCbuagCACu9G3FdS0eW4EmQeepDj8ovwdzNp6Q4EHkXAZxfk
MTWRvsrOSp3WZtW/rYq3AR2PNYFp/yr/RX/fei5K9CQlPy8qL5Z2P7XhYidS5cxX
8l/VKNOrtNo0IGlIKGEZu0IGeGtyw3Oe7Bb5PZOQXD4KfGqx1AvciwOlo3MEYCxd
FMKzEIOoHs02P9iM7hqj7FAYBqv0ChJm99YUeQPazejrqII8euGRQVQHS3dF7uTX
Xw5FYne4zDaNQl1ojaAO0jF6HLeqVlymj9lwCACtMBHefNb/nKWoKZoF1I8pykLk
tWyXKWqj8Bxqsv7yYeQNb1JEkfBEKY5JV8cdCpudqR9ds1a4IbbUZOJACA71rJCI
hcIfpg2M9Vskf/s4BzFJjkbfS0u+6izjxRPUqCkm1TjYu7MSvke90bRKXBv1b/d+
ADl11pKEgYUBqSAlwuzCwgSLwBn0yojEIpnMn0e4OTRoGqW+srONOa3/zvtHXkvM
4mcbIBF94oNjVm7fKQpdZrU+zHcadPK2y7cZQfBD/EnmHjaNW9CoSXlz8TF0YugS
tuGGwhaLEtnAfE8M5KvHHLpgQP2SnhEML7lWjziGqZFN9ooTXO+Hj2wZ1Z2qBfz3
167FcAtdd3ZNgZ/BvRPHtgpASCueOGz6Fs+cjKb33429Y4VYFJ9u983iUpKI1/xh
/o8dgQ52exR63P4q3C4M5WllG/5ScGLtOqNl0ZZ8UF+BdYR3MlWDrylg5jMu5l4L
WmolkHwzfVGDdnX3Mvo1jyk5VQkOi9TzKDyiWFzXv2nJl1RoKMUR+xmcR4u8jQ54
2rRzXC4IFSP6z9NMdf4gJeNEQw2usw2+oThjJVf90VJWbY2Sk6qBfmX2GxjSjO2s
Z0Js+PpptbZQ1DizNIgr9tLwl6MWeBiOgFduwlNFT7QkmELjmgKzADqypkygLhIG
d7Tkk1oqS5E1zDlLRIOX6enNsXM003vBItQIun7gyRKNfoqWsFKJ44bqVPqWeSIS
OawzqweWWiC4Io8q5MztZbO9EnjzVae+axUpGau5gwVTixbou7P3lYUvgUC8nk8k
bWmvxYgFEEaKQ4plnaxg/H9nFmW5Z2dcy/Y6cCifgVZNkYG5aM9QKP8p1+4ljrk7
EUMkQhuWAiM+NE+lf19XEHMeDSYbl+9wiRLxwkdgZoMBt2/dCVgmVng4h+NZN+I4
fwtf9y74t2g1mJzKyoV4YVa538qNNQ4eag06g9d/WX0+eiRUT37uDcMHrGz66xJC
ClF3NbGHZk9dMX6Qzbub3GjyJntbq7vWJntEJ7JD0e14kZww1BYCtCXVrtb5M0+v
gSV3j9RVtxRPNavkKf9DyauoBtm9rvbwCLLROU6oLBCVYA1oyQZILIVngWE9iobd
ZX9WCFGA0puHM4btQuRq2rCX7m4XjSygHWzJCvHv4fQ8Dy1JWGfz2A1MhJYQ2Bot
GIvaVLRdSgBdeXIuOX5mCL7+SjeHizk/SR19dTZjLmfVyx00pHKR7ST63Yql69sB
Qt8CwX+wk00mSsuQznteStIwXwhcsgc8gFOh5MVVfJmDXB1+3zsvgVCvOu6UeL4N
wrLmrqR21p8U7v1BDwLNT5T2fAKhHZe6uXHeWQrv0Gx/lLgWUi5v6gMO/0MAsgWj
xyGVLnylLgM5dMQd7poONemF0i/nYGDO5Sw9qpeKRQUs2w98+Ki56ws4z1dxY1aj
FWJ18WzK/77mf9UkMjzJ821NP+t+492UBjtvhlWAaLhE9pc8eayVTJD6jTJ8BP2A
ukWgJqPr/ZztIxe2M1N6piq5K8aawtQpw7g0X3p3drIsxtAuVNwier5qyP1Q69P4
E/Iq5dkbMcqawJU0v2jCQrlk9itesWUeliLCwNrvqkmU0l51VoT3sY0g/tpOnf4z
eU95A+o5BTTyj+nj5CY+9pWRC0DmsUq8pu9UvaVDOsdUBR2c5IOk/KcAjx5he5Rg
XWOgriI34uPJ6Of3ZaX/hj8YYEzDEaPNiL5FWdnNe7o26gbAtb/Wu5mBVCKII4/v
KZ3VbOCOjZ9PaFgPJvdsCllWYOhTuF6/pP7jlAJRcLCIFaUHZcfhF3prs4QG3eCz
lMArpZhyKEFp4OKQtA0F7Irb/XmtqNgye53EtoYCq4eYZ3FjyxkNg+dXHGaJLx+K
9A52JWcXL8tv46/0TUjTWzZEySqZm0x+JFzvjee41Jsw+BYVB2RmSWmodeM//SB1
UZ564un4qTQAPqjW5Uap2iGeksFWMbhQidu82jhQijxeI5GFAd1wvEJm1J9KGjIR
V/WJU0CjOl/o1CcmOQE4+Spduc3U8fzyj7pXSO45LuNJcRVrXtENSve+SPYI/pP4
cVb9VqTi0Ut/7P2K6WatklGyrcahwWwbHvc0Uq2bVz34sgOhGNbb8w/CbPB04WIE
za9HDub8+WcrqLDQyJE6PBgoKLZDdW36ynXu6XeVvzfntrEbdtg0pFfc7DWBuLtM
uOTbxwXkTdSqDVGpnF/rTYOzFKkkzFWP4gTUyP1O6s4fHoU5yEllFLs80tHRy81R
6jW3Mtpn+Oi0UvhkKqADJzCYQ7yKVDymlVdIhLlxnXpVvzw+HUVj+J7Y68rVcNpZ
96per2lczbM52EG2pBPZuQeHxBfqwlmM4ui+N64b5WgyTQdpw0tSic5Lux2ZRMxR
TNj1R0vMJYdEY8Drh/u9P+9YYnR2SShciA+NeZbl/K2Xcd40j+vKnmXVN/kMju3q
WotlM+tCPE+ySHUQv+jWxbaELiXb3nl+5st1WLYu2TFPlGUeCHjJHmNMxZlwb1rC
x+PK4rRIWmpT4I0qALxFAeEWLc14Q/noDJsrdP98m3Q5N/y+Q8C5ysjdJHT4DR7+
p20RXPQAP+CvcTpiLcL7pZtXAHrjt28Kjvrcc0LQ5d1z3E4KQ1ACVHOzPCSpjTW/
Kwdp9KBlpBkIITFeW5Yt3GAAhUhuAa4AgORyFB6+Mp0WMjQLRlCK6UlLxicjElHy
1bl5gZ4DIvtjQTuos0XlbWY6MbazBYy1j+xIl0DG2uVBr6tIn8FYvfcQrDrwUXfG
T9Etlzomyp6BBtpG9ZX98k/R3Eewniy96xHTju8ITQr0Rj+nopsEU7tv5+HpV+Cx
GjiKT3ODzxG+j7VKDc6meOoG7DXY0UNOnMGoNpVwOHy/p7//9j+mTn0xSI6AdJkK
vKKdslXxmzO8WMSgJPhwfa00Iatpi+P/2VqN9elrUQeKtYShYf5/K3XSuVurlNBU
zC5nJLnMol7a+r1wvyWNB+dS87skNcfMi4sKGS8JIoKuudP+5WrDM3taawWzTfX5
1hQiHlyK0e3KzT0IEhfNjp6BC8l1eQsbroDlPepC+zMEy+rQC2m4tUvLL8XG5kJk
tZNALkNjVRkGrRuHNOyBDiPzxTmCIHsVnpzJZ4BuMHIOgpMxOWMAM1aaElmD+qEz
eGkyRit2V9L32DGK0pwkuWAigFseBym8M6sbu1u22V/Elkwx+x6tTN0fpCyR42LX
1yJL4V+jSaD1D/r/5NhPKFcin0zZYIpo9TvpZLmINePpNOwt0uvjp8+yJsjQDFpZ
7QArAVd64r4cGJlqV+Zciw0nOBLHObU3TAwFlqNcGd7Pk8jguh0AScWHU1p0wHKi
BBQY/3dA45mPIz5WRCtvKqYZMrOxWkzgncGO4ejtUDKQ3kdg3ffhd0XeJheqMiiQ
9khOtf/GLJiwXNxh51tEIElNKE6EPP12bdBbjKmPTD2rFTjifreSuVJiP2zJBNax
QQs06yCGSTh2d32+bf5Q3tO2vQEfRhhEi+9LCCJgInOC+Ir4pFXwfY1dHaIWhiHC
VvqlMmcM47UGrZ5acNipJMagbYUrJ+DeYh4YyAvZzlo9RjZOhiGby1dYEN2j1FTm
15nold7Bxk8a+jMlDEMQ3fHGtaWNAt9IJB7jR612ThMBVRg/XhfyYTIOR/jcaOIF
SIVLRcu63OmsBBywVEaGrnxln5hMqRaXvCmfHzVy1PauImA82moNXDtD7VtXErK6
2X6tZZGDbPOPXe68qqOCRcMULQsVf8rm/zGZfu6ItTk8Og9AQMt+ngxSNMSkH234
vzTt49ozngTNbP7IIztKeLsBMsNhBO0ASny7pBAgLCaFjLPIiFHEWX7FtIiEOE1k
LeQL2KLkfkLjfR07yCW04C3RkEbD4JsCuJEd4NVXamlNXxp2gnv5c571iuKTL64d
AbjbsQZkINYicijgz9eYa82tl61Hsd1LtHEqapisHjSpa78PX6pHaiQyo6qjSJrJ
sFQfjDJXWoAh3C3MNowGr5vZZYYcism2WQu7skaGsUL2vPHX/s8NWNQKpQx4sXN/
ERY7MfhNoixnZTkMvVdb6wtELKEmjE5PW8ENnV4IjJBaZnely0ZDSFtSU7lgndkI
3HgpKnhtAnysyylE0/Pd3oavYsjw8sdumlKagH/iACbcQNH0iJh8tDLNB8MuIBZp
E9qJRrSpIgoHDLJbusfJ3nXCksHs24oMwM7KPALkq5X8JivIK6dx0i8tB4TjCS3n
9/JPL0QRlMkbkZElPaLYZVbkjNXmCqnqnc7TAns2FOeGz/amYzf2KNFoDYs6UD9g
TB02DxayfOnLNwqzPWJJ9TZCaqQjfmZS1v6/TRyF3frEdF2ybp6F0o+H7Ok4gn1X
7pzKmymj5B+OKCBHZ2LIwSgdWtfWsztEFfviGAZxcHWTCQ4ob7NUh4Q6/PmnCENf
IwLbhAdZ9NaX05fVVFH3JVPVheL1QM1tVHiSmu4S5722SwJQ9AZ15oAOxBG7v5Ik
BHwFrlxNQb9Gu1e7AjUIhoXL1UxTfWKigtQKSust3T8NNza1H/XUW2rEpl5upJxV
kGAHcpcxl69fiBQF7QpH4/5jA6HExTkeTusDzT1TJ3BZtY/H+4vvhtIUTQuyjd6f
I8SB1j+WWplzO9zu+0nczsvtD4tqhe/AzdavSuMbEA4lZdwUZ3bDABQuA4zSGot3
zpbTvIbdDXh5eKR1VTL6mgrwXUi2hVD3tY+wROG++iwzzuD/xaG2wOB3gDZEX8pg
/G6ltaisxQBYQ4Y4hLOgevb9YvbaDWhdDhNn/bhxHJxucvG+6lUE0q6HL2p7b4f1
3OL0vkXI04IjsNo+U1nr8DBqKpNKW9Mj9k7CCWWCQ0M2quKqWzM/by+4ZHsfEeX6
62kHk1Hx2kzxczAXzoNApy/ZRJ9iYycbuAPJAjsca60BUBLVa5jp/U61U2RtKRIF
m0IprGOyE15U0fNiDou5BHfexOO11OcfNeJVUr3pNHu5q+z6/YE/Q2Ugrq9o2Lwi
UTTmUoTMHZRYjS+hg2G8WqZeaqIUXMxClRpQ1s5K4q2Ad2eXGd0l/LWExT6C+Rn/
o1wAGdrUp2Ynpci3NZqZcj8yeuu1UkJ46o5x3Ho2bCceNPFv5bLyuCh82OLEHABN
qC8OYmhyq868mjkf8LHVLV7rtifPGFVVnarUWfVSoyPXd11comMlbgMakAGVc8yA
U8j0Zh8C/seoIiiyi8bsI3+L2I/lssACBxnsi/a5UwP+0QFoP49D5zlMepYk0DP+
IZCfsuZhh1A2reax086g9/6UCus7OQ1Tz/msVXC0OP3y0uC2niNK5SWA9oK5OfkB
FGCKMyEdnHQ1cyq/IQo7t+AmCAv8UzjgpOljwURSr4EIJ5BrfMEhFwcbFflU3xCz
cvzcBkNuSSHVM9uW6i6euA==
`protect end_protected