`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1E9zWyekqR6gJIEqoyePTeigwKwItOKg5Yr0rj/Xb/KN
NqLEezaf4d+DCVXhQkBpFfScZmRppd22VWzSl9I1tx2o8e0EX5yw2MBFtCCkx7Ma
KK6yKD6OkVxSJj2YWMIRj1yn+kM1ifpzJ3mgPDSvnhjDwjFBU7sJoqcKGRs9o/w7
7ICfuxlTb1dsi/hcINBfDcoAfrgOVozJQdxl0pY1dwka07EQ9UhZ2dR6SRBv4bM9
im3zEAr4MeYacvpdsBC0MlgVAYNNpvTi5Pq5VqrSGpEKbDVYKJBOhTPSUGuu6FIY
WHddtpdPBnNWJFyDlHnU6AIDIFaueOLrMmprsHMdBDcHPmeFo29dLhdHprz0Gukk
zfGB++5J04C3nWgYtU6JAwZ46qWhzosMiSRCiM4liH03tk/WrnoLHG1099Hh1Omx
n/9fxV9brkDA+ikHEb5D1l3ncqQtzaAr0JoZGDbvBjOpc8RClrHQM8rVUJy4xauo
xzkboZKznW6OKaAGdC2+7omg2cJE7PcDsfdwIgxEuDTUKxdsqf9zYI257Mfyy2FA
0WuynrUFRY9H8uUaBDs3FgeDa6NZYCbsN2krqPAfViC91YR0rNxiUe2wjAmCPRpb
+cajABjQZeCRVfIsovmOfjA/OLH38/3mmiFScSMRHW5zucRUZJ6xTCqNcRHTr9RC
TeaTtLMlONS8MuJDLwl1KVGDN3qh/Qd9UoWj4pxbuUv+YEBZwB1Zizvkuoalhte9
X7v9/FwSVZB4blPd/qArFBRneqCNRThwn7plReiH32l7zAQQmqJeLsi8jO3dHDQb
C5vdaWaamI/h3hm35aURU0sSxXucDRmkr+bJh0oGu0IBXte7cXx7tgHSu+UGUevT
tTj+ZtR2whrEh0C/DutWFVS2c2HK1Yx5o9BWHz/8USOg+JNJNl6NeJfVu12M/4uN
4UQY7RPB339Ntbf17oyunJxCbBtW5UqC/Vi92Za5XUUkp7YEvrvL6YBSvH9A8HMK
qumZkIQ5pKL8Aw3VaUzTEyl/oZXAck5JYEkTnVtl73AHRe8DeZeQMY+iDSy57VQz
csB1SsgxCa9bpdT5XF0L63Rav7YYjB4WrZxjfZFWJdCGZm0SKAiocStjkxBiZMuE
FmUioHJGJEux2+2coqS+rnnP48TrhxDvnQLus4bQdevjEXWiKUN5+tpjT7175UCJ
KuP+SgwCxmbwvWIEtXPSaKW/lWkREnx5k3tFnjZY7TaPCNNf9h7iz/XlmqgsjHOp
ajs3BN2L5ryRsdQPH/jI2vDpTM2C2RnAYC2hX97FuvKl3MFPcPPv4DGgHpA6LVsQ
aMIVC5MjnwjrVadTh1s3lthazPBzriXPKRWJYevYEpZ8DEYZ7hio9b1y7R0YtKzB
3no/WRP4RaQezwbclSy9EYmaruXakN9q6N9kpO/5Flq/FaJwf3qprebr5GPQHo8F
y9Q8+qXYtPH6KTOZN9ri7ES4F3/lAenZxo4mCOshCOokjgfsSdoOUSBpSQNyvdk4
/2w9iHNGuFhx9R8DtoY8KvRUvEU+kvlzvqPCSy6FGCy0TmBHYOLPbe59T/qaNT1o
Vi9g3D2hevV15c3W/on3qGFoyMhdyiCvFHFNj+3rPUCkdBSh23uFP23nu6VE1+Xy
ipGxpfBmYbExDVwmwRUwHwX7cbV4ho8Li8QbQfA+rgwEElG154O+8pnhxvA1Wjzg
lBaOo5YjBBcrdCRW8DxCXTHH23eeC2VOcWtvJF4+lSshSbpX67IhtL+VrbvNcp44
Kq7h7FY8ABpEHixnBQY3NQivwh4yHxYwPbYJ4rsqWZI0dOev0tBlSTAOUWJOEjNT
DFK0ieTX3DOtXhTLAlMzSjykcLYT9Y6z/PJNMYEuPY09q6rsKrZIB7PtJFBG3vpi
GdXMacz+Ri9rWNr6tOUI6cLKV0DafkjTlzmiXUfpAyYlvW2YVpThX9Vh490fgBOZ
gPS0gSne9B3OEcxBlCD4ZmnnA+R1vei8Q31TMmjQgsv2qHyRecFZQ+S3WJCy+tiH
2zMznirGAvNTu0S12XdjqllyU+Z9dUy99iPX0vrW6pexvGNkd55YegGC/AkwHDx0
WhhDCDeNbt+zaXmV2QaGNStEpu7d/wOYdsgV6orLL4DstuQN8jY9B+TljKqk1kRu
a2yusXI/1FqE+RxeRJfecgm2mHaFqjKG0rB8cRF0RQf+diZFIjrZe7fxfy1yjfSN
VA2fOOVb0Xy6YUGYAPR14GbaJKfkflHGXxuOlfn3aIO8h2iBQIXvP53BO577cgzz
lO3QmydAXcgG7AsIgOY7J+6zMrOgpeD4fsUcaAwLg0aMi9VA6Db6fGEY7GFnExkA
1H2ohXztqalWUfwXOO/KACZDHO7ZOVKl0B/txEs4lgl+qUcHE1YF4hCislHjuhiy
ptROBDDZzgdCPsSZqd3HWIB2J67UjD0KtWSKqoCdrbpRQnHUvcJogoJP/8GCgMDN
Cz6Ek6TQg0q0fQVxI7psYBcVofb2EWmlTs87+QKjPLl4IPKVJSBPyhjoRfasZbdR
DWigFtdCCLJZuXgEobRWu6E9SP9T1jZ8k9tk1zNQue7allYAmGuVxlIA7XU8QJtA
oLFGmvLF9otnO+JHnjCeFU+Bwmy5lZOpVvPpzLOe+ZfoLIV4TO9KGlGXMr4nRWG5
MVY4BPvY/Og2Z84bQSNj9fqo4/H4ZKyM/2LyccZerLO4V4L7eH8c186zyB17FOVw
gx4W2bUCTYxnpsYEmD96TmyO0i9NWM+axarOnipB3RmZWEs0J7eEoqvaGU3m0+6M
pCz72JAe8YvmZ4lFkY7u6a9p6Lumo20Gu2t1XkhXPJpDTS2KUORIidwcA2iFLio4
gABiVjrbP7B6zMBb+ZnQ0N+Br+fdv9Vq51ni+dd8WEU4LilHXNV2c6yLagV71Z/N
GtpZuH245fp8147oEwYLGL3nylhP9ajbuwBU/yX+NQjnykIUzcM/dIy8Fn4v3Xii
Sa1QoH9Cx+jr6j7canJ3xL2aDt5BqrO+zjMww7xBjniIposWiV/j0B/+Ui3tyc3c
qgLtY2M2rbcWAPQ8c9gqsTR7AOyVfg4vS1jAG/lJb+3ymz1iV8MnvSyeNypFirGs
+Q7rpNrtpbbTlrhFbXOHV7CVFz7gvU4s/G3dD8jdDWv1tIHSvOeZPhDqXz+iEjed
YWrRxfodcKFE6wWxvvf7PauKZrKYdcL6r2RPgasI2iDtmg+i4WbNiWZHAHQIcHIw
qUACTE+vAKhwTMaqQEMwRXCqnqTst5Hjgwua8nAauCoq7gqFGzNdAJY8LuA1jFXW
DdUnb0CNB+43NwMGy8YNdmpOFr+XFC0PXaJ2Mup5EKrUJCBPCa9Z4JEPyWLM3JB4
6+F3kjszhHl5vai7wC8L+Ho2GNkwSpyujM0mvWCEY9J8o5RU9CELx7pEoxlfjhMj
3Bt3bJR7XthLhdeOPilYBGStNMlOHAuZPmgx7dFDeAzu3dvkRuKRjG7RzumR2078
I+tSAFzQ01SbL2DqhET1zlCIFDtXv681p6bVS1j/9W4OMHse9ClWqS0B5WR4WVFb
hRk001PxWNkPAtbT8z3J6fd0uJhUQ1FCTtkRy9mUoL/wHsm0eGf5a+wc3i68C2+8
wPXGoBBJXIKQ2xo5XnLl70zhyQGUHo7plPrW47RuYM/8iNQzKjjCIfF6ILhwrar5
n6aojDqS5lEH4YFjdj7ECq7GoADoluPEnLuobGMsG1gl32EXZfBDE6eZVzi5QlNE
jCeO0CPY0qA6WZkjCJltpBVMy3OsPHH5QiXLvTg2DunKEeB88JwJFux1otTvAA2y
JEbdMlHYC1OMdz8Yz9ESTBpc/7g0XAAhtt9++HbIGwVa4kyLBJzWCjN3Ux1K06xp
PJTQSB6fEvxjw6TOjxNgpwUsUyw2nTWrbXDzZxQO7EZ1QTu4rVXAwyikuO0zUNPu
2zVUEpmkA0EJXbJtsPrpbepZAvW4zF0OTR6UZ/13Xv94nqIFfCEhcPKqzWsWLBMs
QrrR3uW8d+pAVGygn7RWgHTzm2iQtGRgeZwBW4C5vrN6PsPo1WvTGrLBh4y0e1vt
nEtIx9wbUOI0kCF+Xhsik20K2KPkr88TlVJH4gh4vC7arJAJNGSzKyD0349Myl4t
PiXeUYMe3/WxXaGLTvA81dblhQSm4Ma+9YN1ALaDY4JW2mPWcN12xznd3IKwPDl6
OUe3yYn4YA68TluJJgDXCcZNuHLMuLqZ59x/XIldsKH370NHSsz0i2iEap8Xz1bX
+fvjjDX1KfqMnh9JdSRSGH+h/9fczvgDJZP/hU5aRhCONXbu3qxk2ZLKcp+5OSy2
KceRNZ+4PLfUi5EjQPTGH5UhuB0UFHhdq7Ne8Va0k8LJQdsrrX7na+sFrRn1whb7
uRaB6rN4KTTQQizQPZhS1z6WjIFK0NtGcikHGL335soPmgy7tBTvC/ldZIY3O9mF
nJcGo94CmfOApxnQQkB1PXx1xy6zHYxFR0Ywe9h92xgsoVV4BVW7KXg0YsyTSvf9
gRos34jf3XSoCpFqYaJRLLlfpk8tjztmp6ddEGvX5vNVUPZrcuvYZjWo1jSUV8m7
C50J3NQ8jW5mZ2rMlo/0U2ffltbRBDUtJ3qHDYp4Cpw7AAbuQ5I+0xaSJqcwTnun
Jk5BELkuvV3Zc0Mfe/1YnQsDbZuUDXj1tqYBlRvyXcTURETWGhDYSnfwutLriJiE
xp0G5cpHr5WsZQote/nr5qnCNJtKMjOT2dCX+JpqpoMbK5lb/YnO4hFkPaXXGXQF
iPvRfTZ+Ls+OMdRu5kc5yHsTjqjChUgwYXzCXKf2temt0blCXijNbAA5hJiHkeQt
WFORbr/36qDyDY1lN9II6zv6y5wfvv59Ns779znnfocr48oDIYAXCEs/r76as4CE
XUTvt6c1UWG+dnwKXt4RXc/yqduLk1EDIfm+3WBsmHBbFFxQ1pL32clKsTYaDNoq
wMqUqo2sLvBIY0atsj8Q+PNjQo/R5UB7X6N4qPFx/FSGmWFF00PsBxJWpaCoXCQ5
tdjxUR1DiIVwd3mOMe2DnL5IXuTfbAQNqKswM3OT/DLkZ8G3hKueCk7n59skdJFj
mXBkPAt8hZQli1kPNoWxAs195KvU+GjU9F5p1lQUWcNxXM/DscB+DJ1Hu5iAe7//
at50o/YbdSudsQso0W5ZsBMv9v1MeLHhuNO84XqeeQ5QfjntOwXo+p1ZroUc59B4
hVAqAnYb24PwAgi18PFJsXniA4yBaqPeIUjRRsz6zx6+jAo8OqatDKS7C7+YNJ7V
Txyc2UFVF7DBkpD5zoOLfvkIpoURueX9fhpnW5YzfwuHfEco/PJ7Hsy9qUOopHmu
KGiMBDbNIgZ+SDZ6KlLW+vO5ZJyCNovXGgGkvDviCb3Br7+CmpHhiXEeKbOlg1F2
aSBC0LNI+BimIvlYR7J3XFQDLDf7/kOtnVDclCnP/6YODvAH3uqYSUbx+GRhk2Np
OzUpmzc7LxuByTWCd+kpAXtbDtEVLnx2lIBE7Q+BwEF7e2LsmR0cbEaSu+xuYXJ/
i8EIQxvCpqO4oz5n5bN4v1bJLAPhX7G2a5P8O04qf8BgbwdXZ0aV8CcvXRiID3YV
eA8vk15T4bRo639x74bVKzszRzriH95r/IrXJKqFfVfoAsYGbrLqVWHYZ1MLGPf1
1GsoViajTaIuO0fYTgh1yoQtsuKrCbYFWrRg4y3uXASJ3NUM9ONtxI+D2AWxLbzk
m81ZdLAnY14ut339K+3sJIl+1vTUaHrclc4/B0N5X4WyCNAJwsbaKHaZOaGyMU5n
xOx5li8kGDHyjYYuvB6fFN8zT3ugFMHIjpVPIXdj6bHzKyBwOASVDbyfnRl95iDS
jPDvbT9uVW6SzH0ZqwCp5UqhCF1//d//fpbkNYbeTwUKCAj2YISnFbXAvl9DCLbv
Yz8bI3cHRKKo3ROiS+AvMf2PwJLQkBCKGrQM3qomSCcv5sS6nS7iL7qRqqbL6jd9
WSp4jg+SAjQWBpn5hWZ226gaKTNkm9DRxDMVaR+pdV+1tTTXGHoeTHVEBmxe/uUQ
3glF1ZzNGoAT2hJDxSAhJkp0aQnuEHVPled01a8rOGhpXU3U9YwTOnMv+2XKZPOI
IQSUB0dT/ptiIPo1wVrCH2HzPaDNYajSn0rrMa8SGz13hekiUOVAVAP6A/cKjaU5
40gUSjEQwgVTUUtHENMEspMaheh8DiIZvxPg1/0dWu/ShNsU3CTxoeOcdnHW/sqn
MzE/qYoYj/Q5GYSrWyOS+Mc6G6EEvSjAwjM8Ib4iwfa5eQ6MRsEyDn35fDmWYWqr
AD86wEWtLvGlYy/ex6bStJLcG2owpyLjNe/iGJ/flRdGbcRVsZ6XQIKrFLyPhpF1
tlYOSn7kKSBrJXcaDjyHTkCNqrvhYzvXYNKQl/4qcocG64dvuzNb1gkUkJrDdIwt
ULIR5QM0ZrKNTkXHIAJEcNqs2HAuOT26qcDmSaCgg7wQaIoJMJpUEH5/QnWOFA01
KfZmQ8YhbrNOyrsp/C0b4dB6Ot31c6xjClcJTERNd43VyTyMcnbx9G9P/TET9DiX
sMm79m2SmTL629Ksdb/1fmdZtNkIRi3c8rO/DeHI9aKYJIgO+SGZee7unruvgGof
EkqY5bEkXfEAMdO62P2ASE8Y82bmBj8Qbrez201DA6ESaoxdJ+NL0p/3UgtDtrDA
yTUqqOaH91oPKSsM79WPAxqQyzlDDc8KRJq/PVtm3MgkDb1lgO0EzojONJ/1I4jZ
E3RG6E0peFIDYB+7wh2h3nZXh5PIWTPzg2C5repHwTtIS5FBB8YMIp0q2DSpwPw7
3Wj6SZwLqNKItsv+kPuyWesEqPN+Pt/fua3VtY0KqOYjxQgTNDgqtYn29wyQtto4
eZBQ3F9UPEiIBTwI9in3y9zSX9ADX0f60wpFIR/yWGlpBwDoucr823Tn07z2Ok08
sKEnDr9J+ePSeXrMFwQs3dTCSU9IshGby5ekYVjAxFiTNN3hjlaFzJIz2CgXzlCV
K/3TLvWDCZnFdGwqGEAPIiQ3Mh8U79FfPsx50h4/nf3Njfdw7qFK0Xf2iCSiaZaG
NCIBIXPy9XTiqj+JtutV0phM1ygTiQvkeUYHAUBnFplcBawc3/9K4BQko3F5tDyg
7YAd6zHtk3QldNi2obNsSMoCDAorObxIgk1P/yHxoyD1szZsh/XMZEwGioCkx7h/
5SAsJDYEZtQC7IkVIBoO2isLvl1fLwteY7ywzStZ32/ggCaPabsFKC4wqUK0cSxK
CFRGTIyqV7t6LXG/Z6htzTEdjTgpeSMwuze8i1Y9BlpovUN1HB1fLAVK1a08bxGa
hhlAcPV53JI+c5BRICnDWfFUOY9kgtA0k19YSLl2FnpPpVXbJ2qm97Ztm3lq3dUP
J7sAbmwmgdDYJxalEqV5jmBU/74BJHDPpnuboVK569mQecrO8HmRIVhBxqn9X1lW
FxXFRAyMWz60VdqFrv9vI2aUVM+6fBYmXqljwptvNr2QFP7yMEgVc9eDI1mmXaCX
YppXhh+lveapmI0DdLao3RV1foNAqyuAzWH6eUaKlftj5tI6z42o/XrIvVMA05yX
MXTdilx5m0mRlmm7p6wYVYeT5QNt9F4g6hrfgq+m8RRmMKvWlFkV8EpH/p5u3zWy
na9fTuF3p1AT6vsIvLSx6Xo8wwO/4AmE4Wp0DM4IqM/h+XRsecJhpfNptuUd3g0l
CeOsn2zcqV0xAUpvRh9Ynwv6fceWTjI4Z0hOWuIFGBCRuiJyZjqbgXJJ9FcyIneS
D8tewb0eU2f8o9J7t5Gy36maYA5h0TH1tjrM2x2Wd4YP0RbKTvfULQvdrYo3Acvh
j4bxR7cDXhFFm/URg/RwOFBkwWzv+2ktN45OaaTAxenz2PWlW5ERKLV4P28L3Gx6
H8vfjMWltEQA5skN9ZMlFBXDe4rfMqB30C24kJboPH264QcUEEKzxJTF4S1od1HH
53HTgb/VU9egPWT680LaAuHq2IPh2q7dJV02mq3WYh4fWdffJb14Ywnzus+9VPR8
s8Q4Wr3hAXrjKCLo/GB1G6gTJXrBWVZ+giISOtUwwcpeNDvv7nSipQ3lqI5TO9/U
AxgycSkLVdOx5C3Ls3w7XDjAKYRO5X4XnqSanL++vz1KYXeayKIVqtbZjQl6ICyr
fvxSVvMcT54iHTfOy9HXD1bPvyPdrfjn1WrJEhdxDQMiCwXa1VQjLT1+TPmij8HV
Z5vf6mxBHmhPQ9g8fub/5Z0VTt6w5xyEaSVFBHh7zSi32geRqOiAT54Es1zapE5F
aTGEbF11UFcS0nH+Yn3YrqgF9MoPVEe+0CPb1QtDFxWtu01pgaSDhCrQCdjnie14
txHAWqn4SP74i9+CnPoF/bIWlWuIzselqM3v6j/BuDeJrWvGWg6UuPt0OpGzxjPh
Zk12B3WV0gD8juiamdA0q4HioIC7JBiq5olXtnP4lkj4eQmYGbY2ByJcZTkl+Y60
7iLaEIApVg3TXcnvZ1BPJcxWqTFWeWMJ17bqcyIkjyPQqrBrwCZ2S5nIq77GPM5q
15IbU1Zr2L5rnNwC+Lj/Ad1cfO9gQkISmB7gr6GyQnr0TRvlQgLLl9lFBI7Rp0Jk
DNkYNzOF98jNQVLkPP4tFc0WxYYbeK8DYRjKCiLXA91yRFNwPnWAXBkYH3ViO9yP
3HlF/OTXcZTK+4dVnqTLRzOW/KbPDIb1HHP+kNevrqoErbMZW3a8dxJrT6IZ4YXc
inGJ+Cm+YMezsZ08zgCKLVJl3IY2N2StBs0yZ2ppVIPBThsfGZ2Lbyd5XoNx4xml
jZnlTI5XmRhCgPbW/0OzxgzSpmWpVp0uYTMezkdywKkJyhT9yj8tYkgsit7UCajW
YEui1+IIR+rxYONGM+BJagun7zGfiKqAMONWAm73Txhqp8w218dfd2TGnRWtNJGt
ElgBG4loacWI2eiLFKwLv28n+rbJit7i8zdZlzx9cu7yBnFVQagIO0pavP2iUTyj
319E2Jr+V3KrKfJ0nPBqSKRcIa96BXFMwIEsGUDghcZiGS5O982zvbrR7Ec20BdX
JVYKYgm6itAdxDjeMfewNg6ykfVP/SRxE9D68F7Mft8dUeRuZ/gR8qLiyowe0YXx
VFeftk0zKtGeOrXvlWJmdXnikVQ+5CrPuV+2XbZzz0DJ4nQ7wKl8lrU5tZZued/I
vpToHLHHAJJDMvyiTZH1CX6qKxWQNFHhGCJyAhcdLORHiMhREwVBi5Uphmab6H8y
epxs+fBs0rEsooGw/H14OeTU2vMPjUSBgsVvHd4KrngsfwNzxHR4A82i80M1o9Lj
C5JuEA6BAfpRP22W3kYGD1/CQmcZ47cPSC1llFQacHUpm6I5SVzHbAEkCSllGLsa
eUZD0l6hr4OAuBH9yL3xZrKmBWioUG592AB2rf9W8IghmdQLHmCn+krIpfmVmm/Z
WWG99tmOGOHXActjOwd93KqwBZHcID/4fWGP97KOJg1LmBHwURAlO864afKHNrfr
BJ9BxYGTADQKdYJakNNrMteSnAAYcEqIo8nNcEkSNpwkigqKMNVklnFcqzb3OEWH
QRcZQWKVd+3//yZPb7gyCYSwEQkFkdaQ1NjcmDpdWq2kucmPW7c+Pyy1GLc3ua5q
VKJiIP+6/xfEKfiXTJ64uBY/zcIMzTLfw3YJFHuBJGDRxJUaj9thV1grsOdC+MZC
CqBzBIPvonBarb08f51iDJU8fA1N3y2abKc+L57rndG//PPUz7ojDlDJf9UWiifb
GIiLMX4GLnfE8wuEWTG7y/yuw4upFdv24TAfSP1UiA0ENz0eJW1KjKTxAiIuOLna
7szKQ/TILsKjszKFk+OcdtiuJBk9joj5cWkjQ5KMfPKkAK1tREGN/Ch2Z8PY95uS
se9YKocNrFRYm9E6cgRmU9fwZwFykGda/rCHRqq6TCUcfaF1Ec861i/mk9CBxSHE
1su/1gV5KvIfW3/u6LB6cp12HQU2mc0w/K+a9sSgOGqjk+9ePSlymw+0s2C/S45L
5AIpUcb+pZF0Wtm6UEaCfOA7llF0PHgfeUu6T0PwyhkFiaSredy6unuWEWlygIFX
KeL1dxslGNIX8y43q/qkrCOpXfc2dAmuSbW5WRLt3EZ9nFoziCyIL57D0TIieGVo
M90I4U/3jshQvz0kCfdflJA3Ae/q1VChfTjthZKRWRRg1I3i5u2ImBejr0/KrGsv
l1pOFvl/0n1eeVIZ+ymqBUQB37ifANNWZkxYpL8BPNGIgMfzlK7GXTlYwlCSaXix
OM/Px4yVdwDkmROZJnwEl1eCz/IYdGDm6nQP22B6snsupLaiqR/HF/RmlWkKH9jt
JX56jCujDWJgFmo5HcrJNB8z+nQMbpg5Xwj5TNMMhhsz51ipfoQHhw42rxtrGz+W
FD50yx6Lk7adH2XyNh+Lei6YZMk04vW/+G+X2DSbN25ciY3HMypOTT/3W/vJ0IWS
ziglceCDqrsSpyXZT+rnVmUwc0YPzTN8ethQw0Dol3sIr5dpoeOjHpsC6GJ+x6pW
letzlnfCc2q7+yLVFvyxM/xA+6jmV9ukJlgqlACrpzwPEhfEEWb9xEcxEAEkQl+A
Nzsjj13/I39suc1zLU7+SGZgpb1JpDy5z4JMK74IOzRcOoaEq6RtaDeGpo7LkC5C
f8GMA4AJXQEQ6iRplwDVwnId2g33GrMc7uvl9wN9hF0E/Y9c8hflzWNyj430TsOa
c65pRfCP/nVn0HuyP2ToXbRGACoE9NG6emWa59mmbYWW+4vQadUUyVegn2YQ0Mjt
Zc4HWw1dnQy0dKJ8YO0Fu1n0ZIqbT2HhlAum5fysgP+WcXJz49J4fpOlSHSJh5Qh
4uEKCQJMSXK3p2wdcNTZQrQcsZLx7lBPYAMh00MErzBaApSHzU6WnqJPh3yDDPiS
+8xoVEi5/lw2HNZSiPh1Svu/2cfHKlGFp/TEw+crfxS98MrzlcPzzW7Qy+eFnWNl
3iNx1JV8xpM3fYx9fnleNzLg3aU/MMQIloUPRUI0uZLV04YX7fzhBCUNRuA8O1BU
D5wnMGo7jz+UFSdi9xG471YPQZ/RMrnx5wrVYQ0dU2Z1TyafuOmySC7wFFVmsjFI
t4lebJc+0/GfM04yPbgvW2QcLDhpjpZZErD6jS6uVwFXSNbUeDHSUSRjfoD8qdef
QRQdXJwGXAknB9mSdLsErlmZkK0P8pG1aL+N53+DCOBE9w65KXB+qhXsFd90XiWC
hmtgyK51MJdMDZJl8ZG05L+i3t8MST6Lk80O9coJbb5eoAn0FUst+J5vaVbAdECn
F6d/IEmj8YiPMYFSgqZ6M04LH5VuKeCrQwzxBvPiOHeCwCitx63syznTVeqBTNdo
rcndJywzLjCOYJZPlM5qDzrRu1jeaqQX6BbGsESC6gDs6k8zrPIvKOHCu0VO5jhY
95ZuG/+7E1BLPxP6Ryc/VQarsPZdSvAHvmosNzFPASgUFTq0YW/CbJGhba5kwRgc
FPTGJ1+ZKE359D5UmGK5eg67uqaocmW5NJhhkJjF8rJLR84QwXatq/vxJsVCY6Oz
INZZo1lw2dPxxseDatKcn2iv9Fs/o6SJX7BVWEsLxCgRRU9HrqDt++gEN2X0azlJ
Vq4IgLm6Va2B1d0fNwBdDYDAkwpgwEVQvf27s3UYyzNYl2+czKYf0UCgD6gDh+42
2POHMmIwxrWU0sH4U0MmFb86PWR43Xs/QzxNPv4J0qM+bICkKZZJ6/EZQIHFPR80
RZZuVoUept+hU6Aest0vreeppXGzgqZrRjRRHVZip1SjD5Yru6rzTavFqVBSi3aT
oRsFefL1cczX43DPYWZQ7VlBu1xTGE2T9fVN2mw8IShGgw0UN4RjGPEpUWFuyTis
aSoNeFjND3XLSVOpiARcwJUZSZMkWb5mgNdInibqexc=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
vWaiee8LnCgatAmbQJm76NJlinhaHK78YZ/3NkMUV9jy5LuKOPZEhtbifJNyQBoN
84yCdPG8UkyfCiVzwHg+r5iv5crhWIgek9NvmRdr9yvIJwqMyAN2r82QiLU8E/wM
Mikq9/27TKbweopqSKQltYrxOv/V1L+4iVVAODhSsA8XvfRWigkeRikHl04OV1lv
/vQ+ZDYGwOmxiOXPE6JdJrqAI6+g9E9OErSCAv4/mLfr+yCneg4cmdpPPWX9A8fs
Srz5SUb/0P7vDyVyrcuCzq6uQf1apBdaIO5sp7SUqm8nVVz5GeR2j7EeFgY6QTHP
OrkCSWXlg4qGPzJFy/nI91msrM6b4qQS//OgRvIFS6T5c0MzQqMj3Jde4VrnRFhX
5UC0SaozRt4MekC/oe5zkUJSBk/tf8ubQzrO3WP6MGs6ppj0eQixV5/tNw9mF/IL
XBBriqyhbz5BFZbnRLjj9ILrPUcO19AMMtdNS8+uj9XWeCL0RMF3MaK0+a9/pjrD
6hbMkPzlzh2qYXxiwUD10Ny1y4ySPZY0LnMSx5aXPP+7QI5mShayMMD+U6wj5vD7
j1DpC1j258liLMemipAk2iQ2GA/OqN42YUOs55eRVDtWobZoV8KYnpKZLrBQglIj
SiGuhUwsrHG4Iw+q0qrc6Fu42RkATMJS6PtPnBf/e2Om3ZrvPRirHuNkOSum67xe
xommeqJSR13F21eQF3yjtWkBuS+xG3HyI+f3js1YELe6wXY50TbYhUb5mmK/Uu1M
nd4R7BxmHkzxSYHXKD10uB8cyx3TYnBwOnn/ZWqXAHsn4ArnRPZqV6px8VNIrLFp
7BFaDCtYuOUx6AdD6vKQSY/G2NNTa6QTLWnSkJVSSo9pwLIY7TWFWM2MsQxUfsum
3OhiCe//znuj9G6pTEFkzlROO7aHBFxJV/uA+M8mi0IteW3PhTUeqRPol+TzfFl5
6she/0dingDHh+teu4rgVJdqAz66Ll8XmjBFPV1SA8CcRHSVIw/nt/qJYEe93BYP
4dCOohI9N8TlAhY/Sl/nCI9w3dCXH2i0zf3nqRl/g+rOqZoqzC+/NQdeDnQF3bIU
p51WWNipVw/eSlVEVn+6Voq31MbVIy5WUjeTbisNAYMClJI+ngTugirnGY7P4StB
jrUEJs3qgeKoy6gURFuuK28PAOuZWtIlW1VPsxERpExV5v+qjYuQJDmeUPy0pdm5
1GMv6hEYvE2OIJEZ3zioCaqf3xX/SlFhKzFvajWHkl+i9Ppv/hdm20U4uZkH8NKB
Wqt4Il4q7U38cq94972wrHQjLuubSBLRCvtU71zV24JV1DfTvZbbIXuERpJMBgNL
pxat+lYI90lQtJeYnJKgIfh9eW1XIQZn8ToxBLaSmcXfihT1pcGyUTpEDOnQZfsf
Ngg6KFmQUKIIxvMVAKz4akk7vjY7ZnCPHvSlkWwTiaUuN7z9jMTpXgDVjOsGf1ON
kGwcZgZOQUXdpiKSKMBV0+KJjQBdkuNlfg08JronczTiyNyZRjkICeCEhTYOEvzF
g1WATYV6dIA+DMjTy6maaCtCYOnm2lX2OXyqRlGfAgh6FKMyfdM/73XDqjPgYICg
DWg0rFM9c7a4t82glXXsVyKNZ62yMfshqEl/hRXaLOhWyoU8Gpn4MkOvD55ihyh8
whImSsY4+km6Rw2kpVYur0u5j4Mox/MBYQGYjVi0KTFJMhB4769+t4VHTC08sSNg
PRcfyluwDDRG0o4BONV3Hl+Z5BwU/d+Y44ON6pY9AHiu/pwPJscJ9bQhNTvZ2Wsa
+LNR+3oYJMSf4a+1x0ZJ1zw8EQ+rT8wZQATddd6itM1vNq+eZ8//vY2jCtGhrnPD
rl8zLRQ3NYzXWhoXaIsgp+xJskCtuDPO+OACeo6xTeS+BqsGw7t+F0CpK7MPaD/A
KsYSps2UcPAKGkuVOpeMfGhH7DDhtUKQpvMAxKK91C3a6OfkGEr02wO+frTeG5OS
bTlqWEUFalNojs+amyaLXGATJYxTN+q+Fp/LMpemjxj0JPn5Y2uFav/llUbQQlZN
YH8dBLKlD8Ai3nAccPHY+KM8/FE3YgJ+UN/3mVCNZIyS9i0KrdmGGe4T0j+RtEVQ
7xR7oHv2kwPSzR7W6qpQ79uM/sza1YLwS9u2r04i6Ps9GOqw/0IBRZaRuSjyQ5vK
1k1o2OIu/VksQ1jx5CnauXsGykKnRVZBMqDDHLRrpLxatmXupDX4o7c+0l8KEwxS
sS8noX/GaoedTy7XS7YOSzG7wd3xbaFQIQzoo/M2iPnQRuuJtF3opbpHPUdL4f57
WNp1Guijv55z8umdHUqtAqH/CyleyRfEMNANVr6/Nnb0FFDmyKeUBHomx2nCdmP7
PmTXYa6O4+37TRKMWTcUHOJPfYna0qaMCjdb8xccxHtiB46nZRusjrMNFZe0eDzo
oWp8Htjl+LH7waCZoiu1vWBzyN54ziTcxCCiimZsuOVY+15cv/6FCfpetx8za14l
i2fOIAJV56lQrBfNesRZfLrvrh7wV/UGt2/jgN3htbT6cTXwqRJiP0uV3fYQMcKo
pw5zYO/a8sQ2lPa9VmxFriKZDK97WxtuYlGojBbhRwFwWnYJub+lN4oK/y5eAcda
Zkmi1AnFm+Cwcv1gpKrnwix00g1TcHU7ykINA2tphEWtTC5Xi16HYoZjF1emt+1E
L26PspcjGexMoetqWkIBaaDhqLR7NAeyCUpAYLsPWpFpU2489h5REG5EscjaRd+3
EyYkOXgQTXvYSOrAvPI8gwlJUCKsqFwJJsTgitMGlArSKKELlo5BV1BbE04VylWq
8uuYEYtQSQC0WNJ+qzfI0Ef+KQW9P9pH3PthcMcleXOjYHlXtt2BgXF9WJl1gxBm
nwADoO+Mw85mOGPxltAJPEESTu2Or4l/pvnjIWnR5WBArgmxDMcZXtcyIvMV0Nd/
ZgiXgoepwrov93jfLTsEdOAt7btM8AftjaY50Lk/E21ypQ5Ap7xdBCs+60xrKp2S
Z/HTesCTCAl3DOIYcPM8rEXxEagwQgt4q+UTtakh2c7Q4c8lZNpcpXi3a8x9IFjY
WAx3wwUq7fLV+7c5zhsb0awwk2JX0jLH1gtekDvJ1VcAlkfv3EaH1pi5HGzz45Ss
jVweExTuY4pd1ggM2ME0zsQF8jXRvkA3PQcG6SVC7Rnng41vFFogXneR1GOul5Jr
r7c7QEVMmF/8Q4QTJnNqYQEyv8K9LALwIgnInNRwWDTcsIwfM+q48vSNRzwcilcQ
HY9wPpI9Rcv2ticwAwQVUjr53URPzUFqnnos8DVFvMEMH9QK5unqlXT/Zbe47PKj
6lmpOCx2k3Cn0e/lzKzghW9Jj9u/1dfP4n8OnZfLUG6+0XUu8fohlgjFOQRSTp0l
P6fe78wGXOSuVUmH+X7O4a7zxbAP8T4VPTDSxRTC9b7vDNVE+vSq9WRnTxEkARnR
QYjKhoA1tlkLiCkWjBWff5h2YmhLfg6aqtz89hOKZfdzQrOfrLdUsUITwUbJ3LsB
7nb42tmOFJ7nVu7Q2vM9Q+qyta9+mlZkgl4tE4EHDeqi+ccxdNVIC6CgGCDNdI6v
v5YQ6fwr5zuH+QKJhCanT8IdS/LRsrGKmmGa6E3qX3Z6PEzYwoa1DSOT/dBL0KxX
v3Xycg8BGZS/HDkW2LTiTIDTuhZd4kcm7eZxfxZMPU4gd9vZTcbtFZaHLVwjtbvL
juwhhfvyrVdjp9ZS597T+V1mi7yVweRJ/XqjMLoTdX43gZh11tHB9ugt2iHQ7rN2
40NTayujhJknDdC8HV0y+ehfDluK/BoAMdMoZYHV7cbi0TX4hp3VtCpltrpD1y7B
ztSBnQ64omvZjDZMbgkdItKFaozGgw8gCsvwgvRbxPGTQmnp1LM4KzS10Rf38zRD
DbcLOJNvCa8SfTEL1oQAP+QOIgve2MLJsFoe+BtZi3dhl43aaNrXkT92OXYqElKZ
CWlYUY8P+MWCNWOFM8mB7LJ0NDuQiZ8qZKwvejdp9+MXGkRHGdiAN7sgFKWe8gZc
dWRy/Auw5ZRdS7JzhoErT9FMCvS9zUqt4mmCRoWBL+eTS/3PKVhEmvWUHvcsrFli
2fHHFT4tY9JZv0bZnVAY5d1K/i5oO0rqS8n6vd/HuQ4pRTPJBhou9bFzHhUsUuyC
ycupFArn+EYc8t8hfkbPMwT6Ytu7X3oSMRA6eir2TT2Ez93SSieztYnQf7RG5NHB
c2XUTMfMTgr9ksWRm/Yt1EFPFSu3JVsopZvipzFBBI6VRUwxdctDQa8OUvqbWEit
yi9YjRPuO/l4/fcr/Yag3yVkxtjJ7MfuyxV6feNVcGAr+hRq0ewOuWN8nDcRxY+h
b4G4kFi0JLMv5xiLdb/IU47S4do1stixT2diVHXebbdeStGqAwAp4zOkmzEZTKiY
YCggCXlSi+KdqNuxG1Ki/ERrSaAdQrHwZLLhyBUT8nVPT3z9ZlByWTofWScjpKVf
ZO6WZyo/qPGkmhwYUWg5mUAVeiBhCJHyXZWxFdJ899nu/qPUd/5jEF7Fb2xYMTka
IahVkCn7xT/UZyhSX6abYVb+ljgQ3cvzQlpLHKgao4Yza1L7yN/HzFcrnQAJERvR
JbLZcA3ZbnVJswYz2RrVbTxiRRsVchSPFcVgVhmmCAAIlmLfq5LqucaMSfuXYys0
rYNa6L0AQV8sowgMIBF5ueEQpBjBpwl4DG9KvkBP0QSnAFlN4tKSB/3ZGy38BZlO
sPGb7ki/KH99nE4TPMz04ThNF1B5CmXjbFxcRqAbhdMg8CQIcSYdCxAnoxjXAE6F
DDSLjEIMNK+nB+o3175AkC2EiXjm8MhHUkyeUwHmuXwMvXHRdd6irlBsdhZuQ1aE
6fiQTico0R4sOtxUpfrmGKFKgfGylXQTxDZ5UeeyyJPnOeYjb+egMkMZv/M8heZw
cq6RoWMxoAoBs3QPoY+3LD8xiDHe89hPMlZxKTbINaY+TV2kNkbgb8S0HE6X3BW/
Ojg15Ath2CebZ7vNS2z32emmThybXlio3mWnMTAtFZrGwEYqK0lDEZO5zFgS5Vut
p0GKFWxiZ17Xzi73aCpIHsrMa6XYQDHbOgEtjnqm86PlpawGh8ZnU2ViF0gKus6L
orBLkSIVOYGSXrGN+6qGtYf9U4D5LEwh9r21LPud0O1Q/Dpgf5ro56j8bzCBR2HJ
2N7Rf9CF28QwZ8acIehYn9AcxS+PevLjospC/vTHuzDkD8j0znjWcEhEm/YeVKA5
dxw6A17JJvMyYXykVg0QjSpkERLx7rbDyFXBOjFOBv+eeiwcxGJ4uzD9dJh0fsah
/uHrYsPcab6fMmZVPWRWxH3SURyRfvkY8ysq5elHqbgNofKNtkUFfEaR7pa8nqBz
WelrMMvLopVXyXKctSpq69hsIeEElbbAWRfxFuK0oWoJgaEAb2bPF3jhBLXx7zu3
g2UCJz/HJm9TbNFpWJS/nZCiwJDSgDSal6I13KtJ48+xgz3wbLf4UkKtig0IIS9M
P4qtuKw5QizZMOcZ4aSWacdhxE3B5q3FZd1LFgSBzbJEgEjm/ECjRTnAyUviMJvs
OeyEklv3zQ3GeOJg7Cch3BmF3q1uf8IXaJoGFz9V/dGF1+BliF4CsRDvfqLnvdMk
ZUiLwoAonn+zRguiwLrzVdmwdJD2cY1uBqSS7bjmt5+t4479xmdTAYpGk84l7Dyo
RGJikucXdnT7JQBJZbZycYZS1sqO9ELFazd8YvmS79TWqfHkha3H7QLEYtWYQeCd
x/ZhuPm51puEWyFYOh6rgmhbm9pIGqbAj87mLPAG7w/1SKAaxO3fCSKQAT2foU9B
cFozMVrvAnQG6StSsUmuURczsw3LS8IqvbPQVd6G93LLe2DM+APfueutkNsvQMiK
vamb/vvsl16VTz3DLB9142vzOMVKFv2vP31CjlByLpFyjV9QxDnl3zA+eWCzVVVZ
+D/F29ngQEDhHbICJP36nB6fDeZ8nEq5XdoKp9Dqv/44STI1NlQ6FWtNdtK8hCJV
6va50mSa3Fq1UOgD9yAGIhZ7dZl55JBmMegqEIVNg3xGcUKA57cgSCr6vsMqqxUt
7r2ymMooLFG3Zgq9CPIoZE1fJuqAg87j7hCyTtalLhEWFPk808ygtnor9HC5W3IS
ybjiyabzbM8H1FiqtU6UNNpeMl9dX96tApp4m9J5OIuVcbWGKzR4g0Qag//i5Gpy
MspTbWvfpzfKL/re8ckMqp25gHehkAcUsBvHKg6Wdi5U/RReorpREnGINlK9Xzlz
ngPutsa1AIHEr61DRfAjayHZcUnnBRlb7JXfVQ+ldz2r4YSOCssNNviUC7Ll4FBa
1kukEUJN+n9sNfCrOhA+GjZYYeccwraZpTbT5+u+kzFAzEmxWGuO+5d1QzJQ2t8g
RH6wEEAc34QT/xhz4CNq+7WxDusaq06m/YqU6R42H/4MOPNdtur7M3QghLKRCSXZ
y3obtPaUU5F184GKIHDcrPUkIkWTWHuRfarqjN5r9rl7cmsbfdLLeWJzBYBrnCtZ
0zw9WgEREjCHuBBGAvHAT0Cjl+w4/nM7TvyVGgPjHZZSGbbtFM8Y4uDcCDH0fIg8
fUEASgMmzZ7EA+vPZT12CxE4AorD5d2EvxUZEXSfx+VfZ5kRnU8uL6v/hwPA5MIZ
fiGjI5giGreGzZZamUw6ZCg6gNd4UeTQUEePN2G9SL/f+BMUXJv3ORTvPwpqtCmD
pZSfmAESiSiFHYPr2M5r9CXNzhs42HdOEEGi8TgLev8yBLdDOHC18MyBW4Mg3/NC
67We3645wrwYKJ+ZG5pyFPHJhEmxjBtCuYk5eCTl0Hhlx2iIRXhJLbBHtbNDzIb0
pVxcIYZLZCpSOjkyb2hPTMQtj9TtZXXSOP9sHEjMljZxbiSCN8ICnSuzlM3gl19D
Qa9mHIWhIsVs+nASySkgqxIaqn652KThEMa29+PnGMp3blgHnr4UQYgwl96UAl6V
Gc6UD2cNinRQiZVOHtS35SgHKYUVkcCo5If0HxdQ9anBk9el1gKpZs68WDGqBSpF
pl/CyS2pP8FOa3uaD/mFD10VNVSqup1wnUQdzp4TTABr5cgCrTe5PWsGaXIRmK56
TuP5W3SSOdRoWuL+9EQzV4zee7bPaQ0mGjQ9H3S8oQQku8QW27IeL60Dr1ATHVgi
u2h/9WNKjLOnhAzmvQD4ulPJf/dgR4ZdXgp2f2ZsKumgnr6bk/1FXXarQbiA1xaX
twwNG2z1gU77HSMJZiuzElYJoxgyPK0U07OeNUgfbJHAb9Ptj9DUssPHhZ+RCp1f
KiCthPYlLcDHY6VF6PKBvz+EtElFv7BJpc2vX95eQ604NenmG29H8iisKvYWbBSx
uZ9bmSpIfik0fFcHQkwKyoq4lmD40mqN/uqEJmUd1s7w4Nijg8iA6SUXaoDXMynq
mR3l9H91xqgKJLVezHL0T9iEdjfBWrnQ1JEkbd4p5auqyC5/4UCt5nsAucM3XTvy
2W2UEigkL6hMO6JaaHZm2QR4hsEkakTUf8lvyCNOfBF0fON0gjN5njmGFj9XQPrI
mQ9HJzbAUeRXMnzRk8EF7Q/KNNjGAUNdWNIapu528Tx6E+lD7FVoh19TtQcntB58
y7m2ufK2P2/pcdQVq3DUOL/zgDiCAfD+sV5RFCy0ZkvKQT15laD4UV18cPzs/16d
DbPuh+BfBAdtVIbopyZzOi89XChLlQCti9b+pxwRaAtoQfHyvov5kjjnKnAR4pRY
jk12dzhRIgZcxXd6om8+YtGCmpZi1RaoN63e8wV8NcJY4Q9U8Gv/h8ud7zkjJsQU
dLM99Pj+uM/aqIg8CnSsHyKIuNLjZEIhmif6b+xU5pjv7du+WKa1WFcD92J/JGT6
yfZ4MX1HHyyXvM84sNRnnQu4qDqiseqY6G5TBvhDYqTrogAQOBEAZSqfoi7wr1tU
vMySb9Njiudhu0PcsK8Bn552KKlKSfSuPydULlYxfcT2VIZwdkMrRNyqeyuqxp8A
ISFi/euj9Xlnp5AJSqjkoc5D5nd/JaO0kFFjw45SLadxIuXxiXd3aFltGtSNcbVT
yk3EMyOSStUIi9N4y5ABfzRIy40NdpvBuUTpU0mHOv30QM1fRj7KSmCRWyMHhSGw
qE0pi3MdlXLUjPDNNO5U559RWhE+bIxrHpPLI38KRVwRcVyB+RRyxddQLSmuCZkk
py3hL64Ckq3LqwoHPDPd+M5jePqBJA45X1IkFKl3EEfduMaOTYEN6eNKQPfMVtbg
TcUGtqzdvHvzeT9kSfKX7lTF0nTYTGuRfUBDQPhAzLY84bWB106sibx0HOMupXpM
vve+E7HchgebmyyDDly/Ho/i4gGbJ04o8C/RMZERatZbzd4WE/G88obXpD9e7/FD
SPyNWaX5IElaMQSa8kqcjy25gx6hRt6pnSPL2dduC2aFdnLbm6vXFlDJC37DLOwJ
p0ZZc0aWLOJV1kLetb5EW0//CBxTvHqqrwYI/wlNeSIQTkIL7GC7/eIoSejMfXBM
sBeenhEYj2gUwyeLRYTMslwiPWaty3H5lqWKwPt1vLxLJIE1ELUV0Hco1qncMx/p
cMa3yjH7rwMS06N2eFN5Jx9h1/72+9CemkNVxDjhDSBxgDddVFjH0LacZ8KQrIdA
skleBV93/DGgQCHUqxbbMQoyS+DpXK4C+PU7HG+/p8VJ8KzNm4smGS6FRYBxm5Nk
O1XJr8eDwaLBXIhmBXXE24zNAe/5WViVONrHAZ6THWgI0kY62L+p56BgayTCgd5L
qk34G3iipvJ8FxRz6xSEtWTVZXE2q7T3rVtkbYLFWP68TDI168mM5FrZJwI8DHC1
xBNE6hmcKzJupaFhZ5O8uOb9+ptWZELMi8af+nnsWzY8Woy0yyczIYrb3Dd8VIVg
aFNzaJ88WQQJfSUt/svyMLO8LDmf/USpgYE0t39sj46+jEipZjyBz/kRBLM0Uwk9
13bXdVbvMWs5oc9/aOuCjyWcOrUpRYJ/1ltQBt55EoMd+JHnhKXFo08Qf4FBPd5I
H7tKK43jJLyZ/pQD2J+GVQtFBwKwGxTv/XD1NXMmHNTMYbsSv28RyFlaoa3gSC5h
b7oBKb8hXzusakFdFNmJ38Hu90NXg7LRXWxAh9OwiB3Ev44Q5KWA0XZNm44M4UX0
fyPvMmJ1YR1zsNxCPVTiR2qnEqh44YiwmR6SjZ76LHzrX5AbYwMmRyaa66DbwB+y
GY1AGflxpH9GJF55LEVnbdGqxqyiSXCohd0dOZVXCaMa6LH+RcrVggN03EHI5P6C
LubDNMGWHusVlg7bTw90Guj+jK3qbURhhFsSca20o4kyGoeQ7/nRErnPoS8ZMkOf
36VQjkkPK5IoKdFkr7YOgkUhK8JpqPRKTINoziy2ENGk0PXAVn0F5rPTrA7sC6E3
3YnflmlstxW42YxPI3RR99N3XTu5MGphj1m4pyMAU8lvD4iKY8abw8UKR2pKTk1n
XYz1gWsdRWR3VfKY6OdTxZj+l+KTcTyyCGXYCPTLVxHZYVOsbv7By+TUkQS6pDbN
e4qDIqLUsm0mnYAU9jZJT8BNit//abuq0G6YxH61vdstbgHOVSq8Csz4plYGV9Ed
9zvWfHl0ZKTzL4TflA7CAHUkhJ96nt1YTNwX+0wx+leapWslzZq7AC7ke+kcIe5+
tQ4AIwfZaUga6736vbe2+q3+/3k+3HfX4bfkFnhTG9yhSQy4VmCB5HIDEdt2KlTg
lVyE6EAUvIPM+kT8C3L2nXkzc0btAphyilwD/33q1iFp2XB4cSn9gN9o8O/PanQ7
L8MhNBUyvj5QrQfO94egkWqZy+lEOSxsgqXnMEHSxafivvHM1o/Ep9c0hot5qQGm
kcJ4vEA+68mXuyoifSrUgK9B85U7FEoig25wI8FJs5xyKI9Qk4so9OI32gCyhPN8
3ooYpquNFElNZZtm+jyVgfkyh7uxpx7DwTM4yhRajRb4ZQO1Id8YqV8njynqs6pr
UTUdtpvm8Glxae9mq3NKdn7FFsP8oyYRuFQRdlikXtZpoQLHScQcKZcMjWU+9GDW
HsGRzRytd/p3Y9l54GTr/KPupgxn/2i0xO/84pefu6wmIRebJ4F4DCxyVodf0h70
5dAmVtokHKezYn1kTxTx0B1d8Aj9nNuto0cX4ma35/+wOx7APP8sQPHeTP08ohUq
Txndt+XkRHtKwDYJy9wgyv1/h5TTXjh+P2LQdyPPTedx6ifzfq4oSqvLz27v1J1h
HE5EJrYmegqhKmGxvpeo0/fSZMRzHAk6HtJnpDbYYjUi1ly5fNcBCf522n8pAp8E
9vZIkWyfr6uwsbBDKlw0DWadX1dx1nA1jRfStzIx7C0t+ydiyEE+rQjKa9YuZzYE
S9HbFh1du8jHq6+SD1R/SquHhcnbqGGm/a2GmJURPBTGxqtc4EqwTDcF98EOQqWc
qQbkvIe5rZqKW9569lLNRagum0CtUhJnygso3L5+vWk7rfG19NbkRR9xf6GrSScT
99vimDLlbzzwWlnYLk+slG7bI36Rn5xdT2fIB6lw2W7KfpW3yezSo4UBdNAcsCFc
F8gRCJTFZo8Fcg6owqzadsfDzjqRic/8+nz5VnpHR2fpwiIFRP80nDfeRmdnDeKo
vIJlxCRon25K4RvtaocfcUnMPUJtwj22/j9U4Gu32RFbWe2ITR4k98uO8qWgQjvL
dKTlX1ynUjQDmydVyonxIuh9v/JtKfty6dNQalvpDV9WAE7Anl9WLBRY/C9nzKNv
CT/t4f6CrQKkDaklcEV5X6L4ADh86lSxYt8+wkpVIwDi8/0pV2/oa1jnFl6iY+Lt
Ff9BbqVbF6HrygoLEx0ZqHwWP9fu1ikcpZ9mTktru7y0JYI95h3lNWxVcILgd+Tt
9vHJvAw1Y81dx9DTP+beaZwY867srog4u733cvDSMYbV+ABpDG4+llTuDOluHD2p
7Fo6JgsBSKOPrMWCOiSzemS1VlMEpVgrE5MDbUL7PTY/ajHSUsMU4EJTNINztRkn
psqNg4fAUaNo0OgkfJeOpWBxfEdvvVFdFZuhawaS2/JPjpLZR6CcHeFTQ6YtgY2q
uhxQDQ2bflRiEVPT4rRpJTt78MEmw3qOFDeyNZZoN+2mlBBlUlS7e5ahTAD/GmMl
U0vk6eEXIA5N0Sv1zZMavqPSas/BKJNApQ+8YmZxg8q6db+afdWLKQ1juHm8RLT5
Vk7COLPn/bRzq7/1+t/vwuiqKda4v1kLgWXzu8LFVDhxqCsEVOjnPtm22urmnd5t
NTKKIvRLshnTRzDDBwG9in2iTyH7cCHXjBwiW9BydjHjLGwzkX7A1mIZtLA9M+fD
uKd4HD2cgvGoCPghn+NOCtLFbvWqe61bPc5AfijaZ+/Golv+gV7xIvuRAV9uM8R1
f2NHxvHtWX+PWGgrNli7Z1ycnRvPJEHDCpXOmUg1ClokcY4SyxtrjmUZOIInZ15i
yjQ9NlM7mbVrlxo8waXHyynL5YUXbrWx7AweWMHJswEVuXKh1Lze43JEN2PunYQ8
k7F2zU7DPYWWQlgP9PdJ//sG9fTbtuUUOviTkGaEdhcsLtXpwJAYl7LBLh9+aQQe
XzTyNaq+GEFOUPfDEp9SWgX/5TT98pL27sPpvayu2O86a7YmIWxcEnQ6BMxvcTT6
d5qoIbO3kwfP4vQnYBHdMs1i7ngvYPZYAtY24xypSlndhUj6dY3sxEYbN8Ef/cUG
vevdCb3ZfgZrK36s/mVxVI5cOfN8m3Ncl8w9+2FnXmrIp6VwtS9WOdztDIA/RnpK
N0Yu/gS/n6rmh6LeEAIBy7DIkIqWqmmf0ExAIhhD9A43effyvN2umBLdFJGpnLBB
A5CFE+wuFCCznPNe0YnaeYKbMusKcvkFuwAnq/OOeOZ2eDYE6Y4f6VcCHU6TN8oD
fQpKjhhf9yQkMH8iASRCwHEtGOrU7+SAi461oH0dl/8=
>>>>>>> main
`protect end_protected