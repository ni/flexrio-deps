`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
tZRYouEXCAgDvnyDq1Df8lNJsgp/iMufa3Cz7VXufztZBeBQFruacl+elvk8Phot
laqxoBbRcTF6yEcV3F34bDlElHDibkxl9cR/RtVi+xaRbEo3PhPbSkSMRwoFQYto
cZWEaIF4/07Gf/AMw/2jVc6GhiU9+FUeUZ5e9cT72fFejFCAkAtMdD+hJERX1KTS
xZprkkkOyROHxuMKg9pDORvsNzgCzxuV2XRA8ZVVq5Fq2T4MdCAosj0VtXjxOIFt
+DEOfUW1qDQkFBLypYuMM7YmxoUkuwhg6PUpAOwQQ9fn31i3+Tz6K8/ot2hS0rJA
3B9M7eLbIw91Rj1R4oDpbqkYSaFiaZtMABD2CWvWONDHmaQLt+w7j5vqOm/wavfI
KVF8AQzI7zvDM+K+ayzHgCsoOQq8GA+98Wb54LKd4dbvG0Z1dV2fdRFPiJzdB0+j
RjEmDT0+ft/OiJJXGeQ0hcBIC16Z34yUAELuOr6blP8u10b27YRi0FyKbERPjzLn
sGNF933KIJsYNQiVXEXsPxdy72kcOkmVg4oPTd3lFWgRG4Em2nTE5dTecJxTHCQb
TSHuHskpkuBLNviPvMRQc2gEyhP6kgMLGtozEqYvm7g38hiPppcfmFUPF2M3fasz
piWlp8/loqaKQK2Jakqx4F8yMHj2jAYAPjzFt7B/fSxzmK8BIyuHzsOnsjsUFdGb
cBLj7flMNhllyRP5D6WzbXL6Zka+lm9m7Hf2ZaHVhG0bZAFRTO10kbrd49HEtKKJ
seFNb7EjtSmz0C/z/EHbIqwBCrikm3SbXrSNoFN4YXSd687jZ08mdeieIAQRkoDc
OUllRVeXWhh7MqE2btbwqX3GS0QR4VWqTUNhEnfX9FUtur3PaJc8wuoIbk+Ab1Wc
6nMEs4xM124FASkiQdfz3fXUZ+IwFhH5bT3yVIpW9cOht0ySPIq48f9MWPIckq1Y
ap/UhEyFT/MDsZU/Y8biaQnKttz1dmRcICouuvlvqrpCMJlFIDPtO0xCHQ0o1WRC
mBdfWeeAAb01e4mkB3N3K7vYOsY3GTkVH8jAUFkBq4m+BXLRhJfsb2ClSbNpft7k
KFd//jOyvh7eKRZsDWFohjlAyxcAVRxSvqVL4lyfA668araYecQSA6g1V/iqUgcJ
vh/tPBw/DFn8PxjDEY9tm1ns5bp4+L0dfWhDr5IPdmzYobv42pL3CVRJO5vpHjxx
ynfsD5NaWynuMfLBesfqZOAWRyiKfwNVLD/mTMlOil3dyAgH4a8tYm8joUIbvA72
BbAb8Kn4lf1XVwmOX/IIr3GLmTbkswJ2d3xiq+Zq79Xlp0tvtbWxFGqH61zD63Yc
TbJmJq7PfNrLRhuSxGyeWDTlHVWENIvvXUo1VDrYzATKRYpUpUnNgL1TNBdn9czW
p66RDAKuNVm74E+HBBtYI2Seawp/y/IKq0N/o3wlBsedd5YPAVRbU7YaElD4bbqd
DlxujVxMrkCRzp3yQylpNJp7OnvUPC2zBBmvyfr0vAKM/jqSr+hqd3rGBRnp3LWd
kautQY4W8023M3xsLh/b71D5ipjmtjJUQ0n9HNC248X4vUOzydRPHFfqJ6h549vD
WpQldtdvAqClGxj6pzwBfxPp25/z5N1bhw3F4bwei/nbPzi1UkWqx5bl9xoinDkG
VenosF2L1uCsqMuX17MY3Jpym/ZAuv3Y6pILsFmWf/EZV/OTVvRhEaKM23uIdM3K
dqqC7RAUWkn4ANTxUAjh6DHLWsez5P/Mdz9W1Y9gEX84Ph/Tp9EYN/fV/rNTtT6b
aniOr1po77NAnsjT7IPbHdT1i302tb4QQm2SYu7fXXGBikm437fWPfmRbOU2rDu0
N9AH/kyZJ+KSWvssqkvYzeiIgbfFjoDfbdzvzpzraQw5lV5lEE9QH3rXHRPrvYhH
h5XRjH4M9Hvq5UkmxP3hiIJYXiNNdqAfFuKMaYNbW/VuzuaZMUKCLcH6mh1jZS0b
iWjqyPEsdHmOXz++Nv1UnSK0YDc3Bv3VE7QYyPQFB8YHFXyQbacUZOPLBj/eoexT
drN2qKfNtnCJXPOHbSjrKIgFpbjb5w4G/wy0xxa0D8HcQJAo/uUtkQjEu4bRfMrA
sdZHWIiJpGEfHsGE6jqM9XSHEKN4kclgpu9FT0GfmJLxQnfdpbK+OA72r/r6LcVm
jJ33YaNPqDS5CfIigfNNq39PNXT6dN+TimwwGATASUyY9RJQC06FdDPbjX84QLj5
p1AGr727+JeDL0jpj64+l2qdhtiIJY5NGR0feaoXLCbU5cwc3xzlYLOc76Jw6csK
tGDO1vEgN/dz3j62T9STWC6103QVFBoSBSNZt67o3LiUHf/u3q0E89BZWFGIeGms
MUZk/53rjscPzqkebaxlFgVE9IsUDVpHygluP1pSguLOnooq3yf0CnWvWulIeZcQ
lBBUex+cyR9/ypgRbvAX9wDUJORstUcEmo0UImofUvO56K5IysPoWVeJlC9qmibk
7LQ9s3vV8T2vPbdRku9yQQbZaYbxl9pu7CjbAUlv9bv1LdtKCV+7Jkd0FNbMXD1R
rwvTQy8bV66vMcccCfIXw2tjIUp3/YogtfzZ4j6SVMX3TGob7GfUe8MOlo1mnZkp
IjxAeIZ07VIJCJjsEs8tFmA9L0vHdw/zY6NZdMNkr1Ll4m0w6PPHEQesMVnlyEV0
YZ6D9L24F58ePt8pvlc7v5IE+BEKV5kl2JOFm+Te2MfHGBr7oDLZb2qpF41qSiJR
DXWk9+HZEWQUA8o+gJZTM9+ilQ+XHtegiShKIDgZOSF1Up5/k2gNYNsIajSjo52W
qiO9Fb6Vij7GdtDJcBysev7O5Uh6kcEOnobMp31LnujswkD2BjBKv5qDqWZ2eu8P
Sn5yQsVbp+UHcrlfjrqyUXFkVteqomKdKBre+wk5ZYGMe4NjuT1Bwg6eu1t19LI3
mMZSLAHeeVFzA5zAXY4CcGpeI8wFIVC60nXAi0Nopv75Yg+S/eIgWvXwc4j2Uv/Z
UUBXKSj/BXBPyK1IJbpHbcPzhdHHOyCCDBExF4TpHMQaqrabEhnLYvGfousHLuez
zqQ0glEY/i3C0mKamPel8SZ0a/tq9LwVKyGKSoVnrWk/8BEULspu0yHOX0drKq32
Br91jkm1o11fyCseZ8MFK+m2GuTNrruRVGpuC2WxY5FOoVt4ukrJuGR30z7XQVHm
tYRF4bXUE2dh+r4zOfVmVmCV9mrquyFm7cRRKAZavwuZJ8jSqg5ZIa2aBWOXQwI7
VxRRR6GhcxfcVZQZuuacAbpRNBrz8BozwJ+NxH/VoKKm8tqceFqFi7tXRchoSK44
uTwgMZ4M71nBkehLQ9u+3taBMDHTGPsWaPiMpEUYn7ci7xA+9ZT3klI4uGUdv+7D
Wc+6+ui4HJSY2BODAVjJufjpOlsYUq5FPmSZw0uy9kob7IZhG0kyu5HOJy5eoJ0I
4DJDx9iagFHiAd9Ida1tluVxOpQ250YZstm0OfvXenJEvGRMlVq8xsIvgqLaOJ3N
U6ZjQWNbmqXUb/6BKXm8W39sENBmP+kPFLN2C3tADZqpOHkQ7hIWlACnQGxHKGdo
ziK4+m4x+wnFlE6gGTCy4QBar03ykrMuXOcLggLw9mUcXjEMH4cfAoogYCKzcyUX
Nl5a29301CTBTisUczze4QYyicHbADhGXlM+L58YBqbsGUsNJXBsdqndy+x6XuMw
oFhwm71qnjh7OvykckFXOb0VA3UjH9v1JHXUvfepDt4w4w84sB0+kCBmRuNL/ys0
EGAcVvoqhdmH8DWeeMEIyw/nBp3XPNepm14N/Rkfj5C6w7XZ9S9pjJzWoptCiUyA
fLqE5E4q6gOcm+sn+wpXCI8rDLJVmOHPzyY0slHl/iHCrMvvtr8agxsGx1ngsCrT
cc9EWvFKsSONPwTW91OPSyF2JTS7IrtnBT3uh/c9tTzjHH6RAJZrja1A/aT/cvza
YOElziCnBO8F31tGeaVnFBLMlR8F5Q15Exc6VVDvN9Zp34LXF/qyHqdSc/fMViMM
ir0Dgjru/hi0ZFZRwhdnRup0ZEgisjaJa6G7tXJVLKu+BnChIH//LF9mAdetabiG
VRz+weYga3GygjzEXT1Aw+b+gktZGypUQUgvpx3VgTAgPcfhozBkXHm6MWIA55MS
Daw63GQeWZd5yYMHkcQk8guCvggP9yGJ8E+X0U5vKx9mPGOApapYJSpj1Pd8+uMp
GsnIF+r71OUCwZfGpmxfX+n8Oqp6VIsyBasFvATdbzOTragb5dkNc70b81W+HKNd
+GpzYWkrk5I72pJ25c+U3xrsX60rfkhbxPRrrDq24Nloz5XKwH9YbFH9A7yfEJs2
uOcJvFtaq1JT99IXYt4Rfvv5uxwkDn9/q6pv7auAIJ1ITbvuBm4PK1xgfutInTbv
TNaooT4c+BXy5Ab8f/PZhHGwWKFsjz2AXu/nDSoEugC0hq7Sa2DwslZ2a8C0gmak
OsTbhUyTS6Cw/szePwhlHiI5EEC+KrOSClBbqrcOVL5eAHtVDKZFSNEAFE37Cbe1
L68MZiHSCBbHmeyjuIcHHOSrKx78bzjev6a5upbjp74BAom+SM/D9wS08KX7ezcf
Cu/j7NlYoOHmbD6pyhw3dzbSCawtG7dWaymAKQ91CAfRGhYujpmFA0WkKaAKFvLn
NfFseBYnnLjRzFoRvkZOzqAnY7XuTD01xVP9mXPP24GLQYcerOc28KMEg/6NBqDf
19m6oDtIdpWywxjCfT4s/yaPDUEYV8aDk0mettPyMJ/WkB89ZgC7288jdrgDC9+r
4gO/jr2+Ec25OZ0hLmgQDNhcqU7wnG78LVm2lswRnFVvnaQIuP5bd7mjCKNGk/6l
iuIbNkL3qFWl606fEJtciTOGY3QWp9wlutJWt7c5aN7TR9tSyjg0V844358qD6rc
S7zGbHUcwczjRiB9iRVx2xlMpO8+LpWkX/WNIPULCaUyM91/D/fBxg7GXT2mRir+
XgfyChkwJOpG7U8mR0GWK+CgFRZC/yfJn82+r3K690p5IPUU7EZEqNf+OOH9uiiG
F9xLGGPct+xUpOmf/U2bxROEQ5gI8cFSM+/8xjXdL5mOQAjdQp/Nl/1Tzd5WP6ia
JFHUWglOxVc8yzzsVf7E+7HTiIm2lp7yS+6V8OGyWLnSOMjkvQdqYpbPmQCd+TfV
xD1hjRV9t+C1xim34HIYztahqc9H1cONzo4Iv6zbsB37Q2VPEO52lej6LxfPBtB2
hkDtA99w1/cpurUFNGAcp+UxAWiZL2072kqZl1bl8z+mUCW9fp71tNoL7i2kampW
Sh3t+PB06rkjD/5wlsa5+Ik5mNdTr4OPzND8jXedOgGXiL2kWDV9H/bv2Hgx3YWF
`protect end_protected