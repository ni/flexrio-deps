`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKfyxPA4/qiZ8+Mf4jkKR3IPk1Kf6gD2DwdA2FvEoAnMdZ
qoYD7NN2WOYhgSgg9oe+RskYwqwFl02FGQ9blSBnYq273pOUyR5SMEUKMDRAeI0R
JK/Pj9ZeE1bFAWZxzYALqjvGFti6a+L7SNETSgqUxU1sDhPvG3UpRRDKgzXDNJE6
tg2t4F4fN+sZ/4cHoXrQJ9oI4rZpn2IT5iPQWBOhs0C0ckj20bUiTwGaxslBGSe4
6YctHOIjsE0kBvrL0HjUrup7mpCFj+BfbIBLl7XmO/7O9sUkmE8lWB51dOMCcDlv
jC9A8set1AkovnL8eVBXUtY5jYx1qCe8P/H+OMEgwvfIYNYB3/th9z0C+GEi/Zo5
ffYG0eRtHdzVrj/2/jVOa8GFTtyeSnZCaMIoNYZT71mKRP+fhka+46iRaYWowRq9
GBoxHuST9JkjGfztY7JJ7zJE1MV2QxCPkOHBa31/2EfR+lAKDgKtwfCbIS8R0HEk
m1ri6D/wMX+SLL0SUdq0Aqkm8HxziasrocVqdZuZpwdSSUkP/v2bGyfavEPmpmFE
TkwqKPn2F4qtqEheb0YrsR9+QTshiSZ7yShmGYokKv/fVJfrhoGHrDdLp92PaDya
dipc+ZzakPemonFpgWcIXprAmduW3sWRlFazQUs00m1lgvgsuHlLMg3KF1b27ECa
XdaFvw6akjMSN3T33hhST40/xwhDVTQI307Bawa76uoBHfXW6HNAdY/CbpomIRC5
D2S5vGS/jn56be2b/ZwgxaVTuGWm9F1Ozl9wYHRhpWruhJsmBNVva3ZE6NNcAX1k
OM9KbZbqXGkASgR4Ps+76Mfzs+Qks2DTaG3FfS49CiDxPEdnnfiDoOqwH0xQBTU7
ig47R00RVccjUX+6G9AERnqmDX+BhiY3zGR+2dT2/o4bAMSKV1YLxF0m0y3cHTNZ
I4y8jWBrph7RZjjgZ1c+EwXrgypk9ng9ho0Vw8/EziH3dSvspdTznF5BYkqx9pO7
yt2dTmctWDVM4K7cYX/+2WB73xxOfYvLaPswiwq5yctUaV9rbp+t2M6Lok+Cftzc
WuaZIWOrmKtrDT3Wd8PrMbDuApoBDsHunEI/me59EtM0yPR3USgV8gK70eqW6G7b
6N6YgdsvQX2bAsXzNedTdVfmRbaRGoyao6xU3iudmqcLDEsk5Do5+YZS705B4rCC
aAxl3BQ/c1EKMzcYSWHvXHgZtdCzM4OcMCd8JUxlogsVwCfD+vr45i3Zd2cekKEv
dH4JScOe8nJcWMT/62atP1pzi6v2XFDXml0TzPPXtgx0eV1UQKeuIRiEy9E+BiAz
uZzg3qWkkIKWTgfqcAWzzivs8oSTVyXxbZ3ihJ/C66kmdsRIvRCFcsj13yANF8q9
MQQ7pd/QOgZFb48VAjTK/BTsBbnKlKx30zW+QQGv4DbEudK66d27Pa72lzk84VBg
5dkw+Web447w8oJ/qnfxyVZKyVZWAL+vBxZIH0xX3J8dfJoInNDPnnFUncLjH0Wa
vTjIrfil4WQjGCsrnfWSYbMux0qa+W+dw3h8Idj6APqqw7d6h/cubCymCNdF8SXy
rpfdhUnOVb4I3OWqD2QnATzqoJTJArHgnh1ZKs/C2S401WDE3iZyomfu0xDWUviP
TklTOkUBvkPy9ti/qhb5r2WMPqGFZXZzG6Xpyf+FsyJn0m0YUtOScjmKG784cM7w
jV8Sgz4APckHu1/7ZjPKaQ+rFWKfobrpzOInAfzybE+iZ4Iq3fOyVVLwDRJLVODe
opxFOMe1BD6LUYn0TbDMltMKUaT9A1p5cEai5uNH4RIGQwz6jMXb3ej4pOR1GEc5
PMFGr5Xx5LUc04f7asVgfUOMo24TKWFcVdRnbmdQKz16JlDicHzHL6NSDPhDc7/K
gFoyQW+WnWjy+8/YoT2v/bYONkEh7ja0ql6sg4ucG1ROb9MT+VAlpQCuwIq4ghYW
1wHFsLAeGxjaQq4y+RQI+e8FUD15tguiqeZbozilVzVbB2WxpECW5fArRDxnnU/C
jmWbwACr43owi3oPeNe+9bCWql3zeF/Nzj1vIwvoF+DUQmUAVyLAuhy98LsX3FTi
dPshY9cC87Qiv6YVXT6JIomwwRiqj1BtFZWzJZjoKgr0wpfSwtyaLf6Wt01I81gl
7WIqgQVC7YpPsLapul0X0+ecHq0xnlo7WPzWT9Kzs3/cmMkM6oCauJsDFO6ODIG6
/2r4Xf1+00rMyPrd2X02CEda5wwk8vDyWv1nC3wqGL1iirS3Km3EXQSfHkoLu1te
COy6OAib4tp3jaTZDkAij9qIXEbIxYZ6ZcjeYD4xJNg1mHQXRiU5gZtF2+2nhXgJ
LkWDRasDhWXcFoIUVv18xMGpr/Nf++/tee14INrrBpLZ4S+QEtRJNNUdUG4plrea
HV2wS1bPleL5vg9PX7dMV/j8TKTvz1K8s/C1UNiL94is5g2y58T736uIUlyG+M+V
iIxJgU8//VZE9mCUrkr/pIB2E+1CwIFzdpBswMOibXutB55rFmG3o51R30dl4scm
DqRnJ1FvRkK5X6sqP+Wu9bOXhL9aXseVLuEEGBZENQPsPKne5DPkuTGEOpEf5XyF
gdDM9K+ky2Ypt2/mVi7rBX25JxYSuhhWQ98VlYUocYeoIvP70kD5DgU5fm6pG3yb
5p70tMV/PgoiD+2xNwBeS8uFmOmdRFFRXBVdc9KYfdgV7cE4s9i4W5zSi2uGSj+a
r1NItXnYPxdDldpcY4kifJSKEKN8r8+m0i7iwZZN/t17d1w2/y/vGSdL19tJ0rxV
HbwqCYXS2cR9u8XIXoNuuFrQc8YVSZkHm0SwJj/ZI5vqo4StRygN5H2Ra0hixOej
wkMf3rWqi3A9lQ4ZIz0xWlJ5nN4Roc9U1vEXe67rz1gmKHemZ8I58DW2cSI/u9gn
sdrmAflYJQYFsJhyiHieSPNYtbMuyYffk9yG+HxvbwoWrDL09F19V+PwmgTOZzXl
kC0ceSrC8u4y/T68FGX3USNaD1vbguu1/Nb4dxb6YCJn84fmgtsFuqK9KyGPAAoV
BBKiU7hwnn1K6mi/7FogY+MWtq6bDvSc3VFvBz9/44WSXxjBcx3bYyA/wGjCyPbi
iSwqMFk1TptCI277/CsZMqeZSmHg8pvFHjrQMkMP0cYcsHZLVoFqNtzeV/+FcywQ
T9ANFJ+0xp5P8YQt3CL3N2c5gGn8Qynvdtv3HLCF4TR9xdpMRYWqpcWgHuG648fd
Hxbg0Do4/sy8oZBrDgyozsA1eCt+AhC5RRcGuTJW+uRumAZAndXT9uV7bwLXCKbZ
BbT0Q8ckqGBKgMtENQswXFJ08xgOqOFXcK25XGq0zEgwKEM6MraaK30xYhKzAxSp
a4eAbzlKrribFjbxX2hUdo/ed8cAFVhjZWLdBPESwea3YftEV9ylcujP9C9IMZDL
hcO6PP07JAWP764+8wYvhebUS+xvMiDg4yy2YZsv9rv1fyLwkELAUz+B4S0/35Ir
qPPhgrgq8hxnjIAayxR1VeS7zHl0dU3kUKwpZbtxBsbzS6Z/r1S5zpWlqniUH7BK
jAA9zqztZeGeeCEYc9Al7ToraN7rV8UZtMmAjls3JC5FPwkC1EMNWAHNE1BQU5vr
m+/6S+sIBqJRg9QJxgNk+bSdU4V/mdBn8mtANoj/B2a5nA+HK6L8d/eoAhGdDMTB
z13jPNmIcBTOxjWUQWP84bEEL32xZ7rZsAps6ijW3OZYjYkQYvOFwtSiOIA7wiYy
2PkOtIhHb8gg9I38m37VliChyQUrRDjZ+ozIswJIezFLOwrSeID78s3Dd2D7iMev
pStDZYy60nJ2praIr12Uu/qBw95pRYkKaLROIuA8mryy3ZfRpthAY9c1iuYG3dIv
uSgtm+uMOrZY2GaOXOZDZOsYPhtluTF7jiu7L1yqkWJ668n9lbHiW8fEV24JBtT+
UZR+Uqacq6Jj3mi2xiFUA6qtur9ZnJmDf1iF3nJzES+TZ8INtk6ChInQQcxOJxAf
wlrt/U+zMXS0DHqEng4bU8C5jVNYvpuKA0SCgEMEBxdSm3HjC3RhCiHgbsncHcRu
UWtpgu/9t2nRCKNeNVjo3DiGHYnevGf4anbp7r6aDn3YL2bFPRlz0U3RIcifJ1mq
0K+zPsSyGHcy7ZfP9741L8M734a/ueH2Y8e/RRVazJGN8Kxk35Zlc2cxPblIodrv
MLvkD8mh4CF+RAtr9IqhAd/LUNqgI7hZzO8udc5+Y6zO3u6u7ymoPFwHnCN6wiyR
2Y+ymNWOqwtMZ8Hsyp8bKocfn638Ml/CtcT4hc4fEdw1s9Ln37OnckDEZ9xpVmAS
cqWwGoNndUU+Y+FJiHOq9fOiBWUL6u4O4EeeqWAQMHukkJlpP+LuDaDPto5DbXyR
66/cnNPP5QHKkrlj7vvOHsabwVL4f4Q89Eo0tysE4i9MC+zZWPRB/gMbjIAUpcPC
sa6ohr2x/Begtq5trpNqYjzZr5UyIrg4lk7geLkae0DMIQ0pJAgM8e5tKzoTXV03
HQahHPd5iDqO0f6HdmK1dTc9kMovpEou5GaM7+eQbDtd0m/dV7rcc8D0aJ6l2qhQ
kRQvDRPUgMmQo+JykkJikptj1HysDbyw4K2YU6+pttD5jJQUpO+QnqgNS9SHNE2H
BPB+lQRWfsmHIa/sD1ediplrDr6CgqVrsoqWS0mphjXhCftmmoehmZ8W8KqMOBID
qujpibYsRYp69eoIYBcorTGH3FNR/u4C0uz7ukN1bKbap0ykz3uLTHDJBZk/wpfy
Cjjx6ncLjvQYcVTBTz1QOs0TUBBkgRXYp9biPV8esVnH6XR03sN6key9WyT8xRRL
aTgNJHHmz3BOuu9TZuekV7nJWhg+1pRzn4lkmofjGVyiqa5p1ecLJGaQIRgUjxDO
sx+IGLkd+cONlrBnDU9C3fc4Jsm5OaZxsTDS+CbyP0ixsEd8j33uSIr7D4B6WZsh
15GFXOv34u2z7CRvqvS0XHjXE78T7XYebtqELRwl14qDx4f+M6mvBxKPT9c/vmSK
a13YdCKF8V0tmEXEEWK3bH/pGgQ3wu0/TCNf0rz2Ms+eGGAoRRf4Xbg1JwYCSDSu
JlPaEYTrouMUcdlGO50eQjMuYNGlHjCTmXaNmrOXaPU5t4P0bQ4GBXO0s9LMXcXA
beTM4NiD9vIJIGQu5NKBqAvV6vMBMKVvj9TFHWEiurOQBAWLV7hzgIWzUS4mOimW
IFKB4sWGJ4amnnttW65tFrNRHWMMX7eCZcVAQYdtzeq1XkONESA+spTApjwznsdJ
/8KkQVR8Fts5BB8HwnPnzxAi9LNP5TVCZAHgz3EITOWVHJ54QmMYrlFDJpw+5lnr
KU18j013xYQkrF5+P/mnCmR4TDTb6Jo1gSoYTtzqi9YA6ILizbvCy0Po5wkn0D3Y
r9uSowHVTkCjiBIcGM2hh7oeLh73ZahxXhS+WOg1KbPxOKBR9FebVUA2yXJq3KDV
imDzEGR+o7NgqIzOLlgstQ13f7ivD4XjbIrm9UxiQdyFiRo92+4elo3yyqhBqCMn
UxAaWPksveEtiOWW0CUXsTxNi/9blwTyvQYoLeJW+po1zGmnU0W4YPpTUr0Batgo
IpOGFqHEe1RQuNLT1psAl/04z744WtzGhjHBqj4XN55158DDLO+rP621eoI3fsqH
FlLx4dQZ+D54fwO1Es+Ff7zj6/HazQCsQibOFwuIwpPsYRjKZTE9xv5ENDlaFffA
k6jJsWTbOahsJfpQqZDS28WFg3HdJM8itSh+QIbRg3o/cXNnjbyUjGJdygEH8UtN
QOBQj/s7TsiApyanC8tqQJApKdSVShElCS2agXvRvKvETyyUdwG1iSxOyp7Jdvmw
e38dXoBGLsActi4Jn5OLrveIa8mV+EG2N2OqDfl34HR8LTGzHxQc6vALEnjIRSBE
GLt6b6/20cLCyy9GNYrKT0EZA6DOHGDuK89GVuH7AhPWkXn4+z7tuCeiJjMs54KW
x/M1QR8iTmPpK5YVktRoNH1TOpRguiH5zqcUx+AZvl2sIf/HfNJNJF9Yf52vj1wS
vG/vRcnK5SAy45XVTA8BSK1FErgFMOYIefQN2Atp9CInXPa78Co45WSBc+pX1YaV
5in6EiyVVauYcksFm8A4t1XZBVf6VC7QBfRtwqs2644VlRbaH88KbRtYq06r4K6q
B6Smho2AT7mYA4bS+6nxZWgoq2n5CH/74GqeMQZzjiHPeEOPzrw/ItlGQ9eMPkVi
IzgunjmFPHs1zYK82mHFogHEqCY3zQ3WekLqCjnLXjKIvKT/ehSqxLUkdGIR7aal
RG+R8iIWMRQjoV7cPkhHABUIRhHopUWsxTVj2C6u67k17uAPaj96joUaOYxNeFDe
5aXIttVtvkjKYYrDOw5cqSkPQSpJWyKFoPccX7ECBdqodQFTL/UiZ0kgxsxxSEzq
o7x7pHGN8RKvPJeE3lDWyrJwgop/vn2vlHETlXEiIwBMUD158spwUtsA/EBFZFwC
Z6XnpO88hkklFhZPWEKsBfMFDfKbbEFEPZZkXOg/QTo1MDuB4Jf4D2+KCk8XGuvB
a0cmK4N2TgBpxQ5EYwxd7alIB8/SLlckbP56l8smP4yQB6jcHQiS/gcxjBPhsiB2
cFaJojInif69hBmlB6fViziRuS10/CfrCDzYK3QMdzPasIzAJmBee0y5BGRjG7SD
5Iq48MGY+XKEn50iCeL9t5SKbyzedtAOk7mw/oYp80BtAvM4ruQhph1H+WNipaF6
MAPvp+oVRxJ3wgb532mUSJYDx1aJ+hYNw/NuUCf+LjqZ4NNfG2DNtolp1Syz6pOr
hAJwCD/YGw/SjDZtZj1v7h20CH5iKLz+MX1n8tm75bmM7PkQ7ktQgMrownRb0O6s
H94+PcVrFZ98IP5CsSvojC0E7BJzepcrtyEv+yfrCGpJeykior0i4xY7WtoLqsjv
UZyfRbO2EMNADc1DSmhnNVh4yr4mvgByZyXo2BC1hjWfAwDXSBo8J6tRGWSFeoxN
5pS3t2tjOK3IzwJd+LdkZr8d0UYZF5UbTqyLhFDoIFbmtIcwdnK3rwm1y/2gbYk+
c1y/MEEcKXJgp8gExMvYBLjvNJ+rmd6wL/AYhC1E11mxqMB2EKdl2b6UrwKbphcB
2Pq+g21BkVUc2ad8eiO8lEyilq0wRlyZ7eXIvO1h+y3CA6rngdbXTapTF3XavWNb
aoEX002+IzFOmHWkRFbbjvbVigd6vqF52W63LuBZyaCEbPEJe86nXzt9MlpAaSS1
nxx2RdezHKe8OXuqVSEGtHprOC+FydpuVC7AfZ58igTa8bmEA8F8eaNrcstFPEk7
DxzDJSbvhi2cndM7xwrSX8JlmylNXl/iEAJD2gMB+zivj5y1ENDcL6juseQ1N2rO
ofXJ6i+bSvYsdKXOWsEUD2+1RsgdWAtcbwbEPHMI3qofU6HYFThUgQvdlnuSv1xO
W/tFEg7VcxJDiartmyX9GnYOD5jof652SRinDG/K6XCW+p8dHSd1H/WhX5kS7HKQ
Kj8MVhjkC9qw6Ged9x4zjkcbqQ5+u5g723x9GVBnXTNSRSObBKnQYbOQAyejSRHA
Az7Q/qA2RgEt7215qSJ2Upvigpgm5gHW5QviKDEvozWTNis4bTFGaQUehChA4IM1
2KuHkRwXx1C31/qsOUpdvEO0+xIklB0fwK01fn1g7nWsu8VbihcYDRbzP93bkwqP
mdMsMv45Z5XUFp8cV9zjO2n6e2e+klkvz3MYnwk90TQqLy1tGRbivNBSFVFn7xzY
D7LLOAYTjc44KeH/Zr5KyOEgAL2TtNgpEMI8eLEulC7T7BeGOH9QneUeG+lgp2NM
9YLNIr5WyNjyZvHWWhqyLPAHc9TuifxZbeabvXBf+yeArjxod7YxgK1upSTuXaff
xY6g4MwxlKomH2y3OlHubB0vqJudGdgiYGHYKZC2WffIwV0XVjvCRuxF7uFpJxI0
gxUbQD6oTHlHgpmzoY/UyI4sqrchQ8mjjWeCwA2bDRzIK01X6gO0A0Dn8wAAw/fQ
Xz9imXa64pAXm46C6Xge2n3fSxuSVfnTJrtaKSzfwBWvg8k8PKHchnhAoNaeFPWQ
+cTB5HnWRRzMPo4aG1dJOK67NsjG0KWX3d8dA5n0ZX5xxrO95T/zn87IStPHfg4I
Wly+8WZBNGKkMG+4CpGQehbUQ1XXJEw9onBcz6n18P/CZvw6zFiyAl2d5xCgZqd8
QITP2OnKIlqDeMR4T9IqSrsBZCCzlYgiDGuBMyxQhsP+vafDaiGOJnlAISWjBAN2
QCwtf5HHyI3dZ7WMs9Lx/Eg7iQnrgsQy8WNqBhIrVafHqVuaWgGc1cCsdTYkHZW/
+rvicxdP2sA+ZbYXVh5RlMZd9n6y/2XIPoprwtuc1+2ALjZF9zvB3oEjvAmk0DBu
s/PRES5kXp6u+MdMsvU/QalNYKK62PXJ9ENssOosjrdbuhIVfZmOKm5yY7yBdCzB
mZCEzaxKKX7WN8w9vFkl3QxPAyusxpYBQ3RKBRjHuaFofCZB15FuryMI69USx8ws
0gHDC15uEu+eVm1W4eN4wOV6LRSL0DxSe0vVFYHg8VjWS1CkWk9rpfHk7PqqTKky
tDJwwN73qtS2HlqS/JDHa8tEyDPYuO3xWKx0lExjZTrNYpE783wQ6RRUAVBVArSN
oUhWiuOI+MV/Mj+hqwy0cu97b5oqowXL5tzPc4sSAEwxRjS6vrZGA8iC2fScF+C0
PKK+xBoHoUr/lxDbve/oiJUek//vPAxOcOgZpcSu0Y66AL3R1NOzqU3WiGvhBYIB
PLukGKGrxOu34lGzcpm2EHhJyeBCei2WlOnsEui0lOFbezo8QRSl6yMsM7JXlEfd
YSRcdyhRlv9pYGy+uu/Yj7H9H3/AM9KPlbv5//mI8mqxrgq8o/QnIM04cxHQWgrR
H94fRRi1ccPXvXdtOyB52Cb1Cn2whhg9bDu004GsH/drkeZAyC/eYCA0AJFT6e+q
/WBy47CfYjodx1n6+prKIf8aXyrUkw/ANPYovU5p2q4+ya6Fy3iaf+PiLH25DPHw
HC2r64GUVUmc4zf2XkFw5xksl1JKKog4ph5fUfDE8hackpeuWQeZyMxh6jqfYed+
+YIjKTRBAnAKaxTC9+IDS+oOfs93glOuiJx4/hmQG//CSkZlPeFAZrwl+zR5fEWI
JeusFjNc51cjRH9pcSNQU+1Voa/TPrpzqRAQROHORslFYGHarjJ9PX5myhcLjXll
h/fJmTnWVHN+j3xJraQjH0vjwIffxwz8E46k5K0SxMxeXq4uJcgYhWbwuIIgmNUr
c0XUPKvCeQH8oj589r9LXKBXarasrf87+mLja7jOF2D8RaMjWPOIKzSOp3Rgixf5
4yeu4cEHr3/5Ag9qOghIzbwN5FKkQyakLAkCpiU4vPzziCwXsIH4Cmm+PjShW1Zh
qYRSFhQCwd0T6HjiyOILceqV5Q5lyDFjo2Iny7E5hk+/btwLOq/V/uNlt3fWok3A
mWhe0+AgX5tDtbEmc81JCga5VcpRWdVVr49VWdsb8BAexdTMCp9C7TRo8k+4zkJO
Y83BlsOqd5Fga5I2HoMaWHn0EQGWSmTwEsyXDPw6JFrbuKn90ry2hmEtgQF76HIF
PamayYGiz/uJt8ezmY8L28mtZRmNc8j3IChlJaHjHpsSEvCMbPjTTHibYOOwrE4Q
UKFeXtEUKaOqdAUjCOUyeg5m2LyvX2bmnxDPlICc1QlgwvibBb2yae7TVoc4sL4s
Im9l5SycAAXQesoNWC7mjxwSmpOvriZ9t5Ye+MVHKsxzbT27IIxzp1V9mBuJ1XVO
amVugGBDn0Gn6MqblCctN4/uqGB4Z+5OTC5h7Q87c8sbSGnXt5PlNtwhtBQYhFOl
JGb55rfd3l82dRaTULK5EfJOpRNfU/7M2jJRnt5loblh53nCGKl6WVgaJZ9q6Ofp
Iyjsmfd1HplMZeAG8bDFWbKWMof4dL/svmrWfQiS+W6UE1q5Wy+/tfpr2Hrm/3GW
kzwgADjMcZOXky3KnPQOrhuPMqQ13TMVMiYRr/tDNKcmQidzTxQ8Icfc4ZrnrK3K
xXNKo0MyDRe3ZDunadGdmwbEVJNfS4DW6Va9AYvQm3qWajrzWL8BmU5NxrkCELZT
Un5BNgPRwkr6mxVxhhXT2OXb48mtDHG5r4i26ktpvSF4VJdGxBlKKpU4alYid78P
hMpd1dBKK/5mjlTEuSg6wZSBeTQz+75YGc5LUeuSqoTrqcSb0RM2RkCTO9MspQwt
injeYvyUEKxEEk46SJHJyePy7ps2dRuVIzP74Po7Hg7vXcxCbE6Zhje0i64JSBP0
0NzR1wn7/hjeJsAi3Pn+O+qhHiZdAvb8dHSEM8tJj7NAC3rjoEXpannwvEEGqTEA
C3djtRnuNHjy5ODFOZ7hqSQJ/hLDS+pivPupjntWS4LiCuIeEW9X0NkrG0+5Razj
j05UMiIeOwa5aKZgrQsbk+BSzKzUT3b2qXrT4SOJfJae3huB/uslUw5SQgO5jO7g
HCi8pPRBiXF0MmIiOUDznP22ey+qFpsklrLOOqkmb7BBjDsgqwe+o3bIwTDdvf64
yf246T43QX/rt1OPc53v2uqaqyl1bpZLr/WFbVa3WW/I9xxVrwmDT6WlInhE4ZNr
dkzEZ68sy4NRs5V5kHnWQX8Sx+XeFQItCy4tpc1thkXnMImidfmKHtkvtl2wWqU+
wszQ4Oah7ONmuhy1c0f2Y43MVzUMpKB3qMv7akPSWrl4bp9ae3fcSWQUsOVW++lN
7jA/1EqtvKhd6PQg+jmlkLt6DbuqNlHP3q5oGHNzXOjPBJ5WdAAK5HEwZInvfsw7
NieYC5aRmwsgAB99tnJtfLROVNi6RbCtwDZl0/EyYwIqVIcFqYVzS1qcdhgSr1o5
byxDcKycx88Lzqyhs5o4WPR9qp5yvShsi+irfihB1UqxbpDTTlLPHOiDfSqj2JNh
vRtiKVYDB227SmPbtVH6hB4akFEQUKJuHwhPNQoLadPxVCMe4w0j50JzNQec0Ekd
4wlMsZOCXG94VUg9VmZzS2ZHCSvdNttg/FxKCd5dMD67nJHuChEBsSq2taXu2aM0
M7Mx68xVKgNdI6r5WIyJuKo02VJncBRz+tH4XnrGAAjUqAcUspsygOLyGARKkF5j
DNVuTtIDY1O5gTu+DhOhD2aiYWIYKMZ+wctf/8C8Vw8xBOOYG6YdqqhH8vwKBu45
EjUuy7oN+R7125gKkwwZ8rcT5JI7AT48aOCpq6n0PcIaPqbvMqrsEvis89T+1LbO
fkHOD8Oixi+LXSMIbM2ForPzQUZiIb8TPeRdsKjRRfyPr4wNUe3DbOCjeJVkaRPm
oreD2PhF0EXZHsTyHY1UVch9dtObASRFBwB0q5/L7q/6FUoORPUpKpYAOnOKgVkb
JvXdiAOelaUku4P3MDQi8eqlh1UZp7RDY/Gvw01CmrrG6FLfaxUKGpOjDaCpQB4P
Qc/WZoNI/kw1EZwZIl3JCNvRbrrY3fwKh8lHoR5PYnqedhgYrrvOjUx8jN0jehJm
YcBKv2zyXVsi0nbDZPkBdKFPKsQ9vW04xFJwC85jlmG3JyWpk8ZkmDrJYntn57nU
t41ZqsdxC8XtNX30UzxRCIczIIUWWddzVOeU7Yj0IZK86SOiCbdlGPMluoF3xGaJ
owRydm3Fg2NB3j//rlKphubUmV85R9NMq1RDoQbqU05lTWitMfKM0H/ox/t5Mvq6
ywTLmgnIh1OsBgh3W6DsSIt+Tvhv21Hfd8qy1kGGkBrzgoCWx4d8ESGLAHm5Ul5N
71v49KQf8+ck8rGnHLQ3RjkI6ld+CuevuUqC1+8uOHFmHF4O/o60yA4eno5BNnOA
iRlk2FeurwF/kESaePD+2tOkvjXvt2W4GtTkimh6Y9rMqud18o2OavTSNRSgmZSq
CYncAvvoj7vhTno+TY7LV0qRlf6grvqQ/2cX5Ce/OuTKEgp9IOmZEwZx4TwSUwoi
Zp00f5LtJkiBLRVKdiRPmpOYgOATCsDmyq9THKrXYfh+rDsj+ej1H5OHR8M6jWxJ
0orNF+u6z+BmiP28ZySqkLs8I0HxGhUitZoSyuu6pDkJxB8tPiRW/jDjlU9qNASm
+hR0R5vo5bHtfNC9rwEZMcXXrZJjtXD1yz7YNE+nUHzXlc0VBIem+sZxaYWFP7j/
cS+5PhrINkGPa61CUO9xmwfI+q/xSovg9d5f+l1JD5nwDsKoKQBUQI3IYJ+WiZpu
ynLpQZAJpd13mKet1yGl8nMjS5YoHd8EBMYNRjlvEKZwQneVYIYmyAqYerbizVK2
rtLAr7Q1uDecvVA6MQa/vEp+YM/wgOQiT0UdGXt/0X9f0Y/bt1DuC7NIzraqHI0a
9BN0hMIgZJtJID2DiwyZptzVwfh6mROyjT8QNBTaC7j9WWNSMcDBW//GrDIesRhN
mzNpkV3G8+W3BUTdLUw0EoXV13k/gEka0fRhPm+XyQZea752A6Cvj+JRVo6cB5pW
iNnAEXgSpqL+5D0U5PnGiEOLcNjrgljE/3U+KC1iUXYToYnFGgGAU5yA/1heoTxz
9rFQTrp/5GGntD80Wnv3KW6fEbqpLYzCDA1exYe2jWlU2YrWuvEvwnxHd63Pl0FT
jCM+yq1/eAfaIeq9qwEziPFswkbs0u0ZtGB6GbxcA8CUGu1v/UJH5v8FFI1BSL30
ZmzXYPp/POPQ/uu0Bzd3AyaU91v79Uf0q9XSLL3cpzN7VrKEblXVNmYBkymmeFQJ
GOu/QKn8ReIQzQky3XSHmfw1dRwEZ3IzYDVEpqYu9niZYYwyVGKBD1Fx3QhDncFw
o909086THyKvXYMHo/aMQK6SmpYguT7q8VPimXhRY3o=
`protect end_protected