`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNY4c38GZNaBuQ/jrKCSYG/snsd13MsO7sz9uFEwXdfr4
g4thsDg18rHlq9MyRgRyP4UCt1zsIgTYS2F5xeGWsvDJQdweEorwMc22HiDz86G3
fnQj+hhwaSQ7z/CyUIp8AVPywPlYQPjA2GjjU8e1S828qWRelJF9fCKHaQyfkFHd
ytaXcazcEVbrjR/DO1vAn4p6+kiutCwMtui6iH5liuP/wlm7XSlBLrKxgfTWmUEU
0IzV3P56oHPu8CzhDL0JW2yoYCPVN6n9lACngY0ewhAoo1EwABgT76vCeO7XbtIr
bx5MAe8FKaHlF5Gxv7z2NrWHy1gOaZ+hXtFX+C/UR89W7ha4ivdfzt50lBoqMXvm
G1hH8RIE7SUYPB59XIVh4O9ZdjJczH5nNqE+PrfdQOwK7zhv3nsWIYSNkzKobMi7
QoFYydtefCXesOUhoyv/PaHH0IstVKchr/aQxV9bybHc5F4CCUX0RVIWUMJCEITO
1tAKcC1ALsc9K10lDzBXOMtIVpl4RIZeR/LGAO8TECN0QOE2rZFFOFHDZ+UhE/m8
cqpsE8aBsN4aTnmr6Pu5Sy/uSqUdkhCL1KQ0OWaE/NEAHQbax5v9ZZTd/8baRqsT
y61S/hAwwrfr39B4Nnzfk7NVOzD5H4JIr/Ig6RenNvDmZccecI5Gc7LpqnUQkSvN
YGSq1IgvAlp1AhYcNqosScelNr1wVHSubrixUxr4pWvb6eWCZnNuOZCi+0rRWUyx
tBuN63dtvKM+Ath+ux3i2hU+qx3ZVTiXroRYHB3wyPPyKG4PopNde2NBKlXlUJYr
MYyh5vlCZhR5O4MMX9JEUaRMs7YOJCz9XrocJ5KeLZfc1jkQZySSAWtZr4BYNiOv
OTeEmcUa6apVWxOHk+esMl4NI4Mgc1T0AwHO6izTecyymCs6QaCTyXFBmXjEifX0
EYXvOkwDj99+rcR53a1U+akf6O1MCYIlG5kWqRZVmwhxlr0X1AHk6nrx973N+QAY
V5JRAnDopMB7AlIdsR9QGqSasl/U8aNIiiARb22GQaWfWvACCaEz0ibyvqsEzKWn
Rutw/B2wuhCsaeWb+Mvfbf0LTELwS+4L+3ioB/sktq+6d093dSnu1Ir11sLuLvKX
2VWHY6XOzPQS8i1mLla5fEdmH+Dc2Xn5+CEPwDN+Ibt7vn5teK8kzzPt7tOG5tbg
m3M4fMEAUSCX/hm0gomtJDWyWBm3LxMB8mQecdGiJAlkZB7jhqiKtkxf5yeZFAcB
VqRf2osh6CkgtCGKTPBPdG/aE0yDKVn4ky63N6K1TvlepYH930zTB1LSZXSnmAQW
jK8c+b6fIIw/cioZ1/Gqd3vxHFrXJ1AIkm/bKrHo6lV6SiUiw4LcfsymD2oNuKhr
EGUKjE1TYuILNvHXFbIUwnpNHBuquIpwra+DDaZlfM8Rnc9VaTxZegUmjBgP5So0
UPdDvhqYuBtSaEU2xULbLCIcLaRB3jZ9i/XJC1ODug9EeZ0Oe0j8Is9vIrg/02Ye
eGlQEYhu/jtpBT3N7zmIbFJgCnWVqFF7DTKYKVfwPpUPLQBzin9HRWE0POB3OgFh
qsgS9TXSn1X+7t1NWncVLEkwppwo119K7vbETw6QsCT9qRtR2S3CUgwJYZTQydEn
6PfBJrISVoMwdZ6lW/hShreH9TJ7DXDy1Cou6Rtgj0Q3tdmJbbEX6IA/Xl2t/3tP
XQKRaFak2VtUOBPwNXXxtAZrTtb+pgkhzmYsH3d2BTdM1Uz7tDFUpcQ5AdEU6Ckb
ES9pAFc0oaR8FTPelLTiUkgm5rXZZBmCTNcActoZEx8y1aK0XzuselaHBHLIkVdg
6BVM+wuBV1VD4VWVH0W2AUIbrfQGWFl6Mlc47VnpfnK/3vmM6VTC2CVlfiaZesbt
Chvy/524yaRxJ3jM0v4LeaDZpfChZSAzXJS/n+l2g3NAJ7AhXaong0v6i3E04+Jv
YlaWvM0y8ez7BSlLVDtoq99/Qq/bVfDnO74zQU3+pTlr0tHUEw4bOjQ0YvA56lLW
a0LhdnWUunpnTFuKnuqIgJOsktwqVkfgyN6SewS5I5x7M1wsNHLy1B7ildes5E3t
7T8sX75hIjI4C/hKh/Lu9AGPFgRAYef3KOoPWn60JLD+NViA1lvCAI0G8X8K5tj6
wjpjPxdF3aNZMi0+I4Uoy+eNvuW97yWV6LfLXOjYKUS9HLsU07Yw1k8Hbs1JoayE
u6dOkUHyIJ+Rk7ywphbiKJMS/1RPrfn0bCUr9z4zi2dNnfap6Bn/0vQQrM6BvG5x
wWqnE1fRXcTDUFJ9AqvAXL3ted3lS5CdmsZAdr3vP0EamXX/qzPbY1/l1o/+cvZ9
4PL5porU6AcnIE1TLa9bzkWh+JwEsY2H2PrU4Eb7HnMbXohf3jyxD9BiV3YUvzBZ
v1EOa1IIyvwvcXCw0KcvNfwALTdYAUdOr7Kbff1+VbBMb/izIBtkDjthYc+9aLUq
/i0dBneW2PTDnjviMSLaHZ+ffXzjACD29c+AQyOgtJm4m5MPSSgWF2QmDNnmwd3/
Vk4OTqyrxDka0UkNcJbK9+3WN1xPx7os9bFknAi83aq4JEKoMlt3Ayk67AlOLX7K
V+Me6ElSu/gFwtypsC/zGF6wVceLTV6sqp67CI1t2xNr+4VNu5cEQNS9iR6PD6y4
29KVMkAkncs5Z2IMBCFgrAqWJAhQIewFChtwbdTaTyo+rt2oqpiqUTJcXtisQ/qY
zpP4cDEAo5tLGWETYRyMLvIH6tZjrv0P8wL7fVGDJm6iM/oubu1MjnpyN9h4iYKJ
CAUPRopdfmxVH9sUeX/IHnHh+1KRH3Mnyr3NhHV6d9uACKfeH9IXV+Sc6mu+wVYE
knyjid0qy2ciS0b9DYLZY7p15P7OtWroKG6tHY9vzhBFk669h7fdLl1n3utt6rWk
/XzUrcSbpk+5ciBw8eecNIOm4uk3ccqbiC/xuiUFx0zVL/cROIN2Eqefi3izRi5P
AuSvTESqkkpxoBcCuP0TGjxd0nZ0cY/C5DDsoX44Db5UuyaB1CKmQ5AOeZSW2FuP
G00MnkniE4QrN/TqWRLlWiuCEtyNcv7emr9egGpZYe4OVAdkfx1jFLyv59VujoXL
/o2BHhbT1gUcDJF9vyqgt15bO+bjxbWVpGs/M+9dQ22JsV06RoeAaRQu/+7MFlMG
hOowPjAyfbqW9KviSkBxOF1uIBsyuK0RtXSejdlEBna+6FdRm4Appiryzapl8+RG
WRwmHeklGxS8GeyEnU06rLC5177a0EN+z0KWop9/xDtBY25AWUifl5x8PbeFB3I3
YGjr3vy2OUbUxe27Qvue/2aaukD/qe3bf5WwMSepnKUPlh5Dy6af91lxJ1Po5mJC
Vjo4ixyuDA63g7q9bf7/cx3XYeyrpWLaH3GWjhJbTWwEdj2gWdL/ISiOwkWiVtgH
mgApbTYFECukVw2gASuMMJ3/ND6r/FoyOkBue9Wcy7pRp6cbba4eT/fzLcaBoYIt
OvB7RnlJR/KtM59xTk9CbWUZ0ce8GwjhWsQ/dqeEoxuA17srVb41J18R+XFVyztJ
XvcuL+UtqsKSUjashSyOoDxEc08ZV57uKGKTntvMGgkN4g+D5KqhkyEbh9SESVzA
8LBZHIybLkb3XUZXmuRlcL729XAfFZ7WvfPwwlb7gjqdLUnPPxbDV+9ppW3LGhQ5
0Jd2gDydd1163AjJDKahp6wYDT9q6bX4nYo9zDkq7not8kC7Qx1FSa0hlOklyRph
kTF/qSbp7UbhXZEPcX5bmrEn+UVIRcFZGIWJ5r1oABr9Vo3ibUMs7WNQlAvABNFq
t4pDXwTyGmWjFtpdNX0uDFJGvFWe5r3TsQbKfLNUEYUr97qmoCrcSmPbKkj2V3pN
+AZPjkDeJwPgZgHtEtf6lqGG0f1Eg4PZerE/HmHBJ/sEKE1RF8kXZuz3mD2KDcfg
Q//Eg7PdvkTIMCKl3xjZT8M7+NyyKscHYpIvdwu6/dbekxTzf0Dv3aN5v6BIUdsR
hBL/8YHzA/X4Zb7SbqELrNfMjDbUdAMSNsS6TpJbNrXdFQESGhAs49Mw+NnXUNVm
tU/L2KKvo1Mj7THZAtDRrVvDPEOgDX+/5im0qr3KDhZOPQOlnM3NpDIvuPgRlulq
4UcK/95HCOc32pU3K8trqGdd/yw7qwPtwhHe2/GW7yjvAnJIoSI+9sENX2oGVUVV
BCFDbHuEzhB7zANuArfVf6SToerr896sVACLHtgEbagPjbhrDaVWfifop1rYMnJ6
J2fpbnvUkP3iC2oPJt/5n3jYp32AsdN2yj3/mUfUnN4DwfJynu84ljo6nf/8Pgd5
XDFZf3pmFQNOju+dEoMrMenKyG8jsigCCCt5+SU2Ywf3mDDgBK3ZZyOZECQizpOZ
c8gXn/8lrF30TB7bv5MVerWN3c4Ac/OLsbcBVhnKPnxKbv+vcEGmYFcRiC00Vn75
5z9jE/dKX8D7Do1vqH6KEeviY1sCkhOS9V1YSKfiReFpVnMzdhxdkA1RJDJk+5Jn
rIwX8kCItim776hclonhqOoTc15HXNIuATHXQ8o0Kv02CR9AArEDV+rAsgODXOzP
aNfjv8c4a2YPPThwvOs/RFIT1VFdYuGx57XG2u7utOYWLmR1rDqVDQyY8L113Bm3
5nvmSOfX//1iZl/t65jNSR5azZEAjMPIo31imLjydlwCQ+wVk2358s/wb3vf0IDg
UZQK9PUICHbzEtXUOY2Dy5sErDUxidVUNV5KLlpPtCEiXp3WF2vAAe36y5Z/Spw2
xRyN8Lgy8XCUgytBeRixwdIsI499nW0GyvKjYNbCWlvga2JBiF0g7DqVVFD1Eq3z
Ev/hq86Z5t+GvuS2ptZYrS1c+1Ca7Trv8lQBU58iljXstMLrVSnjdSGAkaZJBJXY
frwKbyP1vTV6JwFT+PWUbyb9sfVlqWYC1LRZATeWeDvDmMOf6UHmXDSpEmub0AL7
/A3n5N/LQQTBLrik4xWQ8Msv/luhP9POhmn5Cx65EcZNxbmpc3c+UD3pwzTGYhzE
kCC2Bj6c5NSNeHUV7AJOeE8u9VTgvqE8D9KRO0kYu+OgHsSiy4+uOqU5kHhXmCCr
GN20zYZHS9a9JPlrxo/nQRF1VmzhE+yadrg3VcbGYZGq/9VapDj5UQkGF09aI9Ji
IsVOJaPbs7vAdEI5Hjli55riiyozPaumoshdHVrwGp4VnOns4xYad7WCrR2JSKYz
1eKCckuPT53i69ZKgOib7lNxApryPKEDmiO5228zsJFJLCE7in++MtNGKXqlJiDf
wUJAENi4O123KXU2iPxCNyYxppxeXOj9NyEuZcpUnvnASoH9j3K4SeayV9enIFIF
iz8/NYdAFvpAMbcCUHn9OPfA0J0IJGlQwp9hSwVD2hIDcy1lbxQyEzTCQmWEg9Ro
LQTPYtMpRByimaMcbBGZXM/hRbZX78+1Cb7BKiY4vdPAIovewFdEzEjgpxxDmfoJ
OqseDbLWoL56T4lLgq/7grruqDQxs2qavPZmP5UCv8WKBnc7j+blBtMAK0P7jsCB
WMD0p4N58IpMkiQ6mnj9Y3SbmgP6fM3JDSsqynnVzfPKrEN1EvVz0c4k+gjVNe+5
AqR9gLQkynf3N/oZEyga52JH9SmUK9Kt0Jm632X3xmta4hKonh58Vs1ufGH4dG00
KReyEi+OZ1rUFdbHtwX6gB3FiPDeFy9mDmw0UsswtFReTXw+aZfTvkxKHQ94Bfxe
yM5fHjFBn2Vy2LlKzM9zFnyVFlizgBG4exyjYe2kUrEHm8limZ8hu1K0plnMYH4G
hd/j152bjsGJaylu08kNEgzKF3DyIdnxZycqHVUWmYxw0ffTflAemvm32bKG2FPv
ksSRA3NxfIuGkq3Ze/76EmzU1ctT5sFvTE0oAAeuZbDBbCrnkuUda520dM7WaIw1
rdZ4Rs1AVmQJYYsxIYPmV3JJj6JB7NX3CCqKFKFVKEL3JUc4tAKINaG+EvhopjL6
tA1+kISaC/8nzNKf2X1QfrgLyIPCLT2gMjbhnE/m/cXPnHB8Mgxa/QaDR9g50yQh
6WptbBktpt60QbOXBWO0/brrTd2cdj60GDwpUBVjFqMfrtp/VjDHzkKefOxK0Gti
ka1E+2CK4MtKcLmRHsBjH6csigP4HhTBHHBfZ1XggQ6i4cc0Wwdf60WslKuu+Nhk
sPxFFP1zINXR0LDChNLFIccvXTtEvGBlmg3dYximeSXURO0lUXO9FEaf9RHx8BaM
9wQ8U5+x0hHFztjijCBFJx7/r5+L2evhIEBkkiUKfcshjsZWPhrtwS6hWOvlvr+R
+h1Aj2+Yi9Sr/Fg3z00Rjwb1SwFYssG8EGpbTjNE4SW4UtjEpw8cwiltox9+zItl
M/isX0sRlszweg3Ei8/sI+VNYbA0pnzbPp9b54yKyXFIjufZ0+PIAJS4lMepkcfY
PjVIKy3UP/baetgB11dwZ8mtkOChcab3dsjwPtzujiG7Atz4An/l2qYMHuU/sD5H
L0PcjJCd5XSUxPsv3RHwgypfkukN6y2Pw9QdCWNIC8+CRbFaM4s+1X5LM5vQXKu8
KFaAQkN4RYoQ/ghUHZy71OScm3g6rZKzEyQDYQebHrYhIUKzCOuMVcSOHjiMwbiq
6Li0qDj7geE++ptQSkQnAr4EAtA2ezSg5ml2Z35GQDHpeCPvmW8y8/2eFYd+RhVi
WZD79yUdlJLCSEpf1o6mWm477etzKtaaRQHeJ39jzdMtgIOkVmLZ2QXiOa3UxZZP
VHLxUpmf9PtJXhvT3keXhNnqcod/xcQJFsUT6hH67nxPPq4j02gXF9EV9xRadYaG
7YocHFXpMc6PhxMSGfHlYOmRu2MDOHoEAOhKZMD4K9Aj8Jg4b5psnRQMx0AOAoAT
yWQHnrCshd1JqQgi4d8S1r0irfYge+HZCZtG3pQdxdeyD8fsOFgVU52tBNZktS1b
wUDowwCQt+mEQa3q6p1VkszGFpJ1JyZsrpxqnMAEi5HPaArHuw4sgabp93imt7vq
yGuVc9e+YxqAksNpD/OMRqZfuOOZLIarFfRTeAK7WUnWylJc5IMxfvE3CduYyKgP
LJCuKJ+M0qdV+fRqU3aLayxkT0V481fjlnaIUrtgZKcBNL+ksI+cJu/a0un8bOIv
BrLUh7yUmw9JLLu1SuyFMGRziLa4DW7AA0zN6NN7MMtOA3AlJQb9YfgUCqdH0KsP
cw5UeI+BbLNqInOnYVpw6npPr+hNi4CVnk5DG2C9m1ChXdxnKSwOBWFn/EQjIpxM
rlDy2xdrFL+i0LRo0/cug7t8sxeVq4k7RH57xt3frKcGVWo/R28lW1lg9ffsdKmX
LyPCllsJ8HNUNX2qLGEXTN6z1rolYoeWS5msH1XbGUx5HxB7lenBZVU5+/XLypbb
KXrA/x7vYnIj1a1UxaLXKh7EozhsKBZt/05W9AxcAalk1B3tdF4k0cdZE/XVTo8H
jvC60nfWNSfMXTgPmAJw2efMTU0f+ggilFlL0KnJocDtQnRUshFwe/jg/3CRgMJA
Vt8y9IUE3pWKqyfcNh/gPcjCRa0KpJ3wvf6WtGzt4b5ErxCBEBmS0OaNhuYSVqjF
cPTFxJS1O0t8g0MGDUiDVlW95jNBr9HX8quMMH4/fLtXqt8OGTNu162rTvMFxGQs
qAyqnslUhTYs8/fCS4Np+uVYykUVIpzj2sD5kgY6W1oD+JjTCHc+1aae0IjJRWDj
w9YGGRKy45JKCPTdF7Pq9D1ANPl9nQyMuybZOrVhsqB/UCJKdn0Mq4UvA7ZSWwRN
lc+gfbJ11NZ+dAKy/M5PCv5suDJuxsrNWSewsvU2npUKZaEkJ/TPg+uXvpQ2V9pv
VY8Ive8u12SRckuuNNlH4YxPqOf4jzIZtQ9CZJAkOrQrRA50JHalpsZ0ssHebsj3
VtCw41H0eja91N/7j8N/QhPi+wKtTlooJEhlvonX8mrexJQOOHcaHXH77gfa47vS
tWZa3OOjAEtuR+DQ1raQHVSqyrghIi5Z8VWpDCTM9wsOLnGa7LQQfqxFkBzIWiVF
JtyL5TiB+Ysm6ReJd27eayOWC5FDyGg9AdvGOYphJ7r1IU0mwqkabpQ06c6Sqx03
8CLUtC2D75k0G+x/5kSPwo7y7vCFbpBYezf5TzcABL5StmI0OHdG1edqTLYwIYoS
en+Ys3f+mtBguf+y71uZRP1okRxWE7+EXRxoA4PItmwfonKBXbMCxLxziyWJ4py7
Nuid5pOP9kWd5V83eDkF6YYVce7Sw5AKhmjJkgNf6d0N3CCYy2AQjgPKPnk7huvc
sszvJtyepKD7zX/jnmv/xvqroq9kSeD3BjNfiFaFBEfhFghmPw2QmdR2WDk9+pmf
mW6RXuUozW7vcmFrKhy0ztad+uJXEZgEf5QWuv9/olslCm3XT/1+c2k+ZiYe4Fa3
VRK9kIYLZOnKJRYkH90BbU6GUaAjuctovYIxvSDsbhM/PdsT3xStEkjjbL1h9o11
sbKd65o6YOzko1cgX+kg2Lli9++9n6v9rw3QCejy/iA0gjNJHojTL/HDsrcGHrL3
WXyWLa+CBJh3UO/ik4D2naSWI8wigsMiyGPAmhWcEZRQzB2QwX46j20Bgaa42p7s
gDoLmcN2TYopgJVd24dbZxSOVRwMtLJo80NqDxPX45dyktPoBqE18T1cMNi2Fdqy
oF49Fk7tkpEDZQSN9jddtvnPvM0ppWJQCHg+d5bVGwmY+mEDjWnSPpQLFL+NXyZ/
YnRo7hqN7S0+/aNB+93LDvMEw1VeYGmBp2vFCxLlaUrv3WRstvtLnxQEE70CtrTq
yit983xFwwXIZ494dFjWfTL9LsKA4czMwdm9MSTv/ZFw+9oQBk6VLCKZHZ2tX2X9
W9crAVIqNos/D60YN0mEXnWH8kw87jEAu1KIkHDj/qpFvmOfwdFBovkNmqZcASrK
cekWgEQFqPP5ryzMTcg/dAvmi3e6O6PN3iPIOcjIg9hBLkun9aMmxFAxQY6hbzZF
wMQeRoTzcpfAHMsNx++OBerWO8t8wbECQWGz48HVbhB6f83dpMjKuwayJV/hyhyC
iNPH+cE9b54NkUJNzQBQABPfh4mbWRCHDIj+TJPhy/3WIorkE6QHJbXKI0mjh44G
cyCR1YD9HA//Il+PC3Z+CF+vyTC/fOx9tCUB2LV0cJgW/Z4RixsMA0lPdeZ6bJzv
Ooyh4Kvrp10/aE9Q58JAWCcaXHzCalnpYG7zZZKDLn0vO7TSbgJQRewL78CA3pmJ
yfTbS/XfTsMMqckFiIm3U/WPsAT8kIcJ32e3QMTgDvwl7A4PO7VajoyuZAvqL4UB
/HBNgI1wddQGFKOy9mWCUejWaTc6xLcOb/3w2Ox9V77gVMwcUgtgosy7hcvrI8R7
htYmnzJUhIXL/ZeuJiXPMdslupBuq0oBvcZQKC4UdrHSWWHZTgJOg1bHav6jIQVH
pTfk2RrCWTEr9I8w2QwKl25vnVaAuP5N2OehRWGfx4TodVJz7Z7jrfvGaoHXDZWA
wAsaIstcsG4SljjroE88NQjymNsJ8pK+eYPofHwf5qjbN+be+rmMQp88EDAS4HtR
q2h+KQuwEY4AVLopP9zq5m5jtAaeY9Y1Hv8I0xtWk+TEpI6LSQ9SJpZ4roSffmFb
3ifNYyy7rgZUpMi7L2XS3+gwpMmEqlB0GS49xCiInebSxP8dUbtm+bC74UU2t5zW
9Uze0onuH5up7JhzFKDPiYQ7FJfoSbXD+WrI7IIEXVp57vfFSZybrJjWvu1Mf/1o
6uNf3fU8otqMVdSc+js5y0opTF51uiM3OEYD36OCgxM4fEadwGxnw4jWemtG5/gU
ewxQu0EjfIW1GPmizdfSv07Yibmt3GuwivnDR152pi1+sIGGekDpNws1KuHwKA/J
h4vLQOTPhbslWX6Z5aBqe3Mu2esBzMJ4kYPoF7I4ZpvHf03aj8R6MsjrsPzuPbnw
y/0HwYNN70C+8omDv9PpJuBJ2vNedjfKZA2S7Q/6vmreRzrf3YB8euymjTLTLli6
TICYkvNeq6zRaoB/bA10ckNzIrL1FPK5JDVYm3MkliaAseFkuuKxsoUvNmHTtAWd
W55CG+NMeLfAgY5839X7Iuh6gPsqu3ZnChfCuGfQ64QtarW9Yd+pkcbtG+4rhUTp
+RjW50IMg9tePJebakP2TyiT0EleK+K51LHjdlTnUMRl9BtddspLNM3Z2tq1zrQu
towl3mjW19BZO+D6Q6Co8j0w0pncQ6PzNQ57CVLBrjmR7VO1PxWEQtb/+IcufnrX
yC07qAeGwkjFiExJ27iVYOZhhCRhtdw61yfx0e7MnfYjQpJVa9Ev8fs6+ptgqxSJ
9ysmZ2RIKdBWpRPaycHzPZQlokd7KGI3FvKR1/xHex2KsHlbwcSh2VeSleVF2pbD
qvdx0FunAJ8oE5raiDzc8RfCmdRkIl7oPkh/vaQRfmoZmEKDibsuuVIdubTDC//3
Q4230369W2JnAmn08ycFbIbGEv9Myj+NXwEj8wX/fvNhxaTiTj8zCIQLt8/8eItU
6xKd8gISLHsRK7Yhm5cN89FXgXUA+Jk8JX42TecI6wBD8r9kiUO9XD6CtHMJENTH
6MSu1d51onaqeq5hgmKay6sHt/BHHfkVSOW9LlfYlOAddqzUuWfftjS5VBXAEgIr
b1dPHki0XC/iG8fMuuwJTrh1EYt4ZXk5sHCeko58EtTpR9bdKwMet4SO13eKct+I
7j9b1MlCIy54qvaTYfYE6ictMrZhJgk9ii5FdVt0X4BkZ6Q3gVLh2GBeXaWnSER1
x0MfycLqVrbPMVhSvyqUk+gFqzc+An3IuJokhf/Nvlj7Qjom22ya6cZgvu4mA5WV
VuBB9D+doPiAV2eTueBEOPwxAzIglP0+ZJqZodnbICY38QmhOOW4dNVLIY+YSayJ
m1GV6BLnGTM887GwQRAfxSmPTNl+CL4xMZ+KT/fpZ/F+rqWj/ksuCRd0kMWilU6k
b2y7XmswgY+jluQQ+qpm165oTkDdLRGuKf/diuRvYv//d76Vu9jwPhg052iVn4z4
5bUu1EisxM4QcwaXUhRkr1WS+FjjOL4CyYZ3gdTZSerSn459qJPmwkDRLlg+tFXz
W6jbI1NS6+t/ueQSjgA9i0TCJgrK6GJvV+2TWyZwYhllUCB6zj3e6ojC6I3pXEAP
7Hx2ngZQV3jZ9/giS9PhzCqaBLq0o3S6j+JOO0ABDcPsB0rcW4vk3oUZrOi4rO4p
3iQDEtpOmvLEilKtlx3DIaSTnngTzGuC9IBB0xFAAThXIbRmKQCeTxBsWsbA0F1R
ADzLPW6ojsXrjIZmkveD4Q7vMxe3D67fk/YMefA0na5pJQIh0sDl9idNQPcbQgci
a8fDtbSiaAvRi6//W6u0fyMvE3T2KZy+dsv+biarB/kqg2hyc/jYSvP5DZJ80tHW
aKUZuOYwenyEDcwNOCaiADYxKTD7C0UqTeCnvCS1/N1FE2Lip3kU/Yo4LL09ke76
KXmVtHHSebG0C92xscaW2te/r3P00oqvjGivrRaVP3BPyYmne5vVC4BTH8HMVJ4z
qqDc0H9UihsHSFmTx3jmTIsLNS6l8H4FL07/HDwfO8AVOS5qpJuDeTF1rAKXrkVG
J6WGOawnvIh3qDPDRv1u6JdNMdgUNbglgaGOPDaUY2CWDMnGv9bE85//qQaUPLB/
+KLVIPgkzJul/DA4VpxI5grkHauxMesWes5843sHYuO0ejJZj4XsO6T8HSzp0MlN
SJzPXbdaUUTIMNSJtO7Wwl5tSJyqBeu4W/Yii6M79BuZw5RTdMSqGOMOmo5+VMgP
yc2X+s8pSHYOmEDot/2/GK62gAcwH3fOCUx5Uv8x5Cs4Au5cV/dSR0w31ca9NUxi
lWEIxR5+QaTb+JPsh//HFQlwqzSgXXkvshSboMLzGVydfbh3HKwLoFZGtjGfWAfZ
GC1RXEKYHRfCRQbIsRci5sdxvqmZmZ/np2FK/W6SGRkfTnlcH4fECxgSTFaLq9dP
JYZbIXj82rneJMXzJk0nEex5yhaFf26Y02s1nWesQv5heHZy8/4KoVsbS/Gqb7A7
CN/nKWuSccLl2FONd15ae5jY2wRdd7qi6MY2uR5GD733j/af6gEmXeANbT7yMZrL
jOQN/v7gusg5fqsrkNPLv0jRNnKnunHJNYHNH0Vkz7QequRfjR+EPKbolhY6uBvF
xjpOFGbagyx1fkOne/DHHQpRs3x0J/bDsrRAilIGn/TiRYjHO8ugjHYS4nEdi697
B6chxJ9dhDke6H90omp6u9g6rs3xvZGVdMSWtZTGkKGIBqcVo8mwd/EPinwR6Vi2
TJujjnPtwx6KPT9lOnapkQyU3/h1RmdqZRfL5XseXEC6/azYjyUea0I13PA7NcON
go2bHaJQ15ITsC/koJBhbR8xFJ5QRxynNKoBcHjyT5bP6OMg8nRS8dS5lDdfzwqc
ixV/ttX5a/uii+1FqwBjKTOCDQim1W+aIzdLnwRgNqV6WJj+2InL9eNW6KaNFlzt
d6VAlFKaP5sFWcSNeHPq0nMoyvezVyaGhiPdfmIhIpyyxuKUAo0q3SQt6e6+qvAE
mw1Ds6EG41GhOPwyTpsCHrBSSyTYUD+eRFo1c12kHOrBbE9DJRFtRECoZVMlueFf
dNekyRcVJhebWryWj1I5vVGKMebgvDdyYEnUTXPu0R9ztaiOe1YGZyJQSbTodaHg
A+HESPPXVxaxYPQIcmF5sm1O2R7VN3Y5CScrz4aKqWX3GnQnXsdIRYCp71f9InZO
6mi6oAlojPL0VqSrFyv/JofRnYgmzrm0WCvs0kXn+sRL5Hs6lFVYZ15x+HhQkYSd
lgQvx7v1GgNPaL7SIC7HJXdCZadOEobAcTQjxrsBtmTUQC+l7KsGwYbzPWKQu6nN
WKSz5wTewKJDpXjlWT9q8SpYmev5tTxm1MaBPvBF2PY0eOu3Ue07FzoGA44yC19S
BCRGg8BzCEbo1+o4DbVpp5GM1iok1TJR1vRbhwXo6rpSzUlF7mbF8P5sFysKNorM
7E/SVteOXkpo/rCVOdu6pnyR0QGd8iSvN9ZmzZXXt6FV5Umvh8S1Bs7iIIKrGn8M
QwA7hjbZm+YXI8qOABNR96Ynk5vKue6LNU0KCMVKwr+Upf8WFxk7CN89F1/zbE3R
j6e3WA89dwW3Zf7lfzs17XehTozWjG4GRcXiQfTtdG4526qfDvYCAFXW4fyLO7V9
6aSGc96W0s60vRUKQ8Cah+rT43j5v6WgrWATEB37iEUuOezsVymdpq0BelCagYHq
s5D95nEs9ZozqJxMIi/TbOUdlMAgLqjhS1YrY4m6An0HJEApidvB9H3qCi//StDB
tdaXXOUfHmFYbW1KiNGYDlSIDFiXDtrkRcVTvw1Yi8+InIpfWKRQnzZpDxy49Axh
MTcWg1zjlLQAVkSIcpxLSXhujAi14nDSSj9FzzGn7Ju2HQfch0C9DIH+vttef/Tq
s2bC1bkdG9UQajDEIIwXIm6m2LG1CYHEBhVMGspVIaQ0oT1zej4dmHxtaqnySX/O
EStZ0L5wGxTS9iCTLQCZU93Xb/ljbk1790i0rq955MvUzHZBFL3r4Q35rxTtD1y3
ds192mscNm+UvJujqdzj808BF/F/i7gqFdjw4Y36WuyjQyj0aZJDBLTC9klAHNfu
tjwkEZjFLYdS7Vk3oLm7UqyHIE1XgNt+IDyI9e0kRZz9vDj+Hn5wo/tVYpYR4Er7
WJXcHCHUPkWlZUxAz7FXlX2ChEn8gW8FINXWgcSReWkxtTB1R3PS+fxYlFCg3efI
d4jvGbnJ/gLhm4Qk5oRZsdOlaTEO6Stpwu3U4XQIGdFDW2ykCr6086Wo85o+sUvo
iZ2Acn2kt0bKF3kLa8f8N6bpYXFZ0uJYb7Lu6KycZvsVPj0hBXI19egpVhrlpyhc
RLVe37zmj00ztPHnO1vSeXbqshJwx300KVdOAfRkHRU+JzH6BDEuk2DjFedVEi3c
uSn9KUfK/gtf9L1aU0nQemjJy32cwiNdqP/uwM20tT0qFElfmu75DWIYiYHtXThK
TyGZbBbU2v2psh8/9h8aHLyY4JdY7Khf9erCUNhKgroaQrGFDAsz3MXN/+zn1kbW
tua/0WE5E0RYgeS3fz8P3WX4wN5HfXu6gpZO9CTjgYaUOU6PZNqhBDXFYAUP1ggU
QTbuIW7YBmZLAv9G49wLyL3IkqFc/0VbKTDXJSX1N+G02pteKSpgYR3Spn9tdpJV
Bt0WZaBuf7kbhGT37yyrZ0UCJMWnCr6vYfodDy25rvfO2Baov+RoIODrJF1lwp9S
sEDtdRb/1Czwx8QUSpO++ILukizcyKtydmtkHBtlqTCKtnosH79xIwaUsy253nBq
3Z5s5EsaXlDS9aGSc0/rGC+5fMgr87SkCFPQsmB7nDklJid1H2nZrIFEToFJQsps
R7Ycy2wLow1wMUCGGxfJhvSc7x2ouNUsdRMuuxURvR4qmC4CzDk+HAJKNkZ+r/y5
UCxTGOzqsiWEYN6zv5s0Ep3+rLSOf8DdzUYY9zN0MbFZwapv4N5r2RehhEXuviOG
fnO7r/M4A/eUIZ0WGmHh8bvi+rKfOrAFyvQCzUIr+iwJVUa8SEFyKY7ckG35mIAo
cNwRr7usuSeLspPJdjPmUT5AGWHMNyYxsLRFlqoaQYJj7FsM8DB0+2Glgt+EMOWP
XfAHxtbywWsoz8hYx87OHpzWXt2omFrLJ+ZiGjkjPfA39Odck2xnrsRAlgi5b4a2
3o8mdjTQzPSaZkcW29edO+fyt/lE+vWf77hpi0U2T765tf0nUSSuv5VUZ6hcAxrb
erDxfufXgiFGZnUGJWwYEPFw9rrVZQecdJqHhHIXMrEpAXFm5Do1o1TNknzUBy5h
Kg59SB6leDMitelyrKTA5qbvKbiPkYNS5DMxDN/EiSHVGIaTeqPxjbqYzb/8r7ox
kbkOTCEIyboWuyGtEKO+lXYupBQwbbk5tUPwSwPw6jCmrcVZzMdcoCQLhtZHBgAi
k2GL+TjSO5cECCJ3G20WFXehIVRxPJbJ4bPr2pEoSx1nV+DpY0odEZ0EeGtLRQIG
KJ3YhO38Z4W7ZKnqFXbJLoB0yF7jsvSfoY4O6D43PkcAaSVToYBZmCnHfiFWS7uy
xEKpJcwaeysh4hubFMCaXIuSFIUsdbUj/AyhzYEMjT0mo7wF7JDQM+ZqU8+H3rnk
KF3vgrzyT9LjFhuh1NqJk6yx7D32UVyQqrMfwMKHbJoRtIko3U/ZVrUKW8X3Igr4
ptkLhdpENUFhH7RQxmvPE0hqt+on30wVVkoBVhgdaQF/Cr9mwghTYqSlOs6bW+kz
61aW/ieaaaOQz0/ewu6yBcyFn5+w+jh3cmcFaNJ0dwpeH5luQ5NFl2MOfP6j9vZK
n0OaOVK6I9Zp3a8vxtz4dONW69L9JPuaVXIvwhY/39Jospgl3KeKYG3Q8zqDGpdI
IwfaE1jF3jcCFwrxYKYhukWQb82y0mQiFbC8SaEmfAA3DX3r8a85mTLaPe/r93i1
CMquNZ2vPabSwo6lWhHfh2YC5kvvQaZk1en8aOnMVXieiBo40z4WSnonDGA73O+Y
zTsH7X8qZMFcPxTTFiyUQ6qActwCQTxkWkBO/LuDdfU5p9J56chD4KJpAEvMimSL
TW3tvL/LD12P9q20JdvFzzIMSB2DjPKmozaJasNfV1u//mrZiaPn4NCw0WRJQ16T
PE7CVzLdgAZqDn1FLsi24Tn6Hv1GTeHJJBdimbnxnsjGTXo48AKtQi7GSXY4xTuw
jQDVFTSeH4zDF+VTWMSmaAnYYy8oWFTRPMU4j511OW2i6dJQrkZmz1PYJ3O5cvu8
K8VX0IpGsf6b06lcqKPVE8pn04OC7oYJZE4RIWLCQOI8Q6d7FsTM0qB0CZs6CbYk
MfKpqtf+GtXc2GyIAynFx79yrtpjnobX9mConiCMvmZBY83FjoC3o6xiJVdz9T6z
L8/ZTlQ5PDX8VgO/wwFsn6RVEnZ9rdY03/oLUOOpV9e0oUcj/UH6kuRsUqVf2Bzf
lliZyOH5vESN4AFCUsYQ45M5LSq/1npCVumTaPpNhXA0ntfK81YHCRTunUgrfBBk
9lNCpKWBybxs5DnBfp9vapOyohVectqDXOaqvD5eVJqMOlhW9+LymBDQeJuosXMa
ba3X9OmJxdomvQCXMc6nSFzSrIrAhEiUgUyFq047CtWqkucjblBCNj3D1fk3WySd
orIVi4w6GvUrKt2fdPKjU7wzzPkmsMAVsJdpPAZrfjQi8LD1huNfDiMQ+9M/S/GI
oviT6wr9QwGFD2ILZn1LCPUTdqKHLmelyWjM2cAN37/39EV1M4CHFLIdXsNiZGzM
BMtUvC8d3y5pggS57s3/Xre0A7Os7/QHtzR6sJACZKYJ0GwHgwcnUlK7tuvxtVsx
3e59A8kdFEFQ4z0wksfvqKkc0EJs7bMDGxBzK4vfoR4uiYsx24NvxM91i89K9gbK
CZoy1Ipo6f7VcIbJj6oaCBvv9Mu4mFd5PAdf8aFN/CFcWDOEB0yG8iN1LgL6z9JN
fmrlXMNHB1FHiQFYBWZ6sfYpXEu/NI9A5mME8Wz6+mqYrY7doXOoT/Z92iBYrklo
6t6Slu3GcQ3xs9oolTpLgJ4sxPY2mv8ALo5HPg3WvEopRHyKqZSBAfXBuTP2vdqp
x9tzSlabyWLazMxclGRavXrHO1c5rp4L6Nhs8mFU8durNILKOPkz0fMgphWfKk6m
Aqw4+n6eyeC31E/J7aM1xHEG2y9RxuH5PhAnj+FFIdumednCmNzNqu6mSOUidZnF
tPwv7+dfhnl5c62hlqRVuoyysO4APabTiRXJB5CRWmlUuCmjY4CVVFBBkaL90lvz
rrX/wHwyrQ83Y3rTVr39jj5F7THZCFy9wg6t0FEUhvq2+S/RJtr4+ivX/hHFzpD+
cYogDv4YML0YsMYRgCiaTs8ujQqw1sz2DkPoX1LS40zENTE9zom5JtMXvnSQeNBT
DMRdstDMMW2FKcJpFl0FsFnR/SLsdEVQ7k1hzZdLWDOZlfsFPgujJfKRsq6Pe/Cx
ytsohJ/xBL0KKKDQid73M5F3Ll6O5186sgiN51K3k4MAZFH5rC2x/we3HuARXvaC
Kz/UttbQSJet/ZzIv9rGMIEa5BM+LQ6IGpULnhhTVmosghDzKijHBIGN6Qd0vEWJ
C03iKXwlvyvAYEBDXmjyHSsnAHVSenuXX2tkiyofbKVZrg15QRYM0TEuHerJ1zas
x50/BvuDmjvVXutKhYW8fhidwfILFokWkPYi4i/eFQaGFDnVOIwOPGOkV11qRyHv
4qGwNvdqvVldf+Pxzn7tEbukUGgACWl+UoZ+9do1H8LU7BSVq2x6qOAqUSvR9qvC
cqQQzWsACWb4DOtG2zdxkjNLW7JJnRzhxYl9slhlyam+f4voU44UUSkUYBHRIrVe
psesoQ7DZnCrf39OL7BaZke/5J6slrWzDK88a4Y+q3ubhyWJ08p6gqcirkFnJk2J
0ZTr2Ai0MW1f2VFNZOx9jerfacXK8R7EZFv3lFDn9NBK8Dq3TAndZgvRbJWqyzjh
EGdXwPx8nXO7Ugz5omPFopOsSmUQMAhwAYf/tcNGjCKzWs6Aq955Vbqze+Ymf1Fd
G8u2yB3+LoqTQesnjyPMLTNKZue/qm9FE4aBhx/q06gPOncExM+Ui7qo0i732LsS
Oy4txF2AxNS6Wp+15hL3C5x49P1yH7YGgw92VI3e54cWqz4ofh40D18lCOxGwPiB
/xNcdoQ0U3FbYHMzqyngdgmOoJenGUlJVYEZcdk6DSj0bLMdHb7Tvu3U2S8XefaU
+IBd++O2P1PX0/25x7nkdbB4D1yfGLCXidvmgyn2uVSHic9L9VEC192uskLT01LE
G9o5qTLuCvhp9kYOJn551ZTSVn+NAeHRfqgEfbjnSubhAUxRDsQDiW0QgZ3kIaUI
9OYMlosKYl9FTIMYWEQP6TGimZeSiSr+rTG9wpmbp/ys3dxX2uxb1271eB4xTWlN
H8VtB2gyrA2Ez0c8k79ytgB2ZGzcPmOD620dMEA1t7PCHL3r488BKQSCDUyLzKAE
N6gSaFRYyZPmeNO5RYIDN27S0ErFQF3sJcJrdOCQPQx1fBbKJ+cgcFkXZSyBC/Is
PZK4Zemlsn2NqidFh2VgM9zRUq3ewAHrJidYzVPA4EGgTNSeY5/tSZUMFZvS+qIz
0eMzvS+6U/nth55dKc95ThIC0Nb9gi6NwGVm87ncloXQtz3MHRKHiljPrPem6cNS
F6micuROB4rvGfuAuD81tOa/n7e/283PiJcIC5Aj838+sDtRntwsipGzGDDUCAOd
HIDYSUUzlj6GyPUZAhg9GKtOXDyTQoAb5WjQI4LJkckFI5jO6fYcqnYSlF8d7J+b
UQSQ+FG9wZVbLCdHRd8FJgEjtigHSWKgC0j141iBre+Cfb6YhorXKKk+2t+lUpNW
Chfkutz3ouYpoA+zNkx6Tnn31WjWeEtqAOpm5aP3mnwug8OVwQfqkdEaGNge2k+b
yDt4qJstBQ7x0V25e/FSi7sD90MKJzdJJRzAGKz6pjVhSHz5BRJyXf162uFaiKKu
L6H8A+S0iAV90mObBMiPFNwKx/6m/3ihGRp0xIvf0dXVloANf2g/iSq9kQ61ZIyJ
Jr+P6Zb4Cq6D7ZfjeimtuKEKS7NYX6AxBwGPFJYADx2AtqzP99UaQUKXWdi1uv3k
wI0IuJUfRSIZumletBZVec4k5FuUfy9/KlUIb6qEqvYfQwk02zEAGZarg4kGUDRt
LKnd1TrPBzoccHYRQw28CpVZr9nlkyDjV9t9vlqmekfN0y7IOQ5AwgQ8Fz7mUDqP
7npg2PBtn3p/FPkWUw5N6n+UMhsVDOnvsvoZI2awy6/UPnADVkF5tHj6Ysuid6VC
ULYxI2+xZqgAc7qp53SApmGzg4hDMCn9R+W5/xV6xzufS4lVPG0rPNV/bw39LtZ7
fkHu1fiYaIdiQYS0PC+HVli/9Q+f1Lq02wnF+85oJqGFKsIQd/pY0OyZMOYRNKXW
dy1CXJQKFKNdsw+yFJwnaDFiEUoe5zod6S+SPPI3WRHE63yfsjcOvEuzlLzpZtB9
jkBWzqf9x3m0v22aGlN9UMHz92NaBFc3RHXvAxllKzsW8Picixb9FUfM9/SQPopR
WxnDedj+c7zeHal9Wvj8mZN7BtAVpumPqKeOMb0sF6WS0F4IDxSXNBzzWxEIHWhR
1p7vcubCOJDJgYTeVaXV99WIzhpMMXCAznsBO0xypNC2qAA73ccMwHMl9dnD+08n
/+/SN/3kNzuJAR9mq50K6wWeBtIlPPZ5Qriq4/C6dY+UGm9zPaF3T+k7Ak+YPhyD
Zlc5l3B713WNUJGSKaeICk4Agb0lQCZ00Dr8UT2rFcQ9kGjUi7jIneajxeqQL2Of
Ln0EI6fm6ZImyDJ+8CWzXrGU8HX3vl46a+heJTfahO2gozosrCh2x4AvMVGN5pix
ugGQxBb9kiSqMvsKUIKbUOCJJYC8ZEGonZBnr6Y+jICqii/uW+UVPzpbYRrulcxm
4no98wCkOQQhSLpmAYxD0o+QP42bX9WOkXVGYb4nK9PpDq4Fpuk4xQN0g8RsooCp
7WgBdZ97mgOXNUTfkXvTEXVbGvkjFPF8l64PsZM17r+M4Nt1IVhWir62S4BT0RUc
+Ktod7pIrQIfUy05N1tFFqxAR6zYfPxwXF+pr0V/8DXSMcz/IcBk+lranmPe9cyH
Xfzmn4+B4Z4EPaw0DWB8MEHW74L84hbSzSXKHfbEvURaXdsyCT8gQB5zdBCLHRLQ
NDbv3N8P7jOdgtj6TlU9aeQH3ZW/WfuZU2yyjp3RJ3m4f9emYLKnpsMNwhJ2EVDH
N0OQYaxcY03U8Bxqq2AMLqhRWFW9P89TORq97wEMZ1XBQQQMSwXqnBbh3kyw0z8h
WbA0iWsab6X5dXNM00bh/lNdhawqNwHI/iDv2wz6EqW/otUTTaGPrLJT8IXuEGcO
B9FxXkXHUWPxn36Zwvn4B0xgeYrrPOi0R9GBW7EkcJv+BQ6fIU+anJcG86H3ew3c
p8oKh56DHr77zhx0gc79dN7zJvBxXJR/ppAMSnUtBBCg+M9LYJdfqvqG2Uk/KfjV
x4xO1KREj9IKFcb5W/MqwcTDbnmfi7EYsQt62sXI5cEgUaqlz10p4WRlih8w5Ojh
KMpEqTEpJfHSkokpG/oI3Vl3Zce1dsssbQng+dQJx8Ms1k+IpPDAu0EjM3ISNzX3
AsdFQyMwUISA2xYTDURoppD85vvwbKYE3mz6u+HcdO2V9s1cZhZXfXOnGMnKtt4M
GYzPE89BkuBLS893mVfqukseg1fFMWpd6zFaFwmY06X0GDuK3pvS0vtwHegdSC2P
/quCMPr0ZU7t5+1JzCukl8SDcz42oOZRH8tEx7+IfwppXT9AXR2sdWpa3ChOBvuS
E4D2H2S+wy8Ep9j+Oym7CTVlPD9FR7dP3LQnvpe4Q7JlLzOXPOhLIgGzFOIlaUkd
Whl3I4VnlBQ1dlRp5OXHk5c/kzQ44vKz5CW+ien3ubbeSKijQPzECTrbt1xdAAzB
4eaCdZQlT5OP4MKCzdoFaXR9BOU/VoemlRfvpOSgzSQW9bQqq9ke/Y9/mWxkuhCh
bC2zJhLkpSnSMiyHVQ/0fJUxRfPF/5ETG1PmP4mjdy5Zt5/iUHF2f1anmbtbOYv6
AsBcfySNXwUEyXn5sX3vrEGlxq7NWkwgmjsr14SM+XFpKz1m3pvUvZkUAppbpY4l
52cK5d72Ilc+m+1VDpSoMTvTq8ld9kJB1uQikhG0GED8cO/lFg26To/lNQxaw1nT
ykBpHVh4RLNWoxYsDh8/LjAFW2K/9AONWLtU52HmDe+Vh2DixrYu8SlvXdFPJIr6
glbKaaYaGFXXNrlaTAszGaHILcIARLEXIHejx2ZQVztp0SO9a3VIyw2llUXuD+3U
EHstyCu9eEMb/eYRk4Wa2nShkhbwqAI+J6d/cTDi/HIuoRf13BuG5DNtgqtuPbha
lgpmI0vI8zmWlURN0xX5kaifM6lcjfgLI2xUiLQm7ctDnYqOAmX2weOety3QbHWe
JYgC+vvjZWjOdG5C5WHnzjGWxVsKvQKGhCwOq3MSLqoJV8Fp1fIFnGGYVib/ju82
kjPpNQK3X14IyifNjKQOm3Ho6KD09FMeHeLatt4gVYiFjvKwePoqeV9ljRTMixc6
IJhzONX14yXTuhhIBmwBjqr8y49ufh+XATNHzSZVS/sYLVFAKr28Fspry4JXnlTP
SwzqpOOhsia62tDCsthmWSgy0JD//IuVyHXbngDZ+8b+ssUu95SIBu54vPMILl0g
+xj4xLWPvvA0uM+73BIzxjl33aF02XdKDDTEPHLEwM+iC/w0qyE3KkMyZ6edatW+
3easzU6atKa78fdzAFJ1AS0my/ucUJhu5P6U8i0L1fWYnPt6Q79UuYfKxd78J5ED
rT/6hPQkS8J0jOzp67qRywWvw1lAARjossaF4IoyTIvAH7pnegXgknnL8w+CY2/l
M0rXUCxHwyDO0YFsKA9pJUTeCi5U6xb/mgSIb5gl1bdAaClO5BVEzmEviIUs4gcT
XZeWwrUWu66rIeFFPk0KwqyC6VpOZeU2YiUpWLg/ucUj4YJzA9GTa5UYYYPLmFdp
oNAJ10dOFbs9VJBoUi5gVfpUkkWtYGkYmCkMkcmrlboTDQKEeuEwS6JwmOpsMpMm
290Ug3UOQu9IOO06NDQM9J6KQIMOMcWOimNUagxun1qkTGq0wYeuKZvglRXtdLhE
F7Eh1mmAen1AVf5UuSlh//ZfH6YyDLYh2I2PzzbS/aCqrUsmNLk65cnUAa99Zrpk
SwJxpsTs8SjUW9VE0sdPjjyvhNNLe7A+/DJgk47QZoYEM9xBXPtz4Dws6XhvJWUt
O7hyEozfebFzzfBhbIv6OG44kClvzPJeslSGlKBXoP3kQzfVMp8cuN/rPlDv1USA
6IhUnvpWoYabunhOX/iP0WPlhF0YSx6MmbW5ruaCOXEevnbfom3snusMaUS7UOwS
Y3kJLpOA+V07vXhlxsv0Em46k7MGY4Co4bDDMLwE9j/0USAUec9t47oXk4Pt0Ux2
sF79chzrA3cAcdbn89URw5pldAVphqVBHmNuNgLkApBsMIbokOLXaaM3thKpX9kR
d4HKZkWIxqcTwSaj35TcdxV26cX64Ju/ZTiA0NRgbk+giQVBjBb/9Y3aUiEqRKtw
JsV7yP34zQ6zBxo37u/Dy+jrIyclPKfi9fnEV+8QKQCOXG5JER7amuAd2CZLH4fM
PZI72BJiWSyAGlFYAQPpQzgPa6UBVvkr8qUbtKxRUAspRhShahQWgqHC67G6ipch
GPYOjSxJ5uuGnsw7m/Izes7YQmeoz96wk71AP6kgTDIxbuC2pumme2t+Dwq2cpl1
6sGUYmVPh6486xmOX1Ns3od++vcXf0TJXV0HBpi/XBTS1FZYpQMc/H0xhu2EiUEf
gZznUv8PuiaTG3Zy8kA08TsBKZqfQ3ln0xDpDF+r3wco9wH2IGBaVL/otpYWjYnV
oCeR5+C9l9TP1PGhjifs2Srmhr5kmpQrSG4pS/zDEwlqsWfsXISYOjhXi96eszFu
7y3/RFTu5H2pg2befU/3uO3ATHQ1rmqsXke00UZTfyvTYnQKCNUx6CaKHbFyg+gG
753nR8XmDZeIcxX/p1bCf4LZcOpIrB6n3w5CDtCyVEIOVDAV6VgVULeH1J13cZrX
S6u1WWuFy0KqajOPKjcu/PO5aPxKvpXVQYR++bidelxFaj+8XiPUpDAU1E2Eravn
L5+Px56ne3CXOEJUGit5aYihC5Z+OjSYnKYnLxhlJBMvZZuornC0ZVBL3QJkJifj
1bbdIRKxLfkAl5aeH8ISjc7RZocvCrTIgFCCwT9RoFTNO6Sq1cnmIHMtbZLVJcMM
s0mhaSSzUvBDOVYwpqrsN5XrIzPKmTU12FuGauA+nMEk+1c+WE5TCU2BjGFPM1eY
EJ5y0zN/Ja4brdYqlQAXuL1K1HJspB8MMev7s+/NjCuCzmAIN9RnRxIkmrFTv3HK
UYXpgNq3BVdelb0jmrc8FDbnZ9OZZG4689Qh/pOpGSaHvFEkjLMxV7DfF3PXyp+O
VSe3Fm8Nz8RrW7LUE8hdk7FDP3Cxjef6/gR+xAuBHGtTtet7AKkuGKuuz92aGyMZ
LiBv2c5/pet67mwc/efDBe4j2m1yDxsO/Nx6WHJKj99djVoJsFI5DZ1mUtMoidY5
msM5lsjaoGE+tnKxdYdBv7E8/qOuZOUOq/PQFVPlG2zPCFfrDrIVmaId+PWT92pQ
Sp6ubEmdpflT1VMWo8BHOSV2yEwFJuGUxPgh0Kdt+RqXoCKjNmpWqOEUYRBz8Pnv
ypYkX765tUpY1Mev9L16+E7VN/YEHSp27nit8if+roaswiCTtldgpTHWGbjUPCt8
zpRqYJAG8CiXGVd86in+JNXnT2FN1lRitMXA153uL/dqo82jvtfiMIkYexP3862D
731t+kXHl59dpZ78WvPDSfjdnjtYUr2dREG7jdzgoeSAtya91FJDTQqMxCICJyCs
o5pzv/BoUvVva4AdqHN/tUNRMS8uxTWhDhmo0TW47VvihvpRBgRtEKNKpCosb7Pz
xnDtXgLW9NC2/nGxDrnHrNHCvferyo8zAcm23KWhNrnI2vBr9/rAFt5dKnsHqXr7
5JWLP1Pq+H5KqmbYTOHyHmG8akr2QJCSItXD1EMHnXtJoDe7Ys/Gih3EN5CjBNn+
17CNPsZ0S8JIgiUGGFF3cg9dPlMgFmfwjtvBo0n7IIWiAxkj4422bPwsikHK4+BA
2hbPWqSgxt/jlq9JqYQIr7YQQo9XWXnzmmXpPVq7gD/K5ylPmcto0HndCIDt4KkD
aiwb+g3CeMAY0UqP4lnUDFunRL7erMyQZss7dpHwux8I+Nn8Gy9+ekqS1Jj2gorN
ox9br/W0RwfC/ToS/tE1dYBP5uoGOOdKUSMaPeO2NceXfNGlz0ptF1ChSZ/tz978
rgjF/0lt46BljSmv7FulEmZlBiCulW9nlH34u9L1hg+WjdGa6T15DvYgKMHrtZQm
CY22mbS5hlWtjhO7WoPhN+H8nn5BbUgijRN6kgWJEp9dBPqd2yK1Y9J9ucem1CmZ
f3zi121GmmAkNyDzdGn6w0dyyV9CV4tQBUsoNASM8V1Bu//7ExO4kxhdBy1aDcOJ
fxZdmf9d/npeNy8V5fGe1ddTfCqbpjbgPY7zm+P6OInvBb3VBw444Zdhcs17e50W
KAXlgpoRYFGXBdeJswC++0685idvxJjVn2AWi9w8G8AT9FqPGXPcG47s+SAAMFXC
S0ChTdTTcyWyKab3pEXGry8BBjAJPxDWxZcx3ixCb8oFlfNrblIUEQTSvRahuq5u
Rw28ZlHw5qAcC11hQyy2kBsK95emfxLTGUvMcpOJ7u0Gjc4Q93rJDnQ4/FNnpmyJ
KqJJwuuRLGgcAaKENn9XX7R4cZX6jIEzpFNrS3/sliW54gvBUPDSzwnUvh4auuWB
SISm+DzyHfqIVjFfxZuCdYfjdGiUvGLIPhjis5C2p/p+jBzbK2PrIPDFw9BeyoOS
eqoPd13yM9qtHswtzn8af/c+rPZwurPS7190QcUHU22pfEl/bHqziF5tGt6cKatW
WDHNirhi1/gJba7LDrTQ4eYl48v7tN0+TzcxdVn2SfDQu7mtZctU63zJV5TXIpKj
7WzzrjqnTgWtEm44f6v/MFX80pnN8rmVDS99rp701fxrPpy31X8MGvj+gdw3kSVy
HgkpSRyCr4EGkLAepTl2dULxH2W+BDXk9FnsMleoZGpfqR0fGQEC3Em/L//qcTnC
23TqPSDn0izmWdGIdH1urI9W8r3mOUVXhfNwadopcqCQw4nyB03qpHJZa7N1lwcs
9DM2+UbQcmwnbboVSXgUB9wKdgVCfvhBXgcajwZ+4ixC/X/qzweVMJOKD2hTfcGD
4FPiRL1P3+8MRuD00U/bwAHwIvPhRScnrDWyp8qE/bjxcv/Rm4QS90J5w4pPoy1f
d38yMI9iJpSq9e0JN1DgNMZvgxCQvzjRHoGAQcWGpk2iuBNd9nlSTopStuLHX/XL
OXaR/KQzzGhZ8C+kY5QmQRaKwNl76Vgp4ginSeDLW8CQ4/qw+vKZSahXuec2/jM3
rBjy7rsdBAxZC+or/qQ3cfOZnok62d5k5Vcu5O6ojnqMt79URk4RDctm36/nw+R8
GTzIB2DdHI6J6PI4P0ROL39rC7WKVgAYfecbMRYP9N0x/n9QuHM9fspyWJ/129FL
zrf8RKrNdntZ9RqIWqwH2LvwXiR2zAEz1YkvVQR/iXfsL5OItW7oWDNu2z6/m45D
By1hPFQuQ/e+sDVk8IueR2SYw0D6cioaiQc0Iks4Z/ibxEE2kdqRQoef/S2j/xkA
1pq5EsH3OPz7lo+Ffco4e5hvTNp9KmSY609UT5dAz0MEF68KIfhmTtWp380SaqPE
9Bdwq7/7L+HxI2s63YHFC8kwm5ljXOm4gyJtsADTsATaiRDY8F/AvVrzl7R5Wecw
rqJhT/Vb/xj3CIZLXSkoa04lmWAz87gcJG+9dkCU1mxxBhUSqIn4B3zlrUYg1ZZx
YBEqXM/2V/ZBQJvSRD7PnNNcSW/W5ucwY3ZQCSfa2vecOXEWPZKQj93pN4PNysip
I5droHWHfmgzN1LzAEclI1UERUov1k9ALztMjlkb+VzhprkiMAXjNokeybd7HSuX
8NBheJ3q1NPXVjD7SB4VjGSRemd+BMCotJ+Fg97FrefDMx6w0eUxdM1ZLaO+ue3q
eJri26o0wsVRalQOtSZJ/BF8GzaULtiv0rjL91zz1ki8n7yywEjILUIL3cVOuNEu
uBfXJFdkAKBwWYBvYdgaUTKLcoV6Pr0TyTbLKwlvMCW9nojU1gfzP6uf32gw2ezE
M8oTfcy4HK53IpmaA8aArwk9P5dPikcTtmwhyOrVvhpkWYeQjUpy+quxh3ADrKUf
D5eOqY/x+xHmDN4aciSyft7LWEd8MFvXbEZVy4v1Zyrdl5jvSqcj5W3eP1SLRTyo
s/Zm2N64cHrm/ImaLt6QHYGGX6sFOzSTioTjIBKDgmW4bx1je2LldNjs+U/yh7qc
KAOBBxSsa7UjUwvA1Omw+ZPDQV5wZtq5GBCJ/W+2RYXqUvNDI0BrxeZa6lwsPrW/
kqA2rbMeDhpcv7ZT9Qtq9ttEwW6Pab4Jwyy3BsHMKpfCpSMtH8xk9kRX0vuOiwW4
vHMd4B4rROppLc7DHQzPjOBfkzuI/Jspbv0Y/Vz6dx1fxCVdXvDlOni8c9Q/sroa
zEu7Bkxa6xl7CunNdN7QjShVeBDnDvPFQooksACnA+o0tnjleyg6kDDynCFB/Bex
x+jcD/EYElBmPTO/KdXa7rhXL1YEWxMEwaXCDAiV/5V2NHMPv4zdKc5S7srioSil
52eYwrS6xw8WcZgd7Lv92YdK5hKO5JOWgbFT2IKXM5/k+Q/qiO78OqGOc84vNghU
8iFYgeAcTH2Ghhbedf1fKmCG3UnO+5J6Z+nNuhwuvfrj/KI3NgZfjhirZa8aFcIt
mchNDKXfUC3W3lYqE6CQUYsk7LG/YLqSfENSxf+a11ET/HVnxK8+FDqSo8ahp27P
1EDO5FUe73KJofkGO6WG8T+TIEC4c8KXepCM1KGygZObkJtYfrOpnrGZc5S/c3PR
2QeG0MG4tZcWRI3LpKMQmIiWf/oq7WvtQoeyi08o8eGE6LJ9YrQf6On4CCjQdLrV
9/zoyxeFfnofRL1l6qvt4I8vYU0EJdfKsFHMgh+TYpFNgrwe1QyP/rCjbKB/iwxW
LWx23K0q0dHWKwTgj/cUQqmhLGiTIqGz4nKGIUEYDA3xBDdzM/JtNCnalwqG8tLT
7/HwOPZRNQL4hLD5uvBD4Uxxzdi9Ofv+ZpUYSGLSLXAmgx6KudJX23Uv23SFHxRo
fII7krgnRLnB8oWzuAsK+rl3W0mkv7GFd1wUX20DvtB+jW9CBinse61B0kkGpuEg
Sq+Z1zxM70S+6aGGvIE4kaACJ3cg+i4e7/8R6Gdnj2OgGNnlSShXDZdIjd9jvEcH
8MzIrURvRNaatVsN60XbuFHFs1eDYH/BbE50oad7FnC2w6h0elKxEMFdC1uWe3AW
WXrqFTtGGwoZ5BHIoXPffIYlfGy4RDmTabu13VEG8YHufXSHEXeV9eD6WdrcbgDA
EEKnpsxJpcHSO65eVKGXEMCQ+DKxxV0xNogxY4FA93/Dxk6zqb65QVpm/IYxL4FZ
/QhshsYLapE915Y08f7mLmhyJmqgtqxigtqm2hZ0Svy4odew3bfkGtWjEym9eLYM
hqUcB19A4/561mlT8BmXV7XQNb/AM/ddXdcvvMn8aKIj17kYu0v90yWwicZ4/Jcu
EXJKZYzDw7Zs5lgH0A4E8N55g5iZTYexMn6KzvJS/f30rzwecys6YbULnW1E5ruT
hqqF/mY7iO+aLjZZamye3dqEBnjw7z4qeUBgkfA4a1wvrt/+dHVS2Yzd7GXvfwgX
hmAFG0ko2ba3tzMQocE0158OxvQBN1RicVMqFQSyZH7ScWTYIi41YKsoPpmCaZtG
G7C6xWxtCSBd7x4TBLVeFBbNPZRL1iWtjquXTr/hk0Vw5Rof7MY/fsQJ4V6Z6oyO
dsVKrYd1rhxUoJ7wZFXxOjrJEYlHm5u44ooUmunHSj88UBI4Z6ny0P5GQr/O2kj2
E+/2SkOvV5nUNxd/CfukdvY9d2n9oncSINdZcFN9uFZh4cnSttT4KYxAwQtIuZ8Q
qXTbusToESe3gyvuOhlWqqW8sTcTGfZPqzgSkHcfgRncaNYzrOancnBmvn1JKriE
/sip8HP2W0ubPLFcCJKZ7zwmPylNt5HRx6l9vyjEDS6wxIe7F6FYeM6DCJjNgqVX
bK441Wez8A2tkYRJgREL6PPA/KQQAoVRj+fiIrz4M8kcmz6+1PpP4C+IRXkiGC6R
0dDuZH3eLE7Q1qAHrX8nJR1RNdLSvQPVOnS5UD9P7DMsEgLDudqBASSdR92LNj21
BkSnQB4DJE7dJab2ZfixKvRUw76Zto6rcaFcJ48sW2sBDahpE2IZ1DF6loQ36o+G
EiaVnpbh7wfbGLSxvroWn9GWaFylTKbxavR45JuvZs93NVWQYf7/915PL6aRQKPK
2cU0U9rjN0EhIR2CmMbKH5cOwI/uP8uBtS7FDDoSUO2ofrg8NseBThpk5lE5vZTX
AhU+fbWXayPoJRlVxryb9baRKzpLRXQVv5G5XrWVpyD1QSW2YS9RCl9X07hXalkH
0HG2MGujjx9d0j7pMssNwHdZahvCTKpswwZjrME51X2MKmAwBymQ63PFQNwIJzDr
tfxmVBG2JSTCRrY57Qdhhu/L9NgAjeAXC6qupIhUfSkBZjlnBv+RVoN+zBJQlMM/
GXVNfk/opUO/w5MQ4v2lE3JwlJ5giVF+XBptpxcU3GQL6BmWwdvqXM7lY7x+bq19
LloZTkASWa2PBhNNZrBhLaBv8C6T2aanrYI2h+zcfa/39LW4zJtIVJnC4k2fucUx
ebI4CMXQBURgScOeVAAuhq0PGlFZILuFomRG5LAD1Z5QMU3A8lnK93+cr3bQh5c4
WYYi1iMPeb5OY+jszd/yKrrjtEbeMqqs3Lw8e9YkvO12+mSjM3bm68q/FTcrgoow
2U/JeN3d8VC0dl6+0NguSSpZEnMpTEDk/mzlikjYptXxEpyxywd+xhfkSvHfVME0
SC2+M+3CcpRkljwmPyHcKQI1yVEoBe5U3YXXgP7T0vcWokrhwkmgFZZDk0KgGJHL
Nwx/Pc5DJDHoCy/JucznHOXLqV5oqWOBseWQcXzqiN4SW4/Yt6tvj8MVZz1MKt6n
FPYnZ5qkBDNXxXoP21jEbNJfv2yxpQH0Y5CmQt04PvLdSSdoVCaDiFTH6SJdB7ad
Kfjeg9Rj1W6uBNKkwKrgaoFqmoHeioUZ5X+zKjQ9Q7zryKV/NpErLaxP+9/BE9Wv
wPRy8pyi9+HIqNew9v6hVDQ87G7uCWioBpocE0BuNk2RGYfYuXsN4GxMCv8hBJxg
uyMe/b9WpDHN5+Lr4HJelSViQLmBXdrtWJKQZ9V+3e3RDb9jK7QV06fib3Hn/mTG
PPr9cmXCVLbmdA3TREiQyHGqILoOs4WkmBfL6D3cjSEUYhGO0EkJNET9Swjufoq+
/JOdOLe2TlAIBmDBEHXoZyAWyC8YlA4e01Xay2MPI2VBKUI+pO8Jr20hjrr2ROoO
pjYOCnvdVVwcTAMc4sj/5u53LOZRoXZpplFA+T/W/2S7Xx1rbyNCunOVlTwCFJaV
2v1ehBSZw+WHqAMJfLjTHQ2QCFWL+iW1LtC107FufCn6rCZ4gfl0MxcTw+Qj77Zh
zmrFv553hrbQpiPFy/hd90Tic/UASKXXNnJM+XKL+4olZ80TQ40SdbaD3PrdlwVR
moJKz6BWDjcuP86jXZ2iM7x5Dp2dqxuTqXcxf5zk23PA5aFLWIaFp3Of7I/P25TW
YT/269EVLG46TtzqMH0333Xqszzt6bx5N3mMg523OFl95WaIz2zg9UAye+y6djEa
8OqqSPC4046XCz7Zj5/RlR132sDYHMNRcy8hCYFfeOS3FKnxSb9LvhdvMr56ujRq
IQDM5CUm5WZBv+IlgpP8xX7iiQJ3vKR4JMTFK0KzF0LEwVZK8Jv3vhlV64JBbD+c
FyiMkwGpMvQd8GDvVCQgI1piwxQKNt3l4uy8IDa4S+ZQJ6cKiRmZ4i4lkOI8pQjf
EE3EN4d9LMH08UubIaDIUtB5x5kbkOudBUNDqRAEjQgc87QhfEbqk35lDxxj0MJn
1za5Iisqqrr9u1j4OO7ZRoM4Xf7aGbpO2HhvZRWCRSD9nftoTmngqxlSJFupNO6q
vlhl9JGumSxpdprKYzzj4fBxpBemfEnnbqajyqpJThK9v9P/eVBZc2zvcKGv6JkJ
7tTAxrL1HKJohnAtc2ZiyMsY5eCUUKRTJFUwSNhMFGzi4xNxF8uwJaEdYikSIBZ8
BvQoN+mV8Nnr/ro0CrcgV/JMdJxcbCxY/nYwU36cbxbgMv5bxwJleJxe3sNzum48
nwMTcMevWOuGCU79LpkaooYhe3Z7FyrBfwDihSJpjdy18zBMrrm0zyN8SAcGPvoK
pN+Ft5BtabugEqcwHZVW/4+G6t8c1IJICwmxSWBIvACvSZkboNwBLXjq25IK2PMT
7X/RkT16+588fZlErT49e/s6xAOU7tiot6jnz8gP85vJPjlvVvx2DN/MP+Wf2HmA
bnVZZCMAni0fBOyEgzd+0vUQiGZ9phztPNGLkcOK6U9+PlZJA/59IrADM8t1Uvl8
giss4szsYx5HlLI72flHj9AgzyNQry0HH/6+QnEbUiD6OINHSj/i7uLazV9MUk21
dHTeGRrXX3ZQXswN0eoFEQt2gbuy5tzC7MKPC2CI9PUJwQJIdxU3CAP3GFXQj8xN
Qxwpg0ttid6aVhuX9zzDHV2thqCyP/hS9knZJVKBtkMvlA0gMGKFhmdOJ67K8gLQ
8up2hfcwZ7HuCNkrjK92ONG0HMSDUwibKeaU53JUeqoe5jzSzbUoWSVm0RJZke6F
aeZcPSNA1EOpXI2VUj82bRcVyxAk9F8IEd48vFTDQhA0baBjf3t/TLXLKoSZL5zN
6A+uST/cabVZJ4Bud+Ch5NvLheWtvu4jQTErgC/MbDd7afWaYolnaj83AhZVe2Pp
SL7UNaoYf+HZ7PFx9CrXkHkbxn2H/3XJ7v+5a/HhbuydoTmGuwjvOdNfqwHiz1Sg
cMhgGmywfIOMWr3cgcNJjgOzQLwjC/UHt2ntgZ/lN1boqzgbl9s9gW6iPc/gA14H
RBeGqcbLj05NfU7jgmAvCQFuAYFmUmgxx4U2WdkmJuuG8hptMMv36XJckoY0erEa
J3Kl+pC3rAmhF19Q4yeuKu+WUfL7jRwHLFKfyNRcB4pYaGCR1Zz73+2hiLY4wCUJ
ERhf9uDb2NNtB3xU7FY0W1PYXEO315Ff+AsBdLy8DPLWX8vY8IPpptPqZ3Q2oRhD
1Vwe9cikNYohsm7AF/z44QCmccMEiUCsEYR7r3yiKabxo3OKDdKwej3gMPggp7Vf
5iiRo+28MAyv0oqWII5qOAeLph0JXMBtLMheyKdFIlDmhXrLKwGmffp7aLygYs7b
euPj3bE6bse2SBWtC8nsKS7dpnwT43SWTAA2qh809TKoXwnDXMBvjqrz7L+Lbzou
NJLNnYNnQhFjRfaO9aPpRF8BZu7k4WD4TKIKMHYSRx3FYe7BX0e7jSOzfP75zrED
gFT5zm6PIasuz59acO8ywjrlseSdf0mCsaoS15aPVjj8/vIC5/UK5GY3C0YBqc1w
t/oEnIP7gDQwJKUHSmKirkBo2KBukAQB7Twv0/0Qg1ry8SWrhwlysWtmAzDSyFYc
hdxifq0/+yVPMp96HJh1IN31mAwJYMVOBqnWJD892hxYigjVjWlKqrQHMMcXADcn
Ge0oC8oJTkUIBIfiMwTQvD33hn9a4jU9scmubqWCsjqBFUt6JQ7LerscWw0p4dTm
5Q0L91NEoBe9TD8aTCek8sgIFxGHZSQ0+BuwF4RIMDZHzeQXlduLKO9OuaCNzOcp
6KPsnXjnNxapV/UbiXTyjKWiriHNiFAk875mZHtsh1K4E+CWKEwGEPlJbwPQqnQn
dvWS6bn8IL/Vvb+2NqIRzeA5zzoUwkTczgsqvWdRq58ZuU6XSKrRwoJ84PIU5gML
2GOz8HGENGpr7TQ2YUvygv+R9hHsP8dqVqZYh8abk3KEiG97fDuaGPUvu2mQH/70
LQ/4KDuVp8bBJZ2oY5RYNmPMR53RgGCUaw5pbNLxbGJ5x5KkLA3k+pTkYwOotEL8
kCtr62JsDI4J1JX1Nw7r0wa6IPKWK8ndJOp7iM1R+53n9rXFCXWhqYAw/drFacyL
s3HI2vPl5DGNzZ7TAofEpf8m5ErlBQxGe+lTJ9K/uiCVN+/Qx9y9SrbRcgGL2nfx
0MhIs+0BdPzLgVrPl/TS9aqlyjEUCvb26WNkwUq25F+dCCR0ioE1lWfPGDFIEl5T
WSeAdHaT/Vie6ppAaeuOsdDN8o3An4F0NFKglIZFqrk=
`protect end_protected