`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
LlZn1WiQnJx96B0dQWSsqk7bDirGWRHiwBYBqRAG1O19z45VzKRHRebV9nn7axHl
cTf559fhVCLLbP7nTZzGST08WpPxccaBiHShehQPIFN6IWvzjcOPHyeXdZ1t1UJo
PPen5Wc4rx1J4xEiKBBPyvwmww/rdDa/5tTCXmEu5qOVmvLxTqsAiLm3NSKOJO7z
hqPRgy3V318XkZUX50C+YDDdjEbwWiRq3DS6RP2SedNwrDIH/krsSb9opJJZsRUa
eiC9dagehRgHdcTYbxIu1tcS/B/kRzD3igl2GTnHSM/qDbmoCUlzlaaUirjBIghD
6djb30guVuXmJHmpUu2iZiz46X1RVkBxDGY34z9ME2BP4wM9OGUviWUUIG5OQ6Ie
0KWCbe8WBwsXqH6qD5CiQ5c8TUAUoCQ+Rfyg8eq+02HxW5f8JoiRM4EASs4Z/Mld
LS2b7WOVz3xYx0oiQQ5yguEccyEZ1T11VL4T6rp03FGQq7pZpZj1OJwpS7MGaCKV
cGUYdwyltb53JAEOGM5cW6wvCp2NmAOB0hlhKe2ns9ZxVzKOOhYdKmmYizDT7Oa4
oGftUMG3T7mlrnUG0AJKj3ob70T4L+MCExyUOYgRMt1neu1+GI/fldbd485NacCq
PGh0Z3xiq42x/kdeWsJZUOmdhkthk4Z2s/dVE9JXHge22Zl8f5Stf61HFIjF7c4n
EaEBgrMJhbfSKMJupU6+I2q7Oa6PJ/3oT1d9agCAuI479k8jBNgqMooRemOoQNXh
A2HlfUeDMC+egizvgMDhWYrwPr01mglvBFs+ALYrxSSOxGraebBgz/UCaRM8lPck
gg3WsQ4NxiFYqULXzh1O9OQz6RwM7wscXPF7L+FsUHa5/EiSXdGtRVoOXn3EP8gV
r2ZneczahrlLcXH++HIyUIQKytnJjAkN3YA7F8FE1/SPImwKcKFET0samrboYcPl
X/N8sPxYhh9Wg3lf63lA0vWX/MAJMgrpWbkWRNMch8qsNhceUy3zeQW+IBkciIqN
9jKSNXRGic57j5jO+TtHt+GTZZbDqBVR6FxkDQXS7vWYGT3nmZd8ppmMyKosuro9
7EX90puGKjXShv4drnG7acivOIgBez91yW0LYJcLd54oy8wT/tos/1C3fAnyxR6r
Ne5SOXPiRL0/2Wkkmj+R2c99+hz3zQaPZOSs6qrbfsdugx7/9eRobx13OgGZg1Mn
Gjo5csL86MiN/BjUwh54ATqroBuOADEdqLlNT9cwMt0bl9C6EcpQDSLVUkZT8U3Y
Y4cy6VgF4nTzCpNEttYQuct8wuDpRe9t0wy+XuackSJvVVPIUPnTasQLMU9V+gJt
T6s/vGu6IyzRkM9X4wwONNBBO/+KNcCA3TJ2KabuD2ufzGYVD3/afN4SBIGUSG5g
YZgN+CwNmQdfY7G8tOQsnFHJuT6K4paEDVoxplMXIdwEnQ1q3hUzUEiXilsjgkWD
PicDmeSar/xiNmql6/OFQpBFBimhl5RoZdS8P4wmA5MmcJtx5B+JbISK7eaRovWK
mNC+6tXrRavZDbJduDE59/OqwiSC+29rYEsvVBNgo1oy9BMvdyEA0BmJlayJky4L
d7DmN6qd38sGd0Io7M2fP4w+6O3GZzqSjHLUoxFsq+4lVcBNha2WjKAlugRMwTnr
+PZP5LW+uAwBzl9Sk18hsGE/lzh3SfJWQOSgPqsljMEfJVO0Rk+eE+XJgXgkRg+P
J4PnNKRQJ3d5CBCwQbRrD4DhnXs1ZYEovC8WmSD7BK3AHqpH4hR5RsVHsVmxDeLV
OjhEz86QtLocZEqU9/c5aSRpBsCmOr5CX6d9+wAjUSBdq9SqXJz4yJX7ao0u7p0G
1ZrHMOySOem7ywBLi77koQh1ryfaBw6eVnroV/qmmwUrV6UIuH+7qSADA5PPdQqI
LgoGUYHz6+LHHd4iZgNTkst4WTalRxq+M04k3GrmTQRc+tYI5/d5QaD/c56O1Inv
i7bBVRNwTN2OJZyrQr91jYm9+AYWgaBPyqPHoeg0nbeOx/U3spsPG8MKeYe4GaLW
HhnSRs9mpDYqQFlFuX+PSrdxd7pWyvVAlbh7kRAN884zad5AcxKTgupU1zl2SgFn
ihAUrmwtVv9B/t6UMwp8g5txZHfV+UT138VzZlIf8aq1vTIf7Uh4A1rm7hiHc5RH
V6bYEo1dWm4Z7VjX/UEQHcHkPMASq3GpCdIn2j74X99QAIUDlKx2ZFqcRNLWvRJp
Eqe13lFVlQ/p7HQcidAp4kJ0/aB0hu/bZNK04LexVkecnZx/fMnnLlbdk82EssY0
F/3lmgyw1AVibYLHPgri84Q0DDvyTPH8NSoNXbevXdKLqkL7bAnl0gMJNW8jieOF
Cld/MfosvJ8f/0qJv7IRZhbFl2brol2ygZ1wMhm8WXS4ptJGL+Fwk17xrr/iullC
URFI0kgPAv97y4o62Md1i35paPp67DyOvzyhURLiDQIIhYzuye9HVXgFm63yBA6C
pBN9FolWWRor5iizG0Z0IBkES8prD6Ou2d7wJ7QNcPyyF51OkleWmIodFs4sqt1n
C0Xrvq7c9y2bmrtk+tVUrCg6KcwfuZdARRxAgM4ei2B/37Ab/XelXz/n/xed1ymU
kFiam3ESohs6OiMjjI0bZGCaSyp5iL1+mD0oKYJiPRDQ7QHaIiMPYEHN07oXOXuT
ZTHUzmJMNsyxETO6tftmvchq8o1zMptBBajyv2itkGTbyb24ucajRh8E+URpEtYv
rCQ/rtpGwzd5o3falJq1yHvLnNXgFeuhUdXp4CsPBecyuZQ3WW0ydkalcU6nIkYd
twg1Y1OwapG03cAAjBd1/9npyB1ndJdM2zK/7y9Fb+5bmCHV814QUbSEeeuUN3am
FU8spGGQbTNbiBN75m5e+r7BZtwBGfaoHK2ROjwdu+SpHEqaDUlsrGb9zHtDvd7N
c/zo/01PPmXch4z9+oYIRrwIn9xcebBZ+qRqb31/4sySPA1vh75xXhP1Y5gY0m1t
d0+50jlxj/gxddKciiWGx2EYP+yyd8xOb7oQLCVlvPSyn7dLNR/k4i+FlQDxmFTW
rYew1Js3Qc7gztA2IaxO2Ww8wsOKBG/cvgOQDWhKgcqZ0B+4Ds8LQUUweZTnQogt
A6Qj2YbOSjd72tabr69o1lE0Tb6vOxOm88ENHwnaH2Jqq5deuN0bpxPXfpkLdPr7
xDTLkKruhmch55B0BE7n8fVMJB6Q9mBezonWcmv03qpjZZFp+PUqcSq3AwH4eQty
jn7qcM84YT73tngR1ijXmbCxnSNBPEzblU+Nca/CdiU0IlBZlrNRszzHXKII9vQm
zPq/nCTIkGU9OBVm0vdMI73jHaAwG2MpOhPLimAayxvxTfCq6H4O2rQIptVzi61F
mRXSYuV9+aO5KseV2y07ss8zMY61lfsRwpSDt+NJg6NRrDZISKqGun8sdcXapjTd
WYWvhUHOS3G1qK5CC6yZTqlK9OY1bDgwnej9scwMUnaFg/t4hyKYrk5QP0JQVXb3
NZn2aK1YwsTZhd6hqvBwtqe6XS3nTgncHNYLFCT5HwfIsei1SCG1r4UE3BTc80LQ
JHQwzMLyLhArSzwqLch0IgwZ169kunQOCuqDYqcGEQv4t3TJrN8LYj8uZuf+PTqT
pTwTOYrY4p6sUC64gckUDCuV/P/DSFEsJ5v8liTflFDz38zOLexchuh9DiADjw7m
cpk65EfCdHH2kmCCZm/44g7XEVQNRx9PTwVRClkr6Y8+gfYxi6vyFE+SK+NG92fp
crZ8amadDeSAq2WMSwmrziN0O9ukNKxFOwXi49dOb5GcDpgj29QU73gW5oMEYdNn
QLyMrsa/3oOphcEMX4d+pdLl4aS3nVCyyb++60p7x1m3KSUT5L8zVJqaf2eDed8j
ir3FGJg59hYN38JMgS8KREWL+vHCIxq3KiM8NTMDGq4aAazPbL7O6bHdSiDp5JrH
TQZ8ZZ0ItsFZY46q9iFy73l6wosvxPrYE3jaOY3JASH9g27bhRvJNKg4CXtM/v9E
G4GPs7SHyFUBcDnV1EmIhD1dFCqqX59SstEJnwW34Z6fSzZndtu7bwNNmYngBm/o
Y65fU/p/e88cUP0QFshbXpi971Bjv+mFPhAmQBms9r07VIW+TCq1AhO/Y2iBD4mm
RTFWe3IVI2wNX/bCauYbsR1mW7keAvvbUfMdofHDfg9512m9VvRg+7B7T9S9uy02
wjAIo0d/C49HY3u5dxIwPfxA3ngpXJaqrQHdEwmwjIxZdjBwM/HFFrQTQA0MkcP8
kdrFmFkcNKzuI5XqkJQnCTp8bivXLJVpRF8qMZtcEQagBx4mn1Vf/2pvks7HIs20
OiCKYMBb/in/+GFP1BAeRKZ8FMXgBjkVL9YYGVrobcFFJA+fjHg7JGt7WoKoh2no
s9JDRrPjoZWPLgoBOP0z1Nn3BUzUJlrqjpTZazLKDKXqyLd+dQeqJZkrn+wy1QLd
6Z79GPXGTchCBtFZLcJOQok5S9cj3GvPPScbnuIlDH4OSosvNY2/BKTDSlr4+1XA
zENBiORJPDu+ZVA0OOhns4HDJj88lD8LsBSIrexaLDyfMxi40SGx52erVOomsxlm
p/pqR+GTkUn7bVI37ys9QLEsZF12okssFs+ALAIOj1KevxjI+ifh6raBXwN6twGZ
J8/ZLRexfzGQhtMFiJ30hGV9KqFXnBPtpcNDZLIocjEemr1qwyiKKhvtlPQ5ID/5
UpvoYRvUbtcfUnnX8YbQ6bxOWgIQLtV13uAN8gaCkAmi2F07bBvs+MJQf7jI/U6E
er23j7snjxM5+pAvC+11HXLoBNiyNeekx9qya9ZAoc68XjewTSPThgIoo51MANzo
EouRbRKVbgzD7MX/9CP+l9rDkB1I3ApS8f0wyoe9Aq+hhL95NYwAKKLgB8Fh4axO
lNIyHeLU63UAoxt3xqDpoffMAPnANxKnzMojE8LgNhP4J+i60m1u1eOhHARi17Se
6OLuO4IpXtC5LZsW/SMgK1oRT3BnygXhlXAFM2TO44vFrXWP0udOjXjYTch9rhYw
V5vRYeZSJHL2Tx2tEDD9LszRDwo69iBQWXPUhM0kB9QzaER12KP6M9XL/EZ2eGD/
B7ssBcUBt3GaLIB/OX5znhsPjM+7I0DBqiBy6J2ILmuap7xXpFf0nzY9Gp+kXxO8
3mWxiY0CqDW/T2aXjh7RgV5S0PAzPoFqdT6QmpZ7lfIQRXPiLWy8zK5JE8AuilhF
H5CTMSqFOZV59aprxt0xewMG95ohGKJhQlBoKedX3qbKTne74n6wwgJSJLgG9kzl
QPfNck86tKdtaedRX10FdPtC3l1jw2Y8P67YvU3WYL4c57/jTTqNTGYiYKKqiDE3
sTf4BnGPXEkvtonlqUgnECPu+UFMeuV95SoKZbv12UnVvdkbWqQX8BqyHWJ6E1xg
7cmumgRtO9B1XG7+FXjuq3OHayg8ZHmV+DKsRSqAX6YvmOH6p2K7BAJ87cBGjaeL
AosjpwKasoOyZIeIOJwMxk290ntabIHziSFB2J7kg0iSWudl5guYkSeMN6zqzck1
6bUzrscMKebp/TCS+P2GpN4iEbgzgQ7rdtw76qIUVQ7/jHcgF3GQtY4+MAfjCIxN
F1fdNqGZMo8XbEdg/baDdWlUf6a4VuK7KMZ8kYpcaQiU3tqithXdwwEfhgUzx0p8
amUTMyJvD0A3TROnkbD/z2TNIHoUzMk9VQvGM6/ryftuzF9jjBbe8NlWVd4I4LsS
zzTbfViYtkYnWIeUWN1eQR3cxUMFc627X23vqOISfrNOay+9PaJM098dl+EFTJmk
wmA9a69Mjcy+z23Bjo9k2sze4Cx9aGZf5YLLiV9W2UPBE5B4FTbISfhJuaO37Btz
f8NPZr4JupDKQYPBBvqozF/j9ijg9wFnVJR73wqtn4EYtFabAoi+UItrmF6Q8Ic0
wUdPHgp7BtcpKdZhArlwUlbDM3qUPNqdLP90xaQTj/A18s50nVYFzQTJ2u6T5gWa
ZaSJZGxDZ8ZeIjgGY9HQcWv6r9Ovc3ozkbWKweRp1AXfjxelvscPpK5e9FgbFXpF
Pl9KwXJSOvmkBqU3umAHCGTmx+9Q7XUICKTirOSPguckHIMGeouyfjF4VA6tUY+9
DX8LmF/KlNAdR6aWQsra9/EpeUgfHqKx0SXqNhqUELub7qfSZhOwp7Hm2L3IuADF
GpJ2jjb1gORqRcZ8ibJ5FwI8kgoK5nAUjWeElW9+6VHZeot5JHCByXYZQdusNpgU
wqTjCOB4Tmg5UjNFyNEEJr36yt/NSx/BGVnGzk5sMo/eD8V6/fNu6mkSVazOCMSN
eseP/gRBPbkLYZB3mYp5TNX394i3KmUE1y/YIsJzoKdZzJhBogJj8zisWCi3kTBj
ISREY9Q1g6Ojc+s84CTbNwA+98ObBz8of1DaFwlpQWBFyhhh0KXdUQPHzTl0PlXj
THvXccGl3HOVk8izIzywX9Iz7W5ec9aCGI8IFEyXQh/SNSG0lqO/180o45u+jrKn
w2DZWz9obJLCvz86j9B7kq6L0tbkb6FsPfjLPlCLP478WQdIjeC46UktmE20ybhW
oRdcvVvQ338NkI1wc4ZO+v211X6/1h1to03j4anSBv5t11AbwE/rQb9elWvzmalS
PpGwbpfDXbX0kFVqANA0zc08ige37E4Xc9cI3KeGdCzLY8i0C872YAN7EXSDjiyt
SIhRdxoLnNTMLmLSXIYv6kf+nssuRw/BjvbiqyECu3FzVO30v5Rzcr5NUy+tpQG/
ZpQszxtzViG2CxTM2c2LscDJSj8GO1EqVMxbTVcEfyOKSnTLx0qw2cDrMOa19GMC
NOU2YOyPoL8S8nJ0upgXE54u05pC6FBPcEs9UN+ldo4YpGgxdXCJxEVqFegHsoB0
lP2LH9lzljc9fHDH0kMJQI5fr3GN7Q4PN8quqpjikN7nGa2WyDjh/usapzh+JJRw
7SZAvrv2+WWYCf/QsT2oPQLQe0Wh3xa2DNLvgPseZ5WEIZsB7iQEaKnMsvHtXFaV
8oX8XW7DAWYcYHcyo9ZwApLv6zcyA6+kF3gpCasHARWVQDAW7QALlKpKl/ZJE0Ac
J7ilwNIF9RkBCM4REL4y7JF0Xe00SzUv3pY3KUfM/NUln8NJlfZg+obmwkfxlfxt
Y6H0bBKiCUHiFq+HveKmZwvTU/hVnQzPTIfKhXEX4U8NtfRLzJ5AP0MEuF3iCY33
NIWSgcMlgBY7Q78Gc1lTC+8YrxgfMVLZnf8LGfT7NFWJ+PhmEbECj+Rxv7ES5HEM
C8slx63YrOLmEL6eTwIzJhgMV6RKs78RDaAqakWsIL56MYO3QOcm4V76YL56tesq
5KLtZoCbAP2bAEafX0EIaMUnEKuxPbl/jgwYLoA+Jbjh5R+bqRiY30CWsiVhBsKk
p/8gsKWfFNjJNRNQ8+vF73XosizvMPoZeZH9v152wTJo+cYQ6DMBMHLlTAT/Qmuo
jDfrOXktxd2m3aZfsg0fdMIz1npDBO9JD0RbMyfWOy1U9Rgh1PVJtrvjQ+AP1bA3
0W6yb1NHbvXnE6FRrkcjjQUyjkTfXd4toeCCRiiUAIJXSMsLJdhoNi94XKEqCDLI
jtODqKmGRbYus3w2iUsSh/9z7JzMON/BwuWaimBzrpByinzzWexzk3gH2w5FbA/K
taL4qJmT8L9Q7dHbcPZNjv89W+3EJ6uRbQED2cm+lWxA8V16RgV+35xCinbX7us4
ZKPzrvXJl1sKI4NIYS7RDNJOMZ4nVFWii4BukVAGvRMrOKqdhxT0kx6e1TFuivEb
acRJTKZAaj7jv5ZhkULZEsOCCCegMAYj2dolwrB7dlmhFBgIJAHfFmCiUbwf5J7M
qh1u5tHizq33cBNrsi4CYH+VVTNSoCASLwH3XuewLuVwySOkqsMhElBFU9P4vuU/
OzIVCpoJF2qT1hQHNTYojNVGq1H7y5F7kp741cuTVTOWbAbQRZ8dQHWla9/OAijF
LOedpVWnQjL3nRuvFcZzakmyUGPHwyF0Uzi+qXmyYK6E+vEaM1YqsP86/ts0L2eV
/XO4hBexB14e7jUju9moxRn/dJY8DjdOWJZcOO7vwUn6FmWe4ajmxG+0QJn4KVoC
araDspHiOjXlYfCPUPbLOU1CyNlfikLsJzIyyiGXuLUEWg5Mzc2CXrwuuqULDMsN
Z/H6pevRFpU9qYvbORbArhlr/lVEtoRKgj1jzf1e7nuFHPH4DJUaypn6LqMAJPBr
EmZlt/FOO6lwxmLfRwC3rKw3ekl5GZS+XH4yNiDSRzWoyl2oh0+UTIw5Ld1WDapu
78qbAusVTLFHuCW2ulrC/6jlfS25+esOddI1FS5lfApVuVHbEuDfYXj8BNHuNZP2
9zzmtWBl1OObwXGn7zS8073Z5cxQiz4X7AJ2aqS+datfSwPxJQatGkkzjvQpxSMj
a7fAvjCqXTIwrDBYPA7Dd0da2ST7TKK/DtsyMdcvbjzhhK097JbsMbOrcvjhZ0i4
lyo0cPnvtgwV5El0NoQ1yVYLRrLMPzy2BfLHZUDVfiEz0dx7TTVqjcL/CAN7zNZT
wRKajFWxPSrU3Yxu+FTo9VWjUiurOb+Y5iVMh7jeVXTHjaHTUhJN/muzROD+wH88
L3SW66FoQPWtfO6WrJrzBIyYkKHHmUOqQvloALoBJ59yrRcMf1cHiWq4wZPoUYxm
or7ASgQflrSk3QlGqiq3AnB6uCqkrr1zP8d6zrKTIuQ=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
AOm0ifrO2lG9CKGJhmiQI5JMR2BN9dR/qzaXxEtOcW2Z2DkzVJpvb5vn1EMxUXbR
d31iqXPkNALB2vhKJahkWE0Mn+r+iGhWo8YO8HoIKDpJvZXhtdAK9dPvj4Vz0gu2
JTnCRDlmNErgz5TDVqTj8umzdHh4Dh+I20Nzi+9LUo2XEqwGaxRxwk6ie99xjrKu
bxhkaBSzN4wMPrmJb5pfc4HWj2t2HBYCTPFRnvpqo9u6m3TZ9tLNqQ+2I9inpk4F
fBbhhf4mnNPL9AAW/Pfs32fgpznyVC069YupgusUXwmse6LEN/nVFOa7hmVz1UP0
zuIR7DmrBSzINqlUJtJDTnQl28Mdy0KdA+aL8afwJIhOUqEsKhnRMfo1d180SDfw
WYj20K2vrcgp+nWaevf/dc7ASwzAI+Z6Q2QcXfc5cyvpGpRAjjthjNoDkn+Z2Ldu
oFq0WwRMpXQryX9y1xw2kZzVjwhrkWvJSDp+8XR0bGgRhvxm86ecwXGpR18hPx2J
T1JHTCVLbDOns+/MFiLtwvLzdKWko667aDswaoLLYEOeAGxcyfZifPtFNbBxJf3P
2Otf+re1HfK4qYn6ZN8JhxnHZjTMc0Y+KXTicgwDkZ+zA9DmcMVWI74/U/H9n4JG
M9ELGgt7B0LUB49nfpP4tLkSZvJg7Nl7VmPKDSXBAD2grplPhwt3Sz5uCfYUw5b+
Ekdwpjed2U7rLjAH5QxxurzBXeCSv/Z/L2yGEggpIJHTNGqn2i6vPt+/0OtJck8R
UYz+5kNn7jJlh9JdENeMAcD2wzMGHJW8EDPOh+2+u50Zf/cD1gVNOq0MazoOrFDn
SKbEWUh+YPf6jc/v5hBF2oQwfJ1m1c1stPo/0+Q91IJ5UorTjJlvotWpcsysSYTl
xAfIQilTWv3NOosrXRje4hN9QSehEOa91+qwvRJRNJd/yTe8MY94QR8RnPCyPs/n
1++JWlXStxTO56nOibPZoMD++JpGZhUX2Z+JMRkyr+zcWbuPegEs4S8Ig4/tQRcF
LzW73zfBRpfvwzoTie/zCngYExZY9BvGTQPFk1cNZuAsyn2MOB3UShnqSwjT3Jnr
+moox+a0RB9gXgWygq5433SwRj3Bze6uaFTCArgSKVflxBvYazAadm2WA0115aCB
3vbX43wss9Feo15hODbcDZXhELO1CjqaC4wm758/z3PzmwNUG/7CTcpP4Hu95px/
75TXFWbY94vLK4sPB5QgQ/QnyhSm4bYFLomcXrSIMftVB32QLNH9f4toUBh29T3Y
gTMvYiMBKTHJuqqn8nG2rwiqwjhcB8Kw17IVctNFAFMexs/fiEw/s+y/Eli+os2E
fZY3pYyXycsOhlttOD4mNiZ/UI7dithfCT0aj14DvI3vhLsMUs1yk2LZIhAEkFcd
sskhNh0ogZEA50xLbaI1rYaUy+vctWwjRDD+JJ22+d2cz3fjbs5Np8PwF/vh8S5S
3ygucDb9FLIBdUbDNn8WYt6kFLHrJIMocrx34QBhXrmVL5FVM1nHilYExanDtLtq
ZP75qLt8oJUOI/insD2kyW4rkOP43qzgiX4zFkR7mUKa/jRWzqE7D8yYBhT2Xzzo
1cxAIk2cnphycfD9NREL160zO2HLRdiei9KpPCChS7tnXu6gQZInfIoCa01Q+US2
dslOTAFMnfNhSPLkfLx+ER7ATFL25XVHvxWmeXFJ8Bmm9EPXMrScaDv8v2bf5zni
8dW78dIngk3sisrptnSmNnE6r6AuDJKZQsIUS9lZUiZ/YgVIyv5oWe6G1Ku/dkz8
WwtXQ7+VZlccJ6SAvJBOgvi0tr8KqWxKnunLWWHABXqoc3MU5YnKMr7MwWXEo0Js
NxinHzvlhfWME/wLQucUqCm3wL2iHLtnNfX+Ly7d5j1rajHJc3IBDrXdfDRrxHtO
w9wSrOqiDVC4gXcCFioSbzG2v8u4fifaOX/9bue3SSWfHABR0Upqtahx6bgb1IU6
lnliHeW+K+T0LlNfqSuy6DqlL78k6zT2g1rHotHEmgEx3v8I+y6waYs4TA6Rt8Lm
0+PpLIm5eybAwiJXLFEK2AorVVGXcJwhL5I6+qP699vOeaFOdom0ybs6KZONqgKA
YKqlAw6ifS16K4MqBIPdgv1dUWdfEcmWKZE3f45WLI1SLnv33InhYd0l7xIDl7nG
TBlDw5YZ1nGGYQhEQ5tGTivt0ulfM32tkEbbRHdtMdBAbuGP/AHG1VQTwo1Ld9S3
nqPfqbp6dcGqq9E4mejJczIN9PPmAXUAiLycH0Nc5iYPOviTxaTn0yNwapbsTk9g
cN46xegh8CBkf+i+AGkLskJ/jcftxtK1DHOog2wOnqe8TrdPEVDy/A79VAqbdxEX
f8VO9BL1ktTlv0mRkONeqg45bTL7HLZbJ2vDMjQ7pOWfhEZzOWallvggeC272k1I
Mvku6qS7ikDmY6OuRBHNHFBMpRcghVGM/ZWJl8iE1PHixCNXbrWzWF1NS5tWec9o
M5F9ly6X60qi7DoXluc+wcv1ait8SEXaTjZsbfYip8TjdFP/h0+gx+tbYHG18lUw
dHUc+TANIjt1LeeqQE5pTczPLIJCIgpMjJgCSADngrkyidrL6wJS2LNRsfSkofG6
OAioB1Hzdy4S//7GDovIqvB4M4/PCJ8907f0We84cPVq0ePIkk8hvwi0Ab2Oc3SV
KP5A5rA9/0BIyF7/DircppYApq0Xj65D+4VCvY7oWdbHWOxCq+kyfjn/6UuSiMVq
ds9U9KhYPyfHnnt6eaKsscloPWV4fT5koGHNBotFnHbjmqFTtUbk2Yk/mca75GNC
6F4DpCNxBTifBzTH4MF4XcCmPFD695/LjthM4850mhZoYnNzJ13J9hCJwUJp/TtP
kzfoo5V+uOPFgUJ+58Z361fscTmpuJ6f0ElUs+lDmAeZ0Alhe/pRqTMNuZdfrW+N
MCIgZ9sWEchaoxj0Ipe3vWI0GPFs9zlIi5+QDu+HIECoVGJBO0NGQKtabWQH/OUa
0UTa6qp0lQ2wOA2wESFEyPkrIAo6EFv7YehdjzA27nugnlxZus0vNHtYhFgfpnGi
MlUOvySfF+mJgso4311j/8MEB5B0lii6/VR+LS4lsExbd56HQ9wJKnd2ArU1geMC
R3u49Pn8VG0+hImkLAfhRZ/If7SqTawmEz/UNdSrCaX9PJje0e9/C1KuELo9MSAI
Zeec2fmsUofG79t5DcolB8PIVAd4JawzpfxK8kAofeOjrIdq7UamCfmtHxjbN0eT
frSp1yTLPPN/yU1axWMrknZsT4ls9+T6cibit+j4OFvQn9RSi2hMp+4SW5h6vjMK
hsTjOlAbZ2ZPr+mjlp3FcZmBC288RunTQfQ3Ucf55EpjioqNk3yFzqwlu5/mQ7QL
de01hVa3nUlVBGvfAqQ2Y33JC8VOXw+0wpJQSPDqFYjfV7OH8knFeuljF3/m15O9
C5GzTB1qxqc5Ry4E448QmWnbhuuV4XAuEP4zy0L/jkzlfuC17IlO28OAUP8570Dv
PEhHR0TeVT1CuxhT9lCTtbfdYjaiSla8T+FBHCZd961IM0yACs/X29XfOYPKqlfe
mNH6ssChayDbQ1mp57gTNSLUTEC/y+F/CFS53R9WIp61lIpaRQJlnj7dxeQuwRq5
v10dewDpwZK0EkO30X8cKxWFkyMyZSBvZFPbQu7AjcwTMo+Lfr0cdL3qlpDMR5WO
kguTbJvNqB8J0DBcFWCs01MoN3IFn8bSp01Q1N+mA+nh+ggDw8ks3YuSE+ByYLqk
yZN6OoIanvCFUQwBmEnElx/5C2bQqWnLf/QmytQLVGsc+oU3Gtoc35KwCgb0yW4f
nHtLvU2Zbt+2EH3S/1F4JmQllyOJ9uxprRiZfUUne8TluSSvPnCVjoFKP0dqRNY0
8wwkxVkmFkVGxicNMjjcFaAFb/JMPlu3hrIfKCi3e/ZDenVA5nIZwFoCu85qRFhz
R+SU+4sSd7MeTiuqm2n+kNWwKWIkCXRBf3KJPWs9CgI4W784VjHvFjUNxnbGYrKR
WMltv9Bq/srbNEfM0k1HsmzslCYj4o71r53iV64t8GGb2EPY1L/AI0Gc9di5yqxX
vwYL/UysQw0lupcjQljt3RYPMHXQ9/N6uns8Gme1zAFiDaGYxtS9GTgObRQlCkzK
zYkLVYeij9d17PyMLcIdqQMUnTymOHJEBQfqP6PzTg+56dxK0RBOUIC8d3uOFUBs
o35DM1kcG6YTrjRYPNx4/h5tgKqQnqFgX32awA/eUIR9BAesKvYUB1xBkrtItSja
+9OvUC9cLH+OlLuaqyrhtwf/Rg32Em35Ioi87tN2wYSS9iP6+0jBqFUe7fUIuK6O
wWGnOVp23JSxbBcB2f5gSLm9U73wCc7sNZleP7IkoZT6US/8F/OcJh9UZY0Tal/i
gh+SyOVSbeM5Ck/pFoYI6uupcvrHl4gPr8cmJW8Or7mfO+coqbm5wbMszsQtwi1s
+6sz3OQWhL3so/r2VTzCfUZqWRFr6lqX7oj1X3nhLV74gsSyymYTRjS11VktR3Yk
Qa1+bfcC6SPE2Ps4BoKkxSY5gpCQvir5d4Lznl6Bsg+edqAJNV8IOaPIRh1yR5jX
HN/tte4XadbabvydFD1NilyCojKu1zV4xmul6OEYIgUaO2YyNJr9k8UTudIGEMBC
R5P+YMByT3NjAAsjd5M3fSFZtcqnPBFJE2+6X+gk5VfQVYz/rhD6mYkgVQSqXifJ
yEhvxozhBs8TIFBuE2fesuHSYs4XkwHhB14jPOpdvNGo9181HiSdOMedxlbcmSRx
HXkKW+QmVjntqjOdTwQvLKykIvGKdhgxcV/BAZB+tkH98usERiaEaak5MRyL/RYM
BNOkMNin1oWh697O+Hqh2X8oUAxpnSSqqQRMQPny2110E0Q3wUrYSCpKFXUbFLKG
jRRsQ94CSC07LFQ+v31i9xTCwPiOY57egesIe4SusC09c9c66fyOQDKiZLduYrag
9HkJH6o1BbI0zsQ0YZqpdPKdpVWsE4/X+sBGOfhubdxzNveI4ZbyYdSmUl2esbg5
S39d3+HXsP7CVrQI4PxthPtZMFjpH4ZnyegUfyRWypfioIvd15Ckzt4uoQj9OqC1
W1bWxudbz5MMW7wH8VBtiCaLD5UdbXbLIkVOE2rOkEZkajtYkd6cMd3yDT5WHTeO
hSfvN27GHSm5jLhaUpYaDEnwC8f+KpE58L0xf/rGjiPgfEt3fL6dFiwlY44BZG8a
svpkZYnterjoJwrAoxKJ9vTHzPJoaHAQnDIJ5rH0C76RzsicUnY60wKH8X1Xn742
ZcoMta2tV4oVacX8hRct2vQgGwd1YsBiPNLJd3FO19edVmRuLuosnHLr1HI6hZrr
ONykT3C7C59Ou18aaIlGkDdh9SxU2iy8WvXP9rXt7mBSH8ZzDTAnBuJwcm0msauj
9QPe5R2ApE+j0P1nfj9HV0TMVqtZjXNg+lLrbqkekHLTdgfALCT6lSUJlyb8GhjW
nbiVzlD7PSN4z3uefksWoR/QAiuhUGPexejnSc/jlWZs2P9Fv8HCHeLIhWZUOx/l
mx4CoVQXuUSepbJorwFW2k5NeBzmex3ITlBJVUJeEX5Pigu2jo4hk3KPhQslCqcd
tn1OzJPMK8j8fIjTbdQ/lxoztbK1V+tpw2C54fUrRH6hX86dboWxwJ4aRwr92TPP
llPlXwmVod1TmnrbYrV/ckdf7ScPUqPhsk+bxfEZFBY1V7Y3I7qFluOrwkfRXdAl
6pBGol2fsaY188Vfa6uXjznLFHatwBvPuscmn2yAmB0iGUM05EaGUeM4jnxWbs2l
mfVLiCcBdOJ9g3+XLRrLTRnns3rHT9E776GMRKA4gLKpdS7G/FPXfMhcVD0agOuM
dXDx9zKUX4ljpr2ChPqvLBP690LNeikwmt+EoK8A2tWoPMZpz9+qIZxdKJ5CtNDc
EAxzUbHhH/Gs8BPY7TMhewmVqZ3zEmAovZZb1grKPm+ILW8RwIAiF3adiLlDHpud
0a+kMkJEEHrH4fQ40CMrkMC8Hmc6FpvL/3pt/44wLzmuKXyuOCBhSpL4YDY0Blmx
LWi7KqxQTABC06/+Zejn+wk2xDM5rvvQIxkygJvEiPaxbbAYvpFxXkJVMPMqTSTD
y4GXKCUyCLXGLwVE5L4O6o2D2quvwe/N70Fo5qeL8QzGiv+4xqo+PizkgIxYyt8d
LucEYIZ2haeOjCSFTsZBpA4gmnRDwWZRkbz7dISS6iiNQylYwLGz6kZCpiCRQuto
wBoOcY7XeNbSexcB/Zcxoi3Xxknnujr8qvQPvBtxJRPevdnQCl9br9ARWn+sCF8D
fVYO2l956tT1bDpcGjPJ51wyxcFL7z8MfHyimeMLkEPWCFPPUq5auaSqeppJ5hO1
DEGm7XsiAIaEx8N91iWcvYMMyJxND1NK9r+4NObQSC0EmqgIlpyYSbhu17kEU1JH
2FuO57xpmk1ixvBMzX92hmWxk8b23rymxAdScie2gTy0Nb5oRFII/+NnCnP+uZJ0
dZE5hvnfhpEUQhWmnKcWqlVBE/qs9AZz1WiBVimgg7goA0ZgaAYMBp9ITrnhN985
c0L4Ee/5HYkCg7DRMIkm+RtaiDoH8hO56WdoVgJ2YbHHM8ZggsLDWo2XJrBHR019
tbxAQIMGXocs+VTr8VYxzZCmCtuBtyph/iqgFg4pXBJBeK5bbAD4gDoMz7J8ydfN
au39gqS/gETHZmuuXkshZNYhjFjYHXAGCLJUt0lm6OTOtcWATgzDRCHuVgqPGj6Z
Xn1PqNVwaN3dtvSom9FN1UcPEBnE/VvPTpLGiE4LmY0riKJJVIkntqz6y+vmSK9z
Lt4cxb/9nLyK86/wexo0mkCD3LFFD3dQRwKrgNjuLi4I48+XWy0+w22h4Qapi3Gq
mGajvGz+X1JwwCjZqBX0oRDD5V7zLUA1clDCDWBuAk/ohPON3wt07b8Md9K1BZl3
srZVWJuSzbPT1sr1CxxHMw3MXf3GaLz7UbE5qlzvp81FZisy6+wClm6Z/3G9GSui
kS5cb1AY04SEqoUvKUX8dVNEZe9srjjbTagWfzC+6bBTqd8wntpfNNgwQ6XhsJw4
QbBakT5IiwHcCcEoRUCcfy/rWKw0C1ehbd/fK7v693/qYdJVYi5JXuXJbo0Ck4GS
8VHMJtFBw+G9wWqhRmDqu1pwm1ot5o1e1v4TvqCySnHhCNPcjNxj96EXVq6vtwKa
lD5qqQP2BImtwte6Q9kRoya+XqPLoIpGqMXNScOWY3NyeVlkggf0tKwnjD6fHx54
rL8CE8p3rS4pRl0Jc3tOJQz6VvAYpUEijNOMremFEX9OLOET2gR3VLqP8Lj+cmNw
4hmJV/ZE2J+zHI43qLIEpztWdcmKKBLojxTPHZmkJWfHVR1Q3eVGV4azas/tG9+H
Z87MgTSVxirFLLtZ3KgOyPUwAP/Z5kY0UocTTpqpUbdbSP3viAV1Ca2cV85Yl5X0
szqqY0P63ZHLfNsE5XkqFdUbr1PCoW3xasNuz1ONXaIy+Y6Wj7//NXlVZ6HcLyyl
GJP+NlNIIbLsmRx3FkTK8wf9SzJm2t3ZEPqSYPHru3hgido9vR5DD5WHYygaBiOt
NhlTiz1098IGGXBYhkafqtGBWIvCcB+nwYLmJKAMjkIZ9IqxSAjqYLAC44fevSSE
VWTaiYmrmQb/2RN8CgfocxgTWCIY+LY3fyziz4nm7C44rSJqSyVllNN74jzTP5zg
VvkFwJIPcYLRxYw9ilhHHUWqVXeVZMbca09o4PPYJzDfocurla4YF72lnqC1cIuA
3YcOzhOyg3g8lliIqamnVqvebXJrkc8S81rBaryxylhZsbJ3DtzipT9y7SQEK/Yf
CMJAvqXehwFtper8nyn8KaYnQFQp0aUI2C727W0RDUue+nkwbvVYkv4fb9zGx7iR
/BDesKJ6QigDKQIUHaB5ophy3grCRgCGz+AakieMHvOAb3qX+5/O5eiInN89HPxy
g7aoodm5jtj3+i1NADslVlPJ4jI6j0fMunI4iFy3DpMH+pR9Cnl3nboFp9EAGHcp
2NiFrlkP02irDusMYdTQX/GY7EbP6mJce7nl96vv9xzRkjovUiDaCUr4S6wNarUR
bTWU8xh5mPfjq1L13FBZFIfILE5v8w+nMtpjD6Nb+YJ6TCiKgKBQjF6QvlyeMHi/
rT9LpBtn7jVYYGM4RDfRKjDyhsEy2ifAKMPrvGc0ahIt/2TeD6TRi5xvRVOMuAVy
eLIBsPgrv/R4zpqBYkfbr7D3QBYVgzt23TvYjl92w4hFk3Ow8mJKc6OXyCSqLGu9
VhZ7jcI3fIoZoI3RQnWpFh6LyK+sL6IJSjX8LD4pPrNhUlxbTo8ndkxnldTg1Na/
MnBL3aGXGhQXevEoOpVbFTmn+Xn8AgawU5fwUER5Lpkf5Dve0XDn1zdIBW1PBLpP
plQ9nza01baRn9ZtueQtyosXqMaHiYqwbNS+KLPZ3JhRVCP45UiDnUdnslh4b8c7
onOOM4IodIWPA7RPD5SULwo8C+oEWP62koMr/vn0qYxjZnMRKJGJdt8/S5tx4b4z
Oe6JRn+mTmJV+w9vwV4dQC2vFs1QDs9SQ1ZAxn0W6yD2etoJ5OrMeM2a6fLRtglp
crVP5zM61ve3Vdowcf0wcvwK973euzX6EMuBGAOKZxndRsNl2WXI/YHmlYkxgdI3
I9wFTamvMDu0GMgrjZ9yhInvsyr5acSaKd79801l5Ng=
>>>>>>> main
`protect end_protected