`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNU0BxIRMWGk/3Ou/A+L5XnAIw0fkhfJoKy6XrHqPZWyt
sUBU1CTUSq0dqj79DtY718tkPLmBBMfF5fUdXr4sxG0GCbwCFzF4DOO9ELvdqwTg
twshJGdutAmr7Pa8tLVPXOKtw4koSnwKxeKfkiTi1ZStCyvs68WWROAiZRoltiAR
nfaMiUEmHz+GCY72hh4B+RntORww4kEDsg17yBGyBRIBr3bQ+NCFx/73QvfZ9X4e
kLBf8j9Xeastsuc5VoKJx0ceWsBWQnHoBJYQLjzS7bVYXnFSKVlGxvX8tVVGcVwt
eW49l86tjQG5CtZUwHTLkdtVsUAp5NKJFWyqWS+1AQWw9KOvG/QZuUQtBds2EKD8
rBTLWZyuGki9Yermqq8RTNiyYApopIhG8UTpSfA53GthvEpHlQUs9fCJc6jy5jqQ
BlAluIXlH2dsXeGhm3+7iEhHvaQetuedNJ7hJkxxdkbnaHH+0wRXMn/rZJCkS+Jb
ZAE/E0uYtO5xDzjpQ3Wuhzf2cH5U9iKy5cjvEmh65Uj3h031N1hbPxH6pEDl3bqJ
xf5ZaEoeXvcsP+6qafA9JvwoumtzhHzugzQilNDfdJ+HNfKOvVTuj2WHVF9JKnF4
Sf/9lPmGRcRlc3IBdeJgxRFoMsMgwbjUq0MXJbwCdNq6QdYeYW4R694Q1NUa8afK
8t5vKOXpwwDFf0ZuyipzHYB6TKk5NjDVtLmquIipv/QiJLtpBa0FbKU+XyIIgy/S
JH1xqg8PPaYzvkQRVKFXlU5mlNlkNRU7zjsJb55YcClu2aDhnO6j0pdYAW0NLyMe
+7eCIDWJxfQfWtdi4kBxUK+4Rsspxwm5KiKYCHGTrRtjyjwc9ejj/rIIZZlfIh5I
mfkUK3kEbN1iVmu8aBhIUsaQdYgmI4IklLpzLgapmFr6MbzLrCriej1DcvjQvXoC
62nZ074XR0ZBUIfwtMLjvydqkukZgMlKBL0GAJg2tH34F/8Mx6v3ApL+P8Ri+zhw
brCMEUXE7qPzQ0Ss2NWF/wpGZZYjU/XOQVCno7azNuHyEBwQRNXsegNTvyuQDFJm
G6WMFaKT09BjTC68r9/xY6YFWFWdK6C9f+QaL3m1/nljdudzYyGdenRDjGqJ9bcC
6qycLp6XegkeIH19184hqGRjnKXCLDqby6cGepztK0OMBccChCwq3Z2hIDSre7ft
fqyrKAlZ+v4dj2h8Q2tYWBRnm/YidopsXXpq9hcAhN8Dfrr6/dDKLeSs4u6231gv
Jq2VM/c/hcnQPbtB6Es86dqE9Bil7j93EIOwc3EPp1TnrX9PM4zBMzIejYvXG4Ja
/62FK3W56GgCM2AbUIKmaiPCtW6S+NhH1uwRqNCt5eGGAov7DuP6YvaYaQpdzmxD
ZOL2qchTavB5D3soWeyBiU25j6iUcl9on2jmN/NIi/yXzoKJio5sX6lVQlj08HdM
McdK1dBo61Myc1C/Ime2k+biEbbVJk95hTODyyBpD4ubG5tNSU1RkzNXn83WvMoQ
+eLXFjcoXuH3Ib8l829VhYvdDw8IgF+d3cAcnBaD/IMxOTBGQ+hwuWnRBjn7M4eT
GKB9NaYKvQnl8UP3MBkR3K5KGu9xfh0hCnWphntJwsINBzIDhDZFDTI9nxQjeEYE
GcIslaKNEFR/FP+azJ8zRn5s3EjWe3yc11DQLlMBttRNPqHPkh9iZIMoxdxWOL6e
1qGcDAsQRfcH9vfctePdeyMmOwvOGBdR/uoqQl+WrL8QpOzBqsuK+aEDqG6Vum2f
5yfR3xkqYisEsldYg3VJUw/HGR7ZVyYmpK7ZcVglAtz/diX4c/QQYSLm+Tg76D6/
1FA+NXmowIUYvNSeMM/hXwhIm1LI9PwuKgqp4Ezw9wkVZYFMmFmN5Vxo+7dO1Bng
SNRtgXHTWp0XiR8xK36nRzTXSAnCSV8xVbRlLT0FhF3X7laPcLqh8xpjXGB2Osi+
kqRyv69IFuHqAGUqpiLcjTFPfUn51xw4yErbH2ChxGhtWZuPG+1AycOP88RIDvly
34DH3W1VnwPGN3SyZJ3r9Kkcg1E+FVKlXyO6kxcsAnnb+JA4jVZwC+Y2rYCS/pRM
Rt5X2VIC9+dJNzRc9DKgNg1seBZWVvuqqgKmpL4z/r8PXtg8ojb9JgM0CXAn3mTs
xJKBAnl4x7cbkKGCJTiog8hYq8TyG3q7S5BxzfgI1UDEzThAF0scQ06SxU62XqPf
+jsZ9CTR2PgGgz9AUtwosrqU1R9n63IPr9PoBKjtBn7TGmBjKr/Bbi3zR/qZ4La+
yR+kb8N078Q8dExpkhIaSqbxkMmatFMysCInXsr95Sips+zM8li6sJv49sTq0Cw6
OAQi8aMPABhmfOfX6HYpClKonZg0BRJ16TfzCgjYbkMZbzzxC0vfjc2Igy3i/k6D
GrTlYI/E84uHnzQiauFRJSV8tAq6IB43F4cWLbrP41+orn/5OThp8QQiuRcECq4d
d9Q//m9M1zt6bC2z2eHO9bFZEUvRfC29ntE9PNljX8JldCIMFS0HZcGbgE/BA9T/
5pwdmzTKPKWmy9beXPvk54biTwEC1VJPV690gtE1ak/BR36EKUgNanIE7n/Y8vVX
NLZ3hnX6u7RstRYiERA+gUAETd4yB0T6XpuVhIKOEFxecI1WwStQr7AYIR3iozPC
YkZFGEl/UXtSziHdzcqRPIfwzd4YGHdHFpDLkYbacn+VLGaxeKjN7y1zmjlHdrE/
YzZLFRQgOch6v9kaltLf5xV+nzyfwDACBAowuJtXIuDsCflBqeuZBYbutSTpCsNw
B95JY1v2v5CP9H9Vznmc+tiVu7b+xJMgWw3hnAAQMnvKg0B+JjDiUwnnBwJUWeZu
WOtTYiMunKW3AxeCPLuzLLKuWCPCa6q+os2+5XNtil1dP0RebLQYmNEhAt7rqTtM
w6CVWeL71ojW7K+lEbS19PeLiu4EnoToXyeeQbRNgqI0yb8PHk6uLddwWbbOQO7S
Lh5EKn/JuF20UQG+9HbRR4sHW7rmtnaPs3+8qSW+R9lLoyOE+tRzloxHPSxMjlA/
CaYqsGxYl1QK3s0nA7hks3s2pdwdKu5WtLVdTfVEIItO3Pn17PoaMG/iv2ybFGx8
Efov0P33F6dkIczpgeGQcJ3V41cJjEKfuify7MFxcCCaHmJ6s7M+4WqmaRhK63R2
JiC590mNyjj/nae1GqaVSpW4USY3s3I4QaFdPKr5+0bMKRYVLS1A3Da+CiC6HZJS
2wqYpSSjbGNVBMVVYiFh2Ex1T1I1OxRKhBTh79kJ1z+z1kfcAvM8mzvSW0obx5et
YNjMsxpJxV2A0pA6pcCLxNm5ndrO+gkwUjKyfM/7DMi9UWw7lFz6UC+V678kCjYn
PT5ngXmuGD3KPlQYfpnEbw8D2tNrPsXJxGZ33GHHPiuEqtYkFyO16EkU5YOGXmWd
qps+mBp6xuhMe7aSkkFokl5HXcoBqBTBnWH5g6Pxq1lIfSyKYcE+/lb3ZXIfG9f6
Ic/pwlrt7OxnjKRg/+8VWfFDwoQhmCO5nAvOGADZMXgJ2a6U25VpWD3VrDC88EOa
ligjALAFIOlfL6rbUuchx3CLJg28HHBEE1lAykML9hoJy+TEGrbh5PnYWo3ArNpe
Cm6L4skApaLLNg0O9pKbXIS9FwFbS5mdkRbw9QWX/7OwhUXmKmZ2mZBuuC/LlP57
fo9x3VUXoI50Wt/q6/6y8QxFRtQoLWxO4LvySouaoCnQQmCKNWcyGglMdfQMHuxw
XrKMLy1CcW2hEUOvJUuY1PxwHRkXrPjLQNBCxYqb8TkxmnhC2J1++5+m1O2Y4ATt
OGKyGDc9ymUUlRtaD7obTCnCctqCeJuwUrHnIRu5gP+RwpDPlZuCovFtdhz+PENs
LY1HK7SAjOVDXyCa6FIHEtEqHx3jxCuabnjNJuDt59H9WNo/RuKsBxgM3RZKAc55
hvm16vqRuV25iJEZ+YvoLxmfxgI9IO9ot9uvCwsDMfCuW7u2tQ4KVVgCZw8JwPHG
bjBVP2HCju2qTjUTZbLVLLAcJ8hKBhWcuxR4LazvTtu7iAyijYxf69CuZzozSr4n
1gM+SA9rlmaFW7Er7acekpmpv2yWluDNg9YEao7LYJ03T1p2wfmeQiCu8K6dKLxF
ppmPqV+U2P6XrCSXU229YWsgcTr7z/bzkoQIp5ngoseBTc90RwVZAF3Lwh3N/Yem
zy7qD5WhtodmlPvGek/yfihAl2j+HGWzvxgL8Xkczoc1zY7wafmdfTxTLqlkpthi
C8PNc+CnEpL9zNoc77Jod0xYGzYkvcUn/x6cra6S/XqYjGYN0VdLkVHB+7O60BAw
8Vl7HxSG+rKUaK4DWVTywBpDTMFaoTvn5N/asc82Em0V5IE+4lQMXSWu64qT08/6
qYT8FhqWhZbOsTXNBH13baYLTYTKv/9+D74kSQMxSfJnS2kthxlDfH1Mbe1KASoW
OFx/Z4YeW816d0v8oqXhhnM1eYTG/JwSQyhOxjMGQJ5QxLnH1O8kjkvDKHAYU9qg
x/UHGOQAp+vblOJGX5qa0POfEka6F3nKlftxlYgvui4REFTREjdo6njYpuoFV/sI
0mr3n6buwMfU1nvQqpyNTjozF29Bgt1k260PrcsrMu2zB1RhSCCfDfYeizukwVns
xGsRL3nyu7Jn1eLGAjnkdwKqW2vx0T9PD4T9+NlfhoZZQVXevaK/F1pkoz3pfTQI
sgn4LT9qSjT3B55GNjp/s7O0r3pSnwo8VQkqQ7dtIzIcU4szYoQbs13jiIV1OtP5
IvhBBqUQp2ke/KrzuJAjvU7NNUDoum2Y6b/56WLD613qyxvQh5wcjD/kxdiHwx9f
w6y3pLHgjVdCeMQurLv8e18eEC8up006CuXIUYsFZ7bKfk2Evx9cUHN0QR4Vpa63
Q/6O9MXCasBbZqIZYya+y7pboKa7GaBvv8fzeD1Yt8MtC7sGKPEhD+xH9KRSTyBK
yYM3jA2kEM2FHnMkPOgXueY+BcStiHcArfSYsIKMKk2sg4tai7FDZg/lix1mehWV
RafvrMdfpPW1nyp3q8tpYYMtMWEiWbudidXW869h66ohythLpjsSHMKgBekWJGAv
NfDwQ9s+MPrmZUAOUPFqs8tg4SlJC9X5fyN7TVTRffqA3cuhKvlDPuLI+FMo4K9G
OEDMqyZSdNz/vwsAHJdVqIQ1MboYLBl6BErFgdk/aPwW3Cm83PgQSAgM0azHnmt+
E3e+wRntyW2dWi/VYP7Hmh8Rjlx/UTwb6HQPLROFQTwmV+NlssZI/lmTVqmmksPP
l+r3Lw8WGZJ+va23AGqtAYg6dJmQ20CnfAW6/xUgTRBGgvhvqMjkPvPIdUH7aSN/
ZUdR4lzjHDK4mM9acvJn5oERUkmqLF+4LO8I/Kvfiem95466BBMGn0BggXmNIa96
cgglhAtN+1k2KszWSVGd3NVn4d+Kc+pUjU/lFgbpDYXSRzAlZzyUBtcCXe8ir8Vi
DO7ZKUu7DNp35z1I2goiAsrrlalGiffFsNq9EHxwEz1kBwC32a9BTs9IpTLvP6iG
9AfSiG4rI8nWpmBBcITg7nRVbnpbXH4hbBNXC9BBSXEmyDsMhSLWeDZt6Peujk8d
0s1K7rpm0HsUtxdtoc1caS2+fNNTHUa1CWFLyJOmYNwB7TXpUmVJ0Hyxg3vzkF4t
VcYzMYhztZ2s6cGtNWdiLQE7Nm/NYVhNu4YYrWXRG1qn9piVBOtW1UT9ob6yImy7
xx3HsG7nxorf/LYw7K6K2KMslDrfPBluJMiSX+9Je6rqf/wjohDZR3xVoWlja9r0
/HgX+LoRisIw0C8nnDevz/bCur2X/Eu3vI405NELV/Uh1vIeQLKfqUkZ6qN9+BQ1
7VK9jQiVhcm9RL1Zb7J5Jk/YChdoIEjv6N2j0cTd8Waf9ZdW7WiPapbNt/vJvbpf
FhWQjgLlNkHNHJP5/FCONZBPaoAniu1XoMHRCpJR/3G3tSGkE/IdG0F9PUioCBVh
EYmUXle06ovZvTFxeQq+KNcmSqM+ZChGGDBIxDZICm3uSYo0fl/9V97VcuXclO1Y
N9HdDoNd/EsO66kY/lh0Zmih2uTigyd1lzy5xCc2g2+Nc5yKAGWkndKxuesIss/L
wuR/4irBV61FyrUA8kP12tF0752Gy2XNxgyyBEDr8Vy6fqRvXFjuDMWdMQwnm0Qb
XBUvUWZSrewXA3pBwt1YTKxoFYQCgn1fkMfKizMWxkduq+Mw6OUEPBUxNm9HiF8E
g8+fydyNWC73bzZKthZdw/tj+QVtxVypVXZl/WjSEELdriwW/3t9+xd1cByb6aPu
bc2NECMA6ykyR/+veLDg4FBcg+m1Nr+DcsLq6DS618KSFhsqWp0GP4E/8SJpBzCG
k5uohIe+uUWAaHTSdcPNqDtMXpHLsWp6iRnsvIs3qkcRNOF7dPKZRWrUPA5y/tcr
J+URjNNF+OzyWCAGPLyixSJ79Id3IOYWfp28lwnNfQC9VVr042Vf5TokB2XZn5CA
Ml7i8/SIonnlvEHG31ohBbew85yidmJ5dF7EgXmQdb93v4S35oef6N/aR4oi/NPW
fUzXJOKfjU5+87QR5JtZsVzW1TAVdgzle1gIx+ur8LD+S1cT2cwG8iEIO1knRAJF
DqUGz1rLV7k665qrGNfeKY1qjZE/boPqGix4vmz67VjS2a33ZKMO/LbvHGwZSpHP
ohEA/O1iAIvZkIRsgFIzo7unCRw+8Dxn20h4HRkOPoHi+LCNgRzLq2GvrZ8Gw8lO
Dhv6KTv4sZFGlO4sxVPXaCtQRcfU61TMEUmKNvZlMF81r/zEYBbapXTn51b9uP4v
IkyRpxgDOoEO+FrO7Syj5yZl4ubPVawp5mizZM24w8r7ir5ggxHxf14fXsc6Hhym
IMZI8CIYPK+HB5a8dgXcGqSDbyZl6dP3ntl/h8NU96jXET9C6/sLyV8igZwsYnNL
y7TlxRgSd6paIKycLH+0bFYTQyK62a29HPG2k+rat0jP8Av19kQohMyOJ74E1kGL
s137r4uSd5nTX8Cqmp/R+yCReiUJElt0sbHqIPNplvqYhGbcfz/3inxfAwuFyb9P
Yvt8SAVpNERiLSnPAWGoVgWp/jbLcyO5K90TkkmF3nyaCr9dMMkQ+PAB1HdGIhDI
g0/ooq5XSBTTCYRjn9ZxhtAHnM+nq2sd7Fdq9sl7V2LH6dF6hOOA9VJyf8NLHLx8
wNFxnDvc5V1Gz7l7JMqojX5OUPV3NonstSRErrPW0ei6WpaPuzjy3/DKH3D8luGh
uK8+ftxjOHqdVxqrrOhArCtYPzU43OT6X5BGCfCzpQFETBsNYsFIbNbhf4DfPYih
RkgPNx2l2HXdBSwL9Wi0VmGXpxpVl+iCc7QdsSvvpi2a4KhxPuCNHwwCoOvGOPHl
JjKlBfRHnClju+Hpp2bzrl2FcvpdGkBFL7bYemTixQJ6y4hNjPcwZfToaNmlvW8Z
eGFFWgJ7MnVvBOOJWh+ELhp0qUX2cWzvO9liOFy/YSGwQZsEDhZ8gwwWjF6eFsMz
kDQa4IwcyNl1xF7ncPMX7/pteEW7qKG458Z6/rt7rvXnaK4YfWKfO961P5xSEwq0
kMZhQ24keQuHBFqRX6nRXkaU2ANNi1qCKHvOw9SfcQ3ZmZelWaoX8/Wqv5BvaHcX
iLsQ/eCbWrFb4wI+MAN0zOQ6FFPZO1sxRTnytKceyk9PS3bxadgpOQjydf6POsiP
ylKpB/6o27COf6F2LBWp6/PpkJ1XtvhXuXpJHHdOWt9CXwCuJoLIXpfXI6aWUd9C
zQ92Oa0LlLZNO4IMMbkkabSMj2vEZBTrr7XmeGqbPJg/MzZa0xEZ9CeEEaPmXGyb
XUOalOKQPV10jpnCUfs2IeKu12GyEgHYWTpN9KzNo7JmWsMBlGM3b5zWnCSYkcmI
t1dDAmzBdBi/UyvBpOXjn3oVhiCikLz+lUcrlfZdLVHNruwM1pmxayWPwn0XrMpk
pE7fVJj6FnSbHTQDw1cwZW8helfWKTXtSuq1CcNE/9QCjsDDYNkosm38HAG0uhWo
UxI30Xi5YWEobPxa1ntxptkWvoKc64TL6Nl8DtCrydaCGjwzM5Gf8znO8cGwd0O1
RtRvexUiqMKa+bLeqo6HkyavjzFdoXPw9Bj+PGK/v1K2ni7Vh66IZLmvyO2i2saL
CBXHSM/DNXH1RdTlq0ExSu/dNCpszUtVxlNzHT0rXFm9DDIrIj4xHHD0/j1WI7Ou
CTLdPW+a+0npMhsB+zK/emf500jS2rfkdMo4QILVzmCLtyNiGzi2dJd9U/OuPchE
xamb8LFk8ko3yPvDueOPICwCaw6e9PgiHx5m0w6B/SJV7g/FnDiEAvzhCr58tE2P
MWm23tNc1lzlkC3M/6QY94xndB6bjxgBNUaMiehGnVQhIE+jet+ka6go59bXMHtA
3ThLn6nqTvw53/UwSubKVyFbvs2URo4VOBEMsGHXazgswfZQAIPMg3YoB1SbnqJn
3SjGTyLFELA5mVkiATte9A==
`protect end_protected