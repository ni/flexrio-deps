`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xsYj4ZwXcxl9cxOXlpzXHdq61odkffdZ8M8+q+kFVwV9XB9LU3CGsyRI5FIQN1t+
80m/BnHSrgptdOUztVIRaN0HaBi6KntDN54vYaUjNslgNp50Q0SQ+wMHBoxBRO7K
aBocoIKu2JVaYvKTGfoe3Dyix7uGXReNtXk4RqoZYtoJ7Lj1EcLUs2K6v0+GJncQ
lcRdnEFDYaYFCTbuR1NWdr4zj7cnpqc6LcEUIoi5XPediwNYNE56bldepcgSE3kq
rk1nO54ixjCLbzjKfdFCRREULZUGPOpfsCL2vxyZeQZXXyTSTG1NkG656lYcCskj
vk2az8bCgvKs0t3Wths2EE3LUEMciSao8tUOIS0oDegx/U7FX/AVBf4OOb/Xfyhx
vzYEVePsfdRPRttPICUjbahuNbVXxuNeZ6dzx+aNI1SgRW+qjzFRpESaetkbE+dy
VRH218CZ1Szj+S0DvXeBh98ZP3TU5ZiTCc3b1eYfQxDJxsON1Ff8r8fx/9S9vPQp
DFjez5n69zNawPo15hiIw4AAT42Pi3WFo7JkRTMVlW+SbcJp8T1oRmjYLp0UgbNE
6NVL6sQWCRsK3tL3r2gFZ4BXMXl5LXoUnWGdAmnVqTFZZbXlNlf5bj8rQGXhgtD8
Wuwwez5O9vZ9vO3Hn1E0AttJHv3Op3qwvgTIHfdKQT9/qG6uTWNcWvus10/Turbq
RRIypa3pOjZD6IfK8pxCuoYCjQ1byNwSOJ6UkrshwUP9Gdqc2Jy3TLKuTnU1fyE/
BY2ANxAbkzfLhCtLuP8de1gkjLQGtdbNniGtRsWOJlEd4aHT+p4scmjDRYmcb/FH
Z/YWxAn3WDJfrA2zQuAVIDE94SfuDQNn7IU3uUtEVQZdFSy6+DjY49fR00tocAFG
23YHYkA7P4x8xkhP/CyrFa8jlA7grfsr4KXGvcPWDFatclDvLmPSZuc4YutI50LE
ryfO53YtprF8uIR2kzeXPfa/8b7wEHmbyGHSy+cGqNwxYydl5YICyZ3uFNgcjSwM
C/tNmXvNzHq8LvjieCIZ4TYefKxCZ45/D1zcMyZJShoS+QwOkVR2g5cwSD3J1FQn
2y/SQSEmOZ95J9AayNAsNKPk0yC0ZwRS6B0dyKdx205Wkrb/uvhcDA6bNbQoFeL1
xSIYGNOWmaONejjDxwE6lUWLSidRrN2CaJcQtsrx40PKCcyw7sjyQyAbp4N3bYkm
XfaPUlIZaZ6X6i2OPS4hQci7bGCWadZFcumzCoWmevRenMVy0COMsws/WbkvLIM7
uvhRELGabWmY0K4zmZtoXMCFlUAy51Lrh7ikvzU/nO1I4rsD5YM2leAfVuADPVbC
9Yd+Fe8NOXityAjkfrDRY9PJDpIW18nbuJhy9wU5RiKXkadFnSnOi47qDAoicD5h
ZNB/ZK20v/X8AQKKvDvwk58EGPGgwg95bTshiilrYd+n9GFn/suWG6pKxIeQCpoh
se7Nk6vkMHTy0Iry/AXH9NYiqIL05x/uqZZkP8LF1wDV11VcY8mTeyUHrTk7Y7Gv
2z/0lJiQnxG8Gwx7T2AmAeC1KuJxVRyFwZDFNT4BPwl7e+cW+ohkDFJqV4gI8nI/
ACOJM6QP7WKc+HKAbikOE5+g6Z3+7Ca8pAP17goiO80jptq4tSIyKRvgYpcNEgo0
7zYahCSvO8ZSLdFxGX9dqj/Q1+UIVtD+ZY8ctzB/muls7CHr5m4PNH2JIdFosmqf
4XMX/sYE5drEhICgJ9zwkvX0fKU2harBsl7SQyAtkIaksikz5y4AsqvNMizm4xpi
7liS+LMjszcjXyUtaZ+ySCTaRJlFMct/zqDAnfyVjrSY1/5ts8eUGhV2JZPuLPc7
RLAlGipyaUBgtcnPt1EwK6AsG4am7I4kewcXQidJqLu+Cz2RkVbY88mEzlirGk1g
/LJpfJgp2Dls4/L+IcarewKc3KGAsy8/OLYOomHjqnViD9NfIypgnA5U1lJJLVHR
9w219QBpxD5VrKT7S4A9fmEnpjV//YdK5BQ2eb2ZSU1HcoX9Y4oiUv8MNVUyNioN
2cPhv2vco1KqXLKXHNePeGRL03uQssm9LbqMk3NEmR1ClVB6B2f7j1txtmjYN208
PmvB9rzQufqmZGFXtAkVIROR9xzAFUnJymQ0HyMVvxY=
`protect end_protected