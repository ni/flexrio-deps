`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
JfUWfeA+KKoJK56uw0JKy/zgsvZQYVYrxUut37zFLYCBOzRS6+SDis+HF9vVFRkt
07aSrmGTcxtdJSn3UCIk9pzs7N5rvfJEb0i1skoptc0TDD4mtWbj64Q2sY1Wnmj/
q5TwtV6gF2/2cuyWDq6yOniPD6h2rxuqfCjuaD0G//syvBKJ8Iq1Twy5RAfg/ojI
K7zaSnGFwUZ0S9BYeVH8gp0W9+hj4cYwfCMB6H4Wcw8co1mErmm1Jk+bB3RgSyY2
NYX/uO/yY3HXGmLA2lxuxwLgvgqYdKNrnuYjz109nJFQdZPrgwx0pCUPS/rWrIS/
7xWsU4V4L79gWnURuX0OGkF7rg6HqohsDiuPAN+x/Ul1clFeGR8GgXLyaSc1Y5mw
cEwvfQef4x8KRfoMYk0tC3tXgLj6ap/cEWFnebsNdJCezm4qJOVlrKoRmcQP2Pqm
vkByNpvC5kjzPxC+Q3jVZsRNSK9L/el0BWqwN+V9ZANP41FXaNDx/8/Uv0chFdEP
+A/lr0QV/0KxfN94w+Glh2xKSyDes/U1xzINOngW+rIgbu5x2Xi310R1HMkIKN1S
X1kR0gZe2l1dJFcHxHI2I9uXw1vN55npwDpQo8aOk6cL4vHUDTjyDrIkQ3fK1WMh
swWMHLe7nshxpZgjBXe4ScB51VYvkM8KDbbrabfBPORsQ9Er7Qye8EeAI8R34HIi
CkJectZdVFAA7MjXEldnp1JB9gEeJ5XAkFXHsesC1IwgGOGdGseVk0QcK3Uh0K/4
OX5eOdqc0UXj1LplYHey5KWWhJAwxRd5ItFyVEBetJy5I4BNW+pm2UPSMZVv6M1F
KoaUQGydFXlLRz3ZGUdIunnVF/iGO5FICVB3URjyK6FMd1flnLfRpMoOWTy/07jk
f7J+HldxH3KGRmcB8VDocaD7t7HtRrtcY0ZtF1/rqUWuBWcna2fziVZXlT2ieSLe
1/ULHc2wWKaJP2TivsL7bgxkQJgGub001pS+Ds2zGyPxbd+tXmdz86xeUpwMsBBh
DelZ0l/oecHZw6OJVlqUKezCEp6wTm1HHRFE485Xd6dXTh7tx5qIf/3z47AdsIP1
AJtf7EsRK1OxtKjwcYGptsBgVO3I0m2onezTn0aRxdhjnxvdoc5q2HA8HlufVZRr
JVN5veEwlSL36bWcuOCInKe8gOhmhYsGFa2ctPWxLM8N0UNI7cRbat5zypa+6O43
oC1rrG+1ADiFlqtzDZCi56R3GWqdSihBYyOLFabsvZtTSkBIZeXgQKTYTroFWAIh
GfinKug8kMBe0M/jNeqEaeq7FgfAvxtcdNlGQOKslqSH0ayZ5o6lEdZCsLY5SqRd
Rv8NEI7rtmJ7KzwLzdO1/mtVfbr+cyX1wCRqNZbWe3F2VU7fubzG4xwyySIBOLYS
KmrQRULyjvD78XgS/w3N9ewXa0jHeA4FyiBtcY1XuLLlu0VJURd9fPXUcLBxiAd6
bvzkJQmij7xuKRXFDXNU/vPH9tDgWys0Bfm5nZM2Dg/epSOQvrAtNT3viAr3kncE
XuPwRqfgsEa+vEgDr60vyIbCOEhQvw+kVxglg6NRlEqmD+uDxTfg7Ib81ZphzaX9
qDS+tVcYfyBC4uw4QJWg9CRF/hAF9OCAmeF8UWhF0xnoZE8s6Uoa5AUzXCP/ju2M
aH1V6iLW3BSMXlrLQxmo5F5KH0Pr3rIewTzHsSLiiczgCRYa+8BVzVBSrFhCxRTV
0xAk1EBgSuk8HPRR4ZIbaPTvaGlx5QLsEDOjOi5Z/kOV2qZp5y13PCFDlyGU9Q0N
O+CD4sBaho69dC6iOgY54Ce3D9uFwbmgiUFzzTcuSTZafnEuGeJB6ngogK0w+sfn
j6o/+lo5wYrqr78cTXlpV2HH5vnGp17Rj546cO4CT3OLEVVkGWqTDTZoPy1bQwff
W2bTQYYJpChX5eK9/+SPQHPmsuXeNoQhcfKYi294BETG65YuljJpyOTJTJNrulT0
+frg90mVbWvJXkGN3TkpDZClTjvYUGE98ZHl8maWjsfHrNMj0ZrKFFnJhP4l883a
eQx/JoUNNamlLP8ISLzhLkBs8a1BpK7mZnjF29sDIbFsS/3ZQGXnS3QFcaXXZ997
AzHjQWiDXGHpaz3Cthx1+hXeWVAu+nsLhSryGr7n9NHcx8xQcmqhT0JGTgnSANhs
92H331Bt4Y3cLX/vS/RyVeIWBNZlCf8dXajr1SuSS/LDPHjToGFjXHp3BxrA8tX8
4P2DKJW8ID4T27xKJAizIQtseqr4MFW+Y/aK49+CJhv8z/xKQyQH7+amyOoJy6c9
/e9y28ZlwsY4+c4xiPVoPlfxBKakEokOX1DtSznwOKybN5CC2K9SgHwT16nvi9nR
H44FDlaDKMxJSy9tomFlcIVqrH9SvU1vrK9UR9W+BvwNoxqJhyvPdcvZWPIG7TLl
JabLxVLt0/kDx1ahnAKwVVgD2kRCLBdyoAJig5iewERNam7e9HgHIiufO7mq/VG/
EcbdBztwbTfks82t3JfpcKHxhcU9C56FBRkXImRBkj8PpyO0LUY2X1cSbBsFFojC
9HpBktq2hxjpj+artnVtqnwn4FHriAJm/pecDFapAPmyI+qTparvFVm3sAZ+pZ7b
qJRu2IcFumNCmqdB5BilK4TY7zWs52ucG3sxu+v+5mMwVlIil5pMC5J6FdZyTTUl
rur0wTVlGF56znhuX8wIQPf7ubrOoReadS82XQQ14mgVopp6KVUVDpnZyLxWOT+4
O4dwbBLNPcc+MoExXQZs4O/8cso75sWzvCABsP99j1fehWRruU8wo6/296JeOf0n
8lU9+tQdUQblbgrk3Xu5oyRXBd4KF6CE/RCZiD1h+3uffWbeFamDCFg6gtQBpKMt
JbuunHj4HqP7acjbdagXMO/TDPuBlRbMErrGoiR/pApmZpzpF4p2jubZR5UOD/qh
tpVa/DdDnfnIcVgQqHJLep6WTmCtQzS63v72SXltu81sS9rNbJrof6BID1R0gxgq
tYQtICwB82JLxCupjuumRzAep+tMIPPwQ1VRCOG4oenibw1X0OSsqL5Jnw/+zTcR
9sFoe5VaoxwYIuzIqSK5pSA01IZiFFnO1hbezQWnxJDaCNFF8f2AmCkJd2mQ+tFC
fNIDn8B6pYCBTlXc256viCR3RBFiEBOGr9p3ZoNWn+UuadT51ipZ3UgaGxW1CIeP
bWk6YYlOObaId6D3Sq+Uiff0XJSebUaqqcfmg4FB6TpbmIPMnNkkZT5+yX8XE2U7
HzfG+pQNhUwk1CyBIlMMptzuVJ68uzwxg67aYV0yoSYBW/M83QjgwaiolwKnjDOf
nGhPFUmYIObn7h89gDXlz51Pt1wBe7WXZGDTVDITjTEQDRW0G2BTKALjIJwP0gTL
D8j4bHJYk9jTjm5TFwoB+JldjfJdPpM5NIQZJCXXGhbymTi0iaEvBnSwPzZHKYwL
DujXIBcbmZd1etgu1At6HUEQy6OC9JUU4Gl8wkvMHVnXbkmPuQ4rgO0DTX7IUA2t
mw2C/BjdGQv85Phz/v6WbKZctsVQDvoBhmB0FEBkGD4TJBpIGMdIyq08CRuScajs
1xqIpvr7aYEdQEzDI/EXaxsGwHvYWYGSXfecAFD4/J6xgIVqhc3LAMfMukF5qL7g
DG9WSJrjflsMWztJQLRqfvnB/JsC1GxGcYS7AecLm0onYzEZbahM+xR6W9r6pZ7F
eifjLP5Ujculic6CGhGd3haa+HlrOGyq7p8wC8nJ601qDALSR+K/HtOsw10dIJey
pH8H9OwoTivgyYGmAZdB6onT1+kHi21+VMls1S7a+ghgKDXlvenJUwhRYqjUSNr4
EJtSl0Th7djz5/gwC3qPVCEX2Xh7+MT46ot3CqOSuQ1cAvDREUetxZShUlFoCzOy
fyupKeNjhVIuqv6oXffvvYM552+P0qBrvtEjyYRKyQTBFemBNI6NIr8TpjCjGkP+
alfoPHvffx1vxnQlTt9BI5loZSMufS6ZM4TDsFJnsI75aBC+OyKmI0B1MXX9Hrur
s4bsgB7bGB0xBRNjy+VneZ74jGDFCJ6wfvxNrDbo5iro8B618Cc2EdQNZXXsvXt2
nDagfmpJnYaX5mpEbW73ZUnR64J9bpLK/ttOVQRadU7vx6Ass+mO5SNvmusof1K7
V2pGBaDPjRE4yeP5+hFKcalOobJoZdiOUQ8dK1RDDEByrkQMi0eqvaihzKyVZB9I
5OHIQWBz6y82Ipe8KYWTjnJcur/J7cqU/QSTg1ZR7knyawbXhBVxyRLPbrubnpxm
80OaR6E9LIC1r262G0Cfm8g5LRWtQFx63fC8kVA9VLaixo0fDVbqNhYJNwgIKf4l
CC+Kh7wZA2ehMTWtmC/uBfCF2azoyf2YCLh1TgdnVK/Bci1SbsHwsMuijkxiYm94
cR8JCBvoYJ3G4/gnOU2vWG/aqIhzjyaYfVj0K6gujd4J1VBEoNq6DhHrT1Jj50D1
DP83FIB7xYjPScnN66YgRhiIAT27x4oNPR4Ji+vosJ9caq0iizmknUrBx8tfvrmW
h1ffx/hdpTzWB8zTY9wx6yqlX7yG5APoLfXMfAPL0SmyAJvUidE7GzVuqscvsUoH
6Qv3UJ4w3OS7uLXoU0VLu2ZqTXfn78oi16mwtMB0MZUOCvIgj8t4G2J/2TvCevST
2Ff77fCrt53ICb4FjH0+0Dldc1XY+dkPNoYUeqjCf6NA1gugichZc0lV6gWqoFbz
BOHkA5JYsLnjHl9Ii+MeiD23xntttBkl3h0MCccesymGs4mWsTThPueOfrqSLQ3R
DtkDMbN9jACJyUX/AvYUj9n7mmlBvFn4ivrOO0ObGd+vZ8iKctcKVDKdIq3oYyLI
ChztyCbEY6VAVj6QOTTWQ3axwzseRG9X3w4Hq/q8SH2452ERiZ3zGQ0F0YjjFAdp
av0yiaXpsnEhcmtRMlUFwrKIwFMETytr8E2joqDnPXzB/OzTFiRNclSc5sJdW5ht
VV6VcJcqvrRdi3z8sseK514I/8VLR7aIvQtFaoDc08u2dDRGcMiyV/w3+WpERioT
jGZkBiwrJ02a7Eb5JwRmCERymi8TSEErJclTsCXkyaKFBdIZ0oq08MKqn8GZcOv0
CysW0TGXKtiDzLpBXy5tCohbKiZloigp4yHqYdLkFarTzTUPv3YhBn47xQGgRiuz
ErZs0mNrjHkuT6y1Av/vQojnRzLSFVXx2jpdLgv5u7peQcOpoFi7Lbi3+LvILqus
h8CDO2Cb0xX5H3ogh+qs4uCz5atdJfziw80j2ukPgB7JZOUbb4mNE7yMmWyiNoK7
OdMNaewY9WV+uncKA17dUz0uj2RnhpqcjXBRrrVLk8bEDGpK6eAPHGUKlQppjLEm
eV9Gw8o9wLEqwP7c+lPlP5F5tCn4fY1r/xI+RJA1MJXnPVeO+12gVpGJmwJ2ZreQ
99fff9pp423lcmOXSp+afdEef+nqxMHrCDbkOCWnZCBNdzlCj/+2s2RlkMbiFn0V
/GzrhF0QzOm7gO90ggC2z0BUIpigJU9BwmjzgRVjRYcHZaHzjHH1WkN/4UgWNNV0
EQS0P4oScdzQ1HJEUOS0reOwCNQfH54RN7iBaYYGJ5HrQOQjHLlICmGyYw0ah2le
aU3vVVvTXkfORrJub4UzxPaaRVNDTzkYOeTcstos48SWcjsjAfZrW89cVDDNJFQy
l39YwYvaDWt8Za0yoQeN9kSi3hW1lTZ5iUjkTr5pR1EgZ6YFGdJWGjmGK75x0maF
Mn/Z/cWmYN/nLCijl/WB+faNQEskHjGspydfZhZSlILMPeBP4Ey+VyPTIIAs5NHL
AODXhx5HFn2kXW7Il3Q2GYwixkObQxuWLC84Q8HwfsT6MeLwXMKX+cFik4b2KkoG
5Fk3w89fJJcqWm+Wo2SlrmQzWckQOR/+wCuk7P6Cgfe/hl05UF7cENZnXJxuGgoV
5+lHw95ke0ul82+EJHwffqwELnVi5z2R1dFrh8CdtPmCVf+7S0P/+ao4VXjBaA1v
2IjcSstdzp9aibYBtvAMgG8aFpXKy/odj8tDp9W/e1nK8OD76Nqeu9mMRxzpgIJh
2wbUFRWSRKWwnF+42Q0otI7Ep78gkmnjcHXvpQmb5gwm/+2f0nqG/ZIHHYOgU4yq
N6ToAIZN83cULe5xyVTqhmZSc9hOdRN6JMFEiLadQtV68aSVUjBBv2nqw9OU4XfC
VHdxCPidgylxgz1SbgkYquiPjaKq59GsdlL8ba9HVk5Q4bvgQdRH2xfew/GoUVDp
GBG7Hp0/YsHc+NRHD41F/P0NhNjBudEyIVRuc8FIYaoAp2A10Wdpq+qPTj2CifCX
Y8qjrzXoC8whcaOKU/Mw+9vjUaxevaecFRbdy45yunrKBA9/RUrB79ItCnt0hjws
Qt9s7VA8cPYjA4TjmDZs4o2mX+ifcPOy4AgeT6ld6tfMNSl9y+Z5L7SickupiHGk
ca0e8Eh8SJEBYdCJZT3bDrxgK+NhjW3bGKRov2mOozUv8ghC2jMZvIZ6Yhulv8cY
aEPLlneIUFxelNXHbkxVDxGU+hwP9i6nkszIFLNogXekgELrIAM6a0Vb/D4iQoxe
G5DtyDm0OQzvMAvBKjtQh7fE6GK72uLxEqVkU8We6p6acNGXb0xTvh0fZ3xwvMA2
7IZ/AcxDRHlp2SOOj54Ex2idJ8iB62DGiKftpF/uNFoJK5ioDOkg0LRlrJBiiK97
+dVb9Ldt2UWVD56se7uGtd0paE9GSIXU9Bv53QE75bYvOKBDqq9fn3X23wrhH6P4
zKLS2RWvHoaZgsKgYzkcXn+dEeanhMojHPPiVSL/9GcG8bcWktJdewrKgxBThrEr
H4tslxblchyoR842g6Ok1TddRNSjgjfVxtkMlNfq95Hlk0U2ye1Z02U+txh3UIZq
gyQ/4Tvoyc0K30kycsiRwJeY/DyQkVZSixBEBO3G/HVvwVwIhup0CIUNkBQifiv5
ZhxifllRbQQjNcmFwVBHGVgmGXMF6cBXjPBnxUAEfiYqmNJiv0gDNhbDdSdgMoFf
vCNDM44rlZ1WY7V/7AjyosDAL0gdEFsYSI1HweHuY2JLy7VyNxqILx4EU5a9ZmMH
ARrkAdygE6xdhDnb/EWYZ/dPFtli2eZg8+LErm0r9f5FfUcBFbBad/CR2wOWWKHy
dV5G5gClQbkfjsBJeyaQjsgTuMlKfVlnKKSxTka1QqNB/0rOBrlDOw8/LwEasPPe
MFr20Ksa2MdYqKxHmCgqnAccmfYIYMayGo2qe5xYUGFwxtumgAMbXmdC76ymMP2I
964Q+D4Lx1qcm5rWhul2Fnbv7TNOtCPv1+IMwq4mjZgj7mpQuCghFg5QReLxRRaV
QeydqcH3JNsYNqlhf9JFfP46kd/glDFbNcZNTRbM6d9RGNS7emQCMLTD2d4zcnfg
wJ2ljX1Dq/tTcyc6UzzuHlQ71ixu+z2xLwhjKhLl+LX08pFQYriH/xYuyO49qmk7
UK71039trDuaqip+QSUXsnkOWm7EjHdb3zEAjB8tM2eqlvHdSNHDnwDvrm62DaBI
t3qtZW49vlzKV1GiuGHY1qNn81soPLNNQP+DWLapxDdP+tQ5MwfDOo7ay0WNyWEs
gPwoMUcxXaUqMqYq8a6wF/aa0zDP6/+HWKa/mI2oD2oHwBrAKTlmDt571abAXB4X
ft4GBYkVc+pldNShtsgHUDk90dPBOrI3xyNtG94mbitOn0K6WozEGA+ScjuMHoaS
eLybmDJOGbM+Eg9xq2j0wkkN77KQgQXZwySQjcXYRC0/tONsurpSTTvDT3aJJD8N
8cLGmXrj/yG1Yaj2wI2A36wDaaL6Wryiw60+pRrmibfFRiVzBzAisoPXX/AQFXgZ
VXpIYXmQG0g5QDrQUGUI+Q5/RZu/VqgW6pQM8dbqsQgkhqalatn5H4L6fo6TdJmS
cLCLoJGyVW/6WK3WhFZIb4+EtaarE2Gi2XsaYk2tPKhNL8huMjc2mSpJml3ddEMo
aNNd8mgKU93PvXMFTRCsxV9ex59UHIbA5Lo8raMW3MHINKzB3LxrWg64lUhHtBkL
ZtLkpLGi4tbshINghUxHggEfoDT33QT1rdcui997G7SUSRS/lGyhsnSikTWF1+q1
dSTabk0DLwx685o7j9SCHabAf86h7rFTnSOET+ipnJYk56bhSEQw9tknDIP3uk/0
IBDp5ho1Wv8ErryU2uiqi8phad1X3WyCDKMBBYEv2YzWW05UammUdpCXpJDH1JbA
YROxkGcdsEuuZsDPlrbJ9rIVRkMr7yceTwb3NXsPuHGzK7OgK0VXpVjgGP72RtGt
ZUPPmGlM291V8oIDYN3sHeCHvIUNuNxlC3AzjvlhKzFxiLHDtfgqgUE5obr44wX4
xkfyDa9rN9mkKbMo/6BoMuTBDxBkmuciyrQ0XkBPkckRVdUlPfCpNY3uG6xNKh0W
r+tmljUN6UMFae0WRDdgsZPzKSAK5PEp0kbMF1j3itkRqjfnIkSpLccu+UOqpDJY
yw35mMzoKaDpB51m3fZXp3B9wDFI/x0MEODTQsob1Jy0dU1wGn0FzrGhw868o/H7
lz5VM39rGUvyuqmX/U7yb9Olq3ZsH+eYagE7uBOnu3PqEs3UgGEKQJ1Is1hlvNpK
pfy8H4Aw9JuQCEdWPWUzqT73woUayloTA0fbz5wla/31Iu7CiH/pJNwDKKkX5Mo3
bizoVvFVht5+bZDMV1tjfRuZ7Chl4djCGmZN7oSN9Y2067nYYees7VF+vjE+1eoE
PeEj7CGWFPWjMwYsWauq1Ao1ZgBZWyJ7v18kBGn8RwU4GP+KHMwmg+LKCSva/bmV
F65e54q8r6S4MtQheYWvj/ONUQbYXHiA1JC7TSdmRL9YcEW3CT+Ss+7/84TTGoQ6
vobcB4Ekq4Rtkr7esZdmOhqFjpyCUXnZhI+UQuDYPeD+KXHHZwZRWcUw3ZNzKddE
cHX6JDhoQQFo0tPaGydYdn4pOZjDSINuc/H7OqdGaVIr4mKDVcZ38g33Z0dbu36J
FcEPIIJ7j8V31yPS7xouunc9Npyxlc9v79xyDeZ0L/tUt+mXZvmAU5xAhkSdCzW+
F2IcshggAgOXWNeMCQLuswf27mLTAcUrrM7TJqnfqUquhT0breqWCoUQunpp4qVX
ZFhXowPG3NYOnAUc4BZfj9sW4nCGsiT/dCdpcQAfv0Bcjv9hhHz9wyE700DP1vX/
aweiNdW3kgx4VVWw1m1I4G6hCg3vUimnAuncYka3OVYqaofd5CTjNldTzS3uXtwF
rCLC0ppWhqo/GZbeFN2iYN6+0NLjjnEUDUW96LKe21KCClxHfI6o+/2cY3fur31c
3f/1XQwUdDgvvP/33hAt05PQJ/u1/NsfSKt5HOKD9oNOhwejAeFrdVOeM1II2fXI
pmUlxqHx+u1+gleSVs58tRQs4CKRX2094Nh1ZPCHfrOaOsh31sYqTlAYNX4oPSW+
0/o5usOSthoy+pQ3iQbAWAOA7VwDu2HwQj0ztFm92mKRSKc4vlyk79lcilHgHv8Q
2xlzF2gqfYQ9U6lou8FaojkQgbeTvbV3hmeF04bI2sg85JbuB2QM4knZsVXJWBul
nomaTgDsBZvBeVm4JlMmqQ3v+DSBjoOPqZ5Jn/Z2Avtu70DB0Aw9qU+zKNTU3kD3
lthuSSn5W2GkwOE+s9p5NkUxrHP1JdnqgdaHvAlqHTwL50RIkFuu3UbbKJ9xtynh
Ms2MDnObY1GhvAT4UFi6DUUv2aRe2WKrS3Ig8H588I1maEExKPp/keCH0tCddhIQ
rvxH52x5mqn87m1K0UsnlnLOyKQdZ26jWWrZeW75S8Uk+iOuK94HKGiB0owsn8Qy
eSXAhAlde3UFarL5Tu7fbT9oHmcK4T8EM8T8Wr3s68+WHQGQguzFgAzCsjm0SJRc
pjcZUSbRCfK4OX1mITQHXkY5Rqrq83J13Im/EQFrZDAA7Ofa898WSHlDAY3Vvw+8
sqgYcVYGf5+aUUKuhYq9JVykeyObzZnoyxVOM1wqx8gqxvdZVV84pIqr2LnakxsF
PKgWv2lcGyQ7mJd6HU6JdpKRf2/LG9urLe0jg3nwh5dkFgU+PessF4frraa5WCGW
Snq9T9sORbpwQxFxJ4oTGhDEx3wjQJVI8jTCJwJCv4OKx3SVegPLnkScu6QS/Hcf
8AVeGzoi/Abn3bLoRCP7IwSRFCUWqX0sAdvVSzBe4AePv6AvKJ1VPKqgSxsNT61N
N09jY3kYJfScRVamHlgPL5dH+TtahpSzmuPVoaQEsa+xpED+skGdJtNbmt6AXY/o
Yga+ICrGwbCjYS3H65rfdlew4jIm0CQFQVZoncSj/qINY6FZN5VlMwQZ20CNmQMd
IyPVPMeOmER/8YjcJODFXTWGO0W77hGopvwU/Z/iRAYiy4mT221Uulty37wTNCnr
VPN9a6StSNjOA2sS9vtWjXxtg1M1iEJ2pWf9ObrBXKKi2ts3WINXlyIZ0SkC7nXb
FxHSbFPdkgnoiQvtcemG2SpKx0SkXqkPy6pnPcls/c47n56jvLa6V8POLsU+DzE0
hHfzNkUSwGBKTkDmo0XqoKklDqCpx8V20exoO1pIGYC7sLEInKmyMROU6CRzp2GF
I634K9juzSZAJQ2hml+cH7NdpgQtV9bmY0RU/UCl+fwelWoXWi32RVKaDZreJqYS
oxfSv6Q2fMr28WALHYTt/LDebE+ptBiFULEiwF7SPuidHPUM0p6kRuoIqs7fkalQ
K2RrDqMKFAdGyTHTdYFWvPpE1PlmX+fMvcofrhhoWYcQjPNapj5rRUQ0MemssNqF
oRqXoGxMeZv1o9xEx0qhzDIr1uLsUenXozQu5eDYOve1FNM++N0VlczLk5JotqVX
ud4OS5o1tyFuUVvMmWRZqe+uZ8Ny6RVFwFJTuNx5mlSrwIdHNoaWFHyH0pHcic2y
ldHNyGG8PAjSTUOhOVYZYEiTrHR3pjdk2ckclLzKyELGLn8xBcjd3ph4+EXbilxz
AYQ2qQrMtBPyZDceTH6GQOTBLR4UzrQAlXrLUTdO+OopOKfkPD7N+p9SJlJuuq6l
sKFftPSA9pCynEv4ubJ6d2E2W5+kS0m/A3imtj9ORwgEpMxgyXg2z0FKr0xo9do+
uMLLLrLGFGBRvhd6Muh7AJbJsdgnyqDqohDiOFtuwNqscX+AUVKnBQ4Gt27hvsCG
265uqOYznozQsyfrWHob8FIidGnACTYVkTGwWr5XdOsVbPrXHI1c4jso0uovXrEJ
ojiaKPDq/d9TKVe+kRbkDZpo1jn0GSB3ixA4fpBkUC96dpPSORddhku+jg2RGCz6
JtaP4dd7+4g6dCx1sR0YGJSnE7yTyj/ICHfmoMcVF/hEyKjOJP5MF6IL4V1fzBkH
e5wI0FAxbp07jomoCozRR+au32D6eo1lJtBCNiLvuHHer6uLcewRH55jHfoZecq0
yncIZHw0fqhEqbwI2CYf8WKOQtAFxOZ65XXmWiivUmJoEe15A7tv5i13dHEATS/P
PvEDcYFZaXalkY4U4cZpEwaj8rosH5/H8cO8gFuMXt+JadbPO6ak6m4o4lK9kULZ
gi6UbiTEdpI861qzeEqMggxXrB4GrlYReU864ffxhUY/O6nBI8icDmUzLT/x1zLm
FwWwJg59/FQNMTVt0OfDormzGAi5UP0q0lDcU+BZX/mEJ5cWvQvZQCPt3H5MqDym
k+WJgzi+XJ3FM1S6/4pBHKkCdO0+2H4KsdhzfCoZ4zpzO2OaVUr/BaTtQZb9mb+6
VJgAVadbZ9VtbEThd101nhp7AqKPLLJ0t6asHNNEJ79yS3Q7dEa8HeY3C89mFbYi
6ymGptytPpY03Cn0+LGdPPfhS+xFNWQHBHl+wg2+Gj7MMkML8FAkeJBHeMfy+3rX
3oHCsAcx1JeiepB5iDd7+GKgLTbPuFsfUwkQyTLjV9MepTh/RWNMJDbue0sVyxPS
FWrlwEBiWKhxSToeuKMtOZNSE4rQOw5j6mqc2fU5dUxe/6Peu2bm1+XdMknEXI1I
zc0aWLqW628AMUbDDhjPyEIXWpAO02VF4YQL1YXFQoeuHJZRatOVSAwneERAaiUv
QRdPbK9Y1vQ7Tzu/St76zlBv+R5y7owe3wn88IeKOx023XHv8gIF1pPzwtiWiPLt
STkC/d4389m8WXclS5hsHFz9QjIbYDQnYCciYtaAXtaS4ydDztGWxA8Kq604ux9g
kp1QZvwJjqhLx6jz8bfdsqoycmZYNFrEt5lCHRY3G4hygsVlPQW+PVAe+U5oMlBs
xXyi2oN7c5YTn0QvGcl9Xq+FImnd7hZjHSgsExURGXlSff1vGuOW2Z4OzGRiMSGQ
FmDtUmFr5QZfj9irdBa083mG+a6WzgDhRdeBpRlXZU056zmCHZM4QlE4L4rggq+d
TACccR1KgzbQd2hXzBdZSCUBB2uWutDQtScYYaOoveYLWJuDcSa6ZBP/jcn5qSIf
AVGt50w/VrDcJTRWb7N0ioT8IoH8WsG9w7imu890cwfkBowgbWY07CzUViZZ/Tvi
6sN8AKbUhPc/xWsASG5xBHomLM7X3ZIJuAoXu1AxEwWRE4Mo2r1Yvun5a1rs4nfc
6yGiXwgsUEJv6Cx/fGswe9FPw/noi6ZKYix+r9csokHv6NhWUKCZSkOxu4+hVEvP
kueiI96VxWyDlZx37LBqa/cDg1WalNc7uDZGQGUXTRpK2TG3BRKLxS3kMOeoWr6R
2UgVC6gfFp8xtrAvblH85VGc0W++/znTYcChxVGlwKMvquRPTPwdJwpRq++Cuc8D
G6CmIZlR4YOtptSdvR+Ns1P2cox/mgwVYKgqWHwZcOU/vVtvsR75A2R2vgqP3FSk
F2QxTlJSy7riFjFuWAIAAooq+c6qRkPZj9s3Di0RCgKePRccMTOSd8hIAIOuQEo/
+kIpOebJF4y9aTzFAT5u+krk31+pmtKNy5TQYNl+JHdsPk4DJo2aSxOW5jalHHYX
kEzc0wq/A4I11Sy7mPCKqmdkdCXF3S21SWaEa/7Y9IX60DN/VFvqAx0PASIIqgTj
C75Vm/dnxOWvWY5B+ingMTKfWfuW6KtOFrknoMrIzvQtr21UXoIAKkVeKgnZG45a
U6j3Xh6C6dDfKKvU53GgZLxgZ2/tvKvgnqEl+IfCOTuFgSZzlg8omOj9BKxyrmyl
DP2tq4OfBOjSjXF2L7u25OMkrta//X90AzOVL7xX5IGW7v3z054YjbwGOapsqkqP
0u1q0wzxckZbCKYVExPQaMENU7fv6hvPDp05Sz5bB7OvkkvLQkKgOT819bjLsNV0
+Qpe8ELfUnSA4epcunEgQvED/Hw/UtVI8BaT2nqAwxInMeMK8Pvc7Y2YumCzySFp
dWrQYBKw3eKNMLQhsL8XahzF6kT4XJ5umbO0k3dXWHALdi55SO/ajCYQZexC2L+B
c8YcWYYAYSwq4dd+cbPMg8jI9gJRaruav+b8GMbTgnjaKr2l+dKpRkS5FE298mEP
5EGTJLcBfW9yqeTzucg31VDSdxwyS/0TWbCTWx8QG3SWR/w0HNuA6RmDYJ4mTnQ7
OJbMnk9Qs5pgLkAomd8ZBNv8ALozXwNjTl1hYhQKPzax953DGcKBtoZKAt5yHvgD
sJHJC1iPBUx56KAfWiiDd1no41+0uAfuasBNkI+WVBY+JkSlZf00ipiYK3JrwCcY
7Cm5TagvpVs6lWuNvhjkCjrFfdjs6IWKyDx5Gb29VL7U14lPvcRy404hYMf4XxmC
a8H86xquy6TUkYAI1lPuJtjXcMWBeGkH0kBMWYH/0VweoYxeX8RKUZ1e2LbQH9i8
+dOSPyeNfgGWQ84W6VspINyAXffkXVZpv2zoZtEp6PYb76Jn8ik3a84/YMVi53o6
XcJaRAFOt3X2HuXFid9QnAK+nqaTQeVPqMPj1SiIG9yJLI8DYJcCFSJYKYoO0B2c
EXeC6N5ABUP6vVA+IUWXE0DpLcpc/hxF5ojH1qNY8sx4CeNd3bx7FfpIQ/15HSSy
HiwxhxxfLOTWU57wr0mCNNxnKtDg/l7KhLuwi4jRJstWlVrSI00ZATGB81nWTG1i
pVu9k0cm7iEu/5eAyKjUQLGxCcfdbwJNoUJVeLG3v76BwurgY6xXJZbVa+zDncR7
VjDMyd6J8iKB6kjVHfqJQF9mqV6FebeUhZMqJH7GwP6MbY+YbZ2Ibvw9lAAgzXhJ
w5fH07MdY7v5oKbRBlyfGW8/eEmORkls4oc2LOslXMfL7ePneDRLsovgDDuB0R0E
+QM6vMw1HjhTr7vxEzvbPmgdtHgzWOJn4YgDDE+/RW0Fow9nm6qWZ2ugvXtF2kjs
mhia3pFqizWUt3V55EFGuXPN478avohC1S10Eow84KGTC2bHp4o+/w8mNQed/ium
6PVLMFZJB/3GoDi0eAT3BSnpB2uofxjdoxmK8TKFL2ILiIAdACSDh0hCImpcHAF4
slfdItgaaGntP01C6JW3dv6mrQtPRuIEVnWOSaFoQ0YClgg96auZ8/r1iPhHiYNf
gjein7yYOq38z09w7IudGWPD60YPKYuGWKDCFx39fXgnzXceXIPGs+DnMQnoUc8o
SgeEFL/F6FGrtp1TruWAX54p6BX4hy3THIUrkjdQBGs91KDTMGxBM5CM0dqhgjHs
bxEpiOF4fG+nVgvHKWS5zztOSSTlRe3/Wtdt2Se8D+hP94C0LSRhFj0cj0D8yiND
Sy4F6DHj/qdIU3LxzAJpSjqh1FfwQPNyLn2es3PkMK1V7AKiRifCdU55kzB+UGJT
FOqJ4pgkH1X28cFuU754sCG3Kzos9Sq00Xo/gzCPQW2b49eAl2Lzakr/aN8mSzj5
`protect end_protected