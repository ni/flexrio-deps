<<<<<<< HEAD:flexrio_deps/PkgDmaPortRecordFlattening.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNbi2tZhE34OOv0XWSzwbOVG3YmBn7B5kG23RxWuE0OJE
C30aB7fIj4cvggH+rJAL2UAXO5uYhP6f/6mFeLnnFa8HxqaHJCgTnFC5RUWkqfdq
0IzcjJXQdDwjmYtytH1qkJuZfIXB9SrOfAihSqCJNk6diQ2FLd9PFosXEZukzZYB
IyD33WEVYiLDrF9FNvItLkEYuQFj6CM8OETEvFSsPkdEXTVlwK9RfaWMepRrARXk
LJn1vUhM7fozONInOmyFnRaUnLYxxhj3jWxIyR7LZQiwoiHKPw/3mqNxre8IBVij
Whwu+iVAIKrHsRfgQEgFmKiaRiythyYOo3wQZWr4eLUgF8migB9fpqYrzRQVWx5E
PjD3Rss0tGwiIfvquspgXqAxaiMqHWo6IFImqycKAePDtfxNcEDylD+4NUsuZHq3
SUztfWjt43edKVMwkvMFx3knqR6HC+npceCP6ZZV2sCQI+m53FuUsiBQeODdFYAJ
1J8BX8/tFVOxeSvhaY6ii3/6LL3rv3gjLi1P5hQEwGsQ1Kcr9TKeQ3in/uT9+ciD
cM6duwGZQxTE4GtYfpe4sgUy6+jZ/WihLq7b7gYY1iuQSMh6GmaTv2UspihZp8Dg
HfvUgw6eb0gaSp7qLZtoMWhRCGV5ncBQb/3blhMbRhB4LFmQyc1fGa2WrP2+9sr1
l/iLrUf+pOi8saTUfvkW2r4R3P63J40aYJEpbNESx6xXTQhFg9mvHKfEH66+8dMa
27bZbeXNdcNeUVfH6jITaaizrM9yMuu6vFQOtQheCtWQAgjn+VpGQL7uUfxWRdDd
X0CI8faxj4jrhgvg5xluowCcfNBIp02i/ySSbW+VUiKBAaGSGjR3iafw83/VHelc
+SIbKJ3G3r/FVkWP8tnXdpU7CQyOGwftkeswlshmiQMJZbSqG7CqnbxOk11vr22N
1BLIFp6ArimtAxNpIEsYv/k5ffRdlaX8jqhWbG22QRd7Pl7j6ycCUyEi9tpaq9V7
oOPGd8YByLkRq6iTp/f2bnTs7gyIlWJ/68McT3y9OdgDuV9mUk6ZxCFNJiGNU101
9h127W1DrByZhQts4ruI6DLBDHZJu7J9bx5mw7FYttBDmy/NZJLxFhAMwn1gtQ0c
TXy79FfAfJmpbyNlJ4FqpTWX9yxbwDUQSBQ2LRwILn+h36dlxo7UZB3XQ2xO2iX3
LFDb6SQfm7KozqlFHlGqAr4fZBwTPY0x2JjfiI+5o7YWA/r48DEMy70Yo8bpkGAK
smU3qJoFDApCPYgVk11MAXi5cKrVz3Zkqriy63eRi7FxEXQZIc3y/DnfWg+HhfDO
kBMCBQUyUDAUEDpHPseAhcHAMoeaOZM9lvXwS8oGDhuA0KGcAnV7huYis/dKDNTu
4Fp+z5Z6KpypzQP2nDMWPY23JFCOg7o+qin2Su10MteKqXUkNoUZSnOWivwYt/Pb
Ai64pOWCCp8Zy8ff87dU14apsdekalYA1kIG5W4NFQMTdbvaD+lxFy33VzTlANDT
/Fs3mYnkCxMClZsHChqbCSjHRZ05tuVzqW+dJQELwBvIgrcBZowvYSHE9mhDqwCr
vZ9e4Fhd+TGklKgSd0vvtWhvdsYmwjhiYMwK1HToJyskCcgh22bRkjt0noTs26fh
ySqUfRRa3jAmtFcWxdTR5EuhcBwgJ/QtYJccQtPuzyF2r304a1a6g65JKvLqXSGL
idpDqFkblZTEcI9qWH/8sFlI1afQGe9ikO5d8cfcQb06Vg0EgM9eOV1LZMmXDdHE
uxqk9DdS0iVLgAtC+9dAVnO9tk+hDT2zBrpMzFJx1rCjsPmcdrkxREjQpoCmx2K1
417Ytf0kUe4QqO4VetFSnBrleX1ZrVbZeOzDs12l4HsfU8foD3oPy1S8LmyWIADz
uAClZbj51rRJo5pfr5tI3KiAtvKyumpVEbvqBjOwYCpKhAuGxxOn6+dZktsH7iFK
cr1P90S/6awh2XwbT6+Z4LfeQxtqEOPBY5aG8LwWCmM9RCRLcIrvTGHrV841FG/H
SVpAHvv1DDzWHNGowj5dchC4XsBMu9NLWgjCVhVNqVZsHwaUVvoWE8YXW6ZhMNam
sU3lBTZcphh3vPu9rkz10YEADF0/R28l9t3Xdtu28koHE3MO9CTE2rdnQ02YJFE1
J2I9u3f1AkihgRG++KhDuGvu6Q892rfMYdVZwtNorA2ukIkyxiDegalzyF989FmQ
mXPSUX1RqacJW00siapUjM7dVWdhcEdkQV91PhTuUMxr9VyT+orrSKdqbghDiR56
irayszz6hWlKB/9vXthwHMr/LYN/vs5zMaZnt56GMsnWGhMgG7urlTarHlhdEB+N
z5pJ7Vrxz7BCa4OejXoYLtmzbpfIZUMAGwKZ2c+mG47FrnE8k8egRip+3Ho1mIH7
kAvNjSfz5tF/xv47nHi7RfOdCZz5IDRxgHh9c1VygVXafaXWgA82wXyPyaEYzPvN
QpXGNyf+tXkcZDy/Ydv893qEulPmvAQTQLBHqJQv//+qsNRtlogAO6zgcbjVVDML
AVteYo92UcXbO/tI7DxvB2MNgnt/4gdMPBkjZgAFZcJcrs8IpHKT9Tr9Y3RR4xlx
mzKF6+gXS+wJ6eYCBApS474FuZJwSTZk+7GRgXP2ZidqZHjZ72uveMemOQGCn6nI
AfTxpLngjSv5m6CPXRPnIaqLwvFMbnpVgnHp8POqZYVM13AlWOqUH58qtSpaltG6
9a9EPK9urRcBBq/6lcuh3ovpb6PFiWZWLP+ejWLn52i3/93ERb8JjHIDZzXU/U0Q
2wMKbNTecYVnu3XgfuxFtteF6EChaHoHK8jk+vYpM7sjpsuT+i47p0OGkMDfc5n+
9CH0BTrb6+jxiYeH4e4s+9zgeB3ItkLvzHv4mLa914mhF2CJJsXprNC9UsdN20Q/
QWIXd9zAlYjuIk5kAKVuWzV8aTf0LuXWSSVjkxeq/yZlWb4pzRbtp2/54mxE79Ys
p5zbCtFVouFLqHDvdgoK0JaXtTHIvrENotwFm2shkIk8k8exsJZqdloqTwyKmGGE
VSAgoJDERKirSzWsel00TpjfYJIFMyls+Fy2r6G8kg/ya3qxgeufRzRlJjUM8kxq
nrGDgxMGFkFKgeYzOnv7mS4B3p7rmmHQA1UZQenKyC9hPtoXv+Hk4NoNV1PW44a7
/ZU7eVkFnAydV1c2UhPapV+JUXD7yVHq5iw0p0Mt8WG1Gld0OgcGbheLU2KSCnvh
GdZ0OCwDFIV4fjolo6MLiNFShNAOH2Ob8Cr+EGFGcQAD6hcn/H4QKFO/RV1I0Ydh
rP5ikL6GVFsNJmks0vn/F8JgDLEF+trE0DDl8I9BnQc8gGj3kAzrFi20qiNJcEWu
2+xQTm8YCx4/21pUEoDC2EsEbbGYlNL+UBsQWsllep82nMQFiRjLzejHlDqw88T9
3Vd0GWKsgnJezHC4YuDwB8/eQJbOgZxhl65GGixz3aH4r9JA9ImZmh03Z8oBJbCG
BNCx+TFskrk4Vr+7ssx1Be29Yati3z8gyuCoGGuHNkSdeTNz6wRBbfYuE//d2jre
QqDHv07mDpB4/WQVgwJq4dnxwM2OnBhvHxbT7G1UtfWt82HsMgVAB4W2CoEctWx8
r6jlGYTHw5yLQNoP4dTrXN7CZFmsDcRWvpzxZdAxBBKOlBoLYeEdFpQcHGhb9F7U
PC/Hvn1V17NMQxmu67US4igtgd2/Ujct9Ba2tWOXoqM+h6yC2P6hBIaNz1gago9H
lL40zb3epnDS/1oEePaOp/1H3TT88lybFhqyE2hjSK0EcNiLZ2KyJqKz3Ntx9r+z
PodBPKtL9nCNITHmpfA+DeymlhV7IYuGB/3j/gz3vTmJAwDi2uVWGC9/XxY99Nsr
OkaWTvFKxwRpSY7MOVQUqn3HIPUhe2vj49uK1T1CBakNJpkgTpIs0THh0jaSq40U
NjBE1Dpt1YNYJjelkKO54Evf1Nu4i0aFFBXBiFBrZsZwgsDt+0fRbBDI5Oc2hHkh
GzUK+VCiso5XEwhiiD3fwWOVsvcNTVjmQmfsMnHh8bbN4jK0C5uArIjeaPwbMip2
fP3WaLl+AAo6ijlEtvM/TlGMeIe9VSadSEEsTUE+OvzBj4EjJ/rLXvbHRe2LGg+C
kSfa+Co0aKLHmEaGOeYSJkEF+D51rQ8zMhaa3FYEGBwRHEOhu+g2ndyHGkErxyDH
txCGoQtoJVlXVcUrUqprXWlTsqbFearW4Lzs+Hq4O7KmLY2evw1r6hRiTuMNO2Vo
z0KS86z6LS+d+TRG3Gk7rGDxSKIpP9oXOqrwR+bWHWW/ZpRo+z+WjlyQ2WL8ijsZ
IIDUmZNUxlT1sOS0vCDadPIJo0T23FuvuBjf5X/8B+oi0lL27gxhgssULgKTmsGP
648fQU4I6us0HV+hw7PVBt2Pa7/T7Za1trHTD4D1KWbqASgCdMaGdr9woSY+TqvP
t68d0xpRe+xt23zQAvadpB3myGfRlLuj9Dht/Zu8j/c8W9gi+20tpqT6FFe/tiYC
GlUrI11LJwm5eSKTKJ4zftr4s3ASmXplEUp5fGJERoxDgvccyX93/E4cgsfRIR6A
GH9ZO7exC2cMaliJL2lVTuANLM2IiyLiGoIjWdxdbKJw0QmqAyPJHmgnU5GOQAC3
oq3jaojIXu0cnT+CIRKUaJzOjLhwaKXzGXFJs8GLI1KbwbmfcG+8uIVIMSBViBmv
V50+45qooy2kxVDzORKUUQdqGnY6Idwp37qRHfDENzC9ZItNFv8xAZdgrR9PfPel
eROrhNXxJP8b8yqzFtLe41sU9e6GW3pwYTQTIMBLUkQ/JuH0GcVxuU1upOTym/vI
gab5tcbpkcGdExMsjehZwYvYJsjWtiRg444K3GU72D3ZDmjK8XtE89rOUR9HFkYk
ObpYwEkBINv5H7g5YQc4qkNeOn5lPLpU4gP6fJTErg9z6xRnrb1hMgrQXeQQOtNi
xWZVHltq1E9wqtTE6Br/NVkhDvbW8A0XDth4qZddPT9e8NVPC44eG4AX7V6vRQHW
jqg5h+FkPbf3Yit5QgC9AwqI/abTvEz6D9G8iMITDt3vkCWziUusaa8XySJrNwLK
2qOPgP7ww4yKjYApQsR84XZdJ+y9+CPr1nUMnMjux6Ley+aCGqiGyJvJjZ1Z6dzd
5cr6d9HDeeuGNWErLB6YjwGZzYrLx4UEL65dT7pMNX+3PpNrTvrDBhyXrqLpfzpy
8yp8YSbu6FKF12PCjPFQrB1Lc0yv5T60dvBAwHUSAR1km9JQWO3ocvmiKTSyA8lP
MfaQp2sGshYyc2zDhOJcBnqcRW8TDwhYX+Iw0PotYxYDfDGWuqOBeQ+0s7WUp38c
j89xljlKaRcVmpxW+zwTM4MGBSkoQEJjGueR3AyrMs1vRiaR+eq7j7YE+3jom1lA
gEYbR8cYmw2RCc1e/mkA4ZJUWOTw/SY2tyVUnQKjZ17bIINJCluLBSt2lZmnoRwF
atmF1c56KHN0UoiOt64IU7BxNDiQ/90V6GmtzRTnt/fuJgOGfo5CSwsShheg4Yv7
RP3kq3JQJfenAkQgJuBNOY4J3IBMDZ0cv5v9M2Q9wNkFiumLcIpqzDj2G5ryqy3B
58xTk6sgK8O2HcWVyyxGeDPs5lb26uitri1VMSJGabgy+1jEGxD8n9n/rp4Vn8MR
B99kar535J6iX5u+Yc5C3N4qx1V6bKrkkmVq/GWlik6g76sykbuQXAChLSkZqCHw
Cr7DE1hiy6DXWMVH9BcBcyw2pK07BF+9GVVHHgbbAk6+1QgZlgu/sAqen+9u4nkv
gUWYcCU20UXQgXBKaW+VvG8dAUlRbEqjJPs5OXhAAOJyN6d+5e7gCUPBbuxTWCTG
JPQuSmA5vHZz5Y3fQMPnox+DHMc9jacViT5jND3WsKNCYCmQ7cisy0UjsH+uuPOo
M9b672T0hSwaRjLoBox7ZlpTCxV+nL6k9kTd5FQ1XTi1CYKMPnSSFn65lJvxU0a/
b1bYoetXKaKpxbgBASWKvQxPzKJXuaYL6UEtaWST3xRogwfO7Dc8YZqhf7O7DX4v
gvR0CAXOvxlzlHvByldpREdgryKDl3uGL0WNYLHSGukWHEgl6XWdIt6BdvbYL/pA
eSqc6lPZWW6aNV+Oh6CGcvxFmAsVMIs38tFWTTskjQ1BN85S9mzsNlnDuuI86MLD
GuAfg7SmTE1JXfd9V8YFeIiTBgYtN24V++nGWoxcPzoDuW0gUADpAjJexHxeL/DU
FOdZH7W5SC/99iW41Lf7xgNUZGKVcu8/iui5K8pN7f5Evvfd2XMBZr+fY1edS/qb
wIieI3rxAqkBJjNSqXb7RzvfCuOjIEfPuKGczntzntiU1FAmyYL70mGTzqahYN+8
Zf8TiB+yS1cE5BVp4MVGqo74G0xyCezdQE69GVXy+Onou1ZS+kUACC/VzGW9v608
ffqcDS2ormb1nUnFb1QiMrBTKCFQJYEptwqaxJMdD8MqmpowsZlSbDXc25FR8uTv
RiJO3rQCSXN+TbLTmZaMEbZOAsKJzzC2kmPJlej776CV8WBLfC8x7hIyxBAWMK4W
sjoB+y/Mrvs5jWvGLovQZcyTAn/Yji9Go3QUvN2GNZvNurBGdTgb0rHgwghEzs1b
TIscrIx59H+SDsh/r6fJp+aAdqGA5EoJqtzhzkJSmNKvAGQfm2rlX8WQhYvxMBsz
eDtNlJkv9i/KQL7PJsSne41mqdjY1DHFS5UZWmdeqFVNQ6zufT2bLHYetIARyBD0
Oaif3zSxXJfYv+XlKEBj8lexJSMDJD2YA1rSazXl3Pgtg5O2eEMA/cVmVAulKLpy
5/kQWVDMsLO7hSTzlR4hAaAC+0/1FX1V8TTwMBFsW6H074Glg+Z1SOUhvnjR3EKW
VJYzMC4gIQRff70dLJx3Xbbo1i0oF4E9qfWM+GNtZASEgXIlLq0jY47hY51vCvDC
zt8rDX4Wyn4wCZyAIPkQs6CzCIHGeRlIfx9joqfkm6YJOB+rS+XATYb9ZYwIgAa4
WO7g2OUwH28EaNS40HcVGac6gF6Q53Opr2jHyGDq0pf4SmrXtP20bBlpqPJXT9FB
oDHf4+QETnm7OkuOpjRj5Z5oixfFecGLqL0XUQX/fvB5amY9TN4OErSvE2PFwkne
YCwohp/8WxuLfU97YaB8jChuOuH1PonFPcR8vR/6S7hG+LrvPXfUw2lWQ0M9IjIL
6iW/Ub5n4bDamRlGaDVaL/FjlOdl04FdTyhAktQHjpQqEN7VmUJlITSh8GC2/OTA
mTmVfyvFYd3FsaCzjokECQWnjmr6UMkSwXZBXRioIwGmUHIgdT/AEnsIU7ul0sjL
VrntWKTpVxsvNSE8krLDgD1dfvbe8NZOi0pRU35WivRMe/kKc6/LZS3fyrAzdYEb
gqC0Na1PHs3iR3A5cJJg02bto5pnomND/tQZlvBC75A1pASbR7iAywDJ6XrqPEZf
kz6akKCNydbTGQmCc9OkKW7mIwYgIy+znY/U27tMEoQ5H4hFH6gebbaq6VyZVK9V
th68KjNHGJZc+xdJeyGKnN6/13n3QGBNIEQCMFtceBwgIVviA3uG5NoTvarYj+p+
135cBxTRX1H4E0NNcbmynFTXvP48n64AXhin2JVzh/GNh7Wy2Gw9aG1L0QVqDDNN
8bSI41BMibhlPhh0U+dulbX4A6rfVD87Gtgqw83mybBOWu9hFXUP0FRqTZ7vHPU4
judEaTI13HaZvX8LyUt7wMaIDqHy3fzhqKeesYeZ8tI4My17M+fJWkguFiYRqK21
9xrxgx7Zew6wopuoS1m2xRFI7LciCnsow9QMtvcvtKLQKd19URbwTQFVo+sOnOyP
Ad2qC2oqAiBpkfOjqjSH0iWH0wyyCx7CwpKN7fpTyVVI95aAEOJXosOk5nov/VnH
AGMHtVP9WHUkAxBb3OItcehw2FOTch+TyWPugRJ+241RdainFp5GR5PCluE0wECE
kDC1Y23tBLKDXugpXfC0ZU29yI7ZuuEICL1WiimlZ7Av3q6w1AbwVXJd3vDtiGIP
AgUT8VFa7RniD4eDoII9KilAc3M26q9V/iBHxWWMsnR3O1kqUtakckZe/TcMlbnN
0xl5LTen/u47IuaBPirHApgkffxLXLh/yHOnCsu5QvA2nacCGL0VFGJ8otDdPOLT
tGsmDzRATce17FZTnSOZIllLFCgNko6nZ+tZD4x9g8+iqQtJYmwoUJW3WQPkgGjP
h14ToZ6XN2v/CM6WOZqi0Nldy3T8L2lXHduGIMFYA6xkDQfwPy96usvbUJZunQad
QvYtXMMXzlcS0OWaypsCjMPN+lT1n1YrTKOFaYo7cQ9T81LRRk54wyW3HH797cZ+
EWI/B3GG6pZg0srt1++4qujcG9TWT2ECTdkSRh0ZWxgbXOE3RbhvejQtolkvwcvP
D9ESRsxbJWu1GChB4Vl8HRZGEAmZirovYkwJeO191Kf2xBYU/uIZpTo6fsC9HPQa
aVWI4NBPglORtfkEVRCiSTIBKvLZv1Kz8UHPc8ahZfxaC+zPP4sXG5TSBbM0wvMJ
EtjoSMeIMlax1HGlTJN7/H9xNEQ5h5xXQvUnOdwDxSvAwgzI/q/tcbTDGTu053IO
rPqRc5eV0ssbaghzD0t1U9J90emRqEryeAKL9+wDuGXVjecbD01yQBrWjsd50SqC
M+scTLscR0g3eoqrXFYHfJKWnJQ5aHfETx6duQY8U2QqLgGD/z7Ke0UfuXENAkGV
Tn3NnskwgiesIiMghaT4FgbkiJByhIQMPJiMe9gBmTphVDXGZtJi0adGOLS/ZcwS
iEw79ajKvHiaE3XJu9ShuuhSj9T2boDZppvGOBs0ptPy7s2Ro5cjjsGn86Ucci0A
yR1e6xZXpmTJrql1irgOoxB9lW2DfAQFd4+jpgjPDbsFn1efY5ZvTthxMMRjUMD8
GDLiAubaWt36H56MDUMyWmgbBPoLIUVvE2kUaXP3gN3T3qsPS+spEZZNyFRfg4FZ
V5Lsqt1BO+mY/07yksAjdYG401Axns7rrhDQNYJ0HTOMNNd9BRZVrHyAKdd+4CQf
hEsKc4yz3aWLd0XrQ4v1UREq/Wxl90FzDILhRUUPBkD95vn9o9DMxjzkbGXG2cP9
PumKbT5WzsXP+NNe5SDcoHPLoGfq0A/VUg82g5NROaR1z+f7lDsrGuhvxFF+gBum
ZR4xRlquyH30b85cI65uMLPVah5Cd7jMwgL1j7wtTFgXTVxdGTZQNRHVd1eNH8X7
iE6BI4o53WuZ0ykgrapZ+hYF9/Xet10ohHoSgdxw43ZmbunjPYQxtzb51T6x5OfQ
tKo3LGSqrfO8ETiyRXFGiBavxsXcbwVS4bPLWzsd5cQkXgIK4iQMu0r3Q3qBpM+S
4KF4oRAh+A/PPbo7J19b5bGzZKgfRBQg2Mc5oeW9jvimAIykpBS1zJ7akUvPx4l4
qmkZu7/4l6MsdUYjJedUQHnaNiVvw1l87PnrCAnNFLO3h7QimAcFyy6IHaRKrAu2
HD+0y1vGMYqezat0nvuMbQyy8vpM83UpyIIUZBy760WsRT2Cf9MXon30AH33lNix
4y/Q6DFYDB188QPF9gRpj5vp/fZjZ9ySIUWn39RqflubPdvWXnDJRzx8YLOVQZZF
uVLaqihd+Cc/jOkNSlX2IIqXxg6VL900FJvqmSYHfetb4uFWXc+nRS3IyrH6eNXm
fyuAso9Tm3kY/QabAsbllaya2BGMXdFz2wQxW/BSpt9A20wkWHaQika4MoAghvmS
p//mDsimPDG/zmDH5tMItSOT4rPuRdfypHKSCoM41vX9OYFprdu2+zKnVuOXaVJF
FPI4+qZpKLsRgXI+QaopOyyT3crPpnXNlh9TJD5hfRzwa4mm7A4DY9bvjEZipp0p
RKF9Nhd0Gnte0uVlE1i3LuNlji+M+CS6JCnCpP7WoDydoLb3dBc653bdQP1BkN0M
HILXy+I+ro2SWys2cwyBmFXUhdVq9MQS5Dv8KWVOir0omJgebknRvU4/w4WG2B8x
1O8McjWVm7lY/L1SayeL2kKquV9inBd9fRW0otWGt4qQrJs0/Vck/7qOuWc62CHS
K+/snWZefmkMMr+XKsaYRPY++1HEwq/eK1+knca47RR95eCjKSSV1eqpcXEmdL6M
iuR0zvQdqKYvhl00BBL2N+TlkW8bXFab7h9MGvGBMqfZAKNXh7HcWLYaGqKQMJ/k
GalhsKCJ9/ebTll5IqhIq7svdjkKgUney62UIBPW0GA4kNcxY/RLYBCUhBse/Lbk
UWnamPjAMVV4ZdCxOgOEhbRzBOzgufJa8+xrNCL2R6D0KtxrY+IdZ133qwS9oiDx
tAE/5d5gDQX3O/UuIGzr7/qsU/XJ3deXPcP02Uq046TMjpNgWa6iiOXN1iSZszbl
XEXM7xqoVQ8ACyFtq6BTGrMTWl9TsKgYaP/vLR5fNTJ8N6Ek2Yc+rog4XFOBLWHu
E+HAqw01qOwwXWaK9lEJuPUnlwYymEpT1LY9BJXM3rZsgmQAHycyZnvD6eMyFtVc
ge/od2ms5r/F2REgbJAHnhQe0OIO/zV5GP8h6EZx9xPeSxn5nP/Batn170r24XzK
1iIMFmRfEaunadaXuVZi1Hsqc4jL1eNH9gx19AKLvcu7CxZa73cWf0kGDxyOHWUw
vBBd2k/K8hJ34LHBPW+AQeMo5Dysf+5yoEbipqy/8CCJw8/UwiSKJ8ASOhIe5k3F
Hxg+d8C648csoU/drdcAnOnamlzxqee8ADrNFvWpcO844NP36IlfE5lyQGfQ1GwK
nSwKJ8sd+cxHPy0a/ZVsPq74fdCOIo/qUtKFuNn5V7VserDwgzRpwfi6gayN+eYL
JTUSLRaf4uafiqb+eG7q0umttb53hxP/C+H79aksVQTExNGHPfNkL/pmlzGr43iC
Ag7Bc6Fj4jTE7S6Z8yGEOKazBB3/KmK2pJCtzSQMx85KPO5LJ5q7MXqAholYxOeh
aBb0UjIGGUyUh/Ajar5smUF29e7tR80GZ8H2FCzNL2efb0pA4Ri13vIGojfW55Pq
p7TDUygq5UXPbzwwkRAepTTfCHK7h0Coa7+68BTCc0XqBNCzM8iNnF8Le0AxycLp
Am4EXNGt7lu1EqOrX9yx2/HaUCT8NLHF5WLynkR+WGljWCTzv62380z1OQWyR7Mr
2tXcGIOIcDJeOiGy617s2SQ9OfqFe0SFPBQgJYMrbQJzs1WvWds3OVYP7TqWdYbE
g+Km5zHik4qrI/GIksWbMfnC45aYc6XvQcnwPsYO1M4S1dy6raTdC2ndwCIAMTdm
ROX2uQB4SUfksJU2A2nRXloe+zAwMjJPTXL4enwpc7d4mn3qEE8Onn4Qaclt46Wv
AF/7xXeZbPETi3xKxo53TmRPFTgUk/sjqPLk0zb0XjuDGwissnNmGfjQCGRnB2jH
YlLBpVyeR4acYItpU0dCmxNxKL6FaknqDelRo7tamtL/5eZduFcDsIKdjoXpdcCY
FFJo3WtvnsI018AwfzKV9zkJ9ysvXwVpef+IeKDOI8UF5XawvPIFzcTsyCcXujF4
wH20bHWrY4lgG7GWgCCjFICbIAf3npeaNth7RkFtIWdQf6Dnya8n8sbwFtjt8LAU
eaAFxF8oJcGGr+v9/sSMTGmGm+UU85uff2mUOVZbDxltAqRhV9jn6J1WyqX5MSwu
f6uW24BhlAnI21b3+jBJtyQurR7YGtjtmgBK4oLPDG2kuOaErg+a8S6dP72cZzWQ
K56laXFzrZZtonXkVj89KeZs893ao/tlF2NqzQm9Vs22PF1OhovtFgf+ow6pJ7jg
lUj3Wd6q+ceMjEF45D//J80F9HpZJy/1B5d2a+RQeADZj5iTroAI4ZcHbT4syEQa
H2rPO7trODD+vRThA+Boy0CDPVDu4tH3IpLpVmkUg+fmiunYvlovzbo7I/HPOsGO
tJ8mexJh5INbEasqnIFYXVpKsjFB0FYfM5xtECBWCvYKDs4i04rwMiUIaKyDAEEj
HstvrdhUkbv2XzHPRmjQ3Kl2k3g1lekhSRSJ7fZdU4CwJYy7WZJKCAU8eYTVQy34
lqey2hAmMeVlAf0vcERrE56fiDPyQGZ2iT7EnpA7xvQJgUXZuFh8mR3Kz9ZClzJI
bjCV60ufMxoqwGK7duuQ2TTxGu2keGzafHxcLL9lCc8DqB13gqPz9Ce7Z60NDHCV
0NLbwGbR7ud05U0T9OeMeC/KsTYWHzWn/EQHZy41IrjBs7ETcx16+PMP3B8S3mG/
jxeH10quOg1ihH33m3wd/Dmj1jJnCaOVCV24kSYhTbK89aOq9W9iV4usoZy9ji+t
5G0VRZENZitM6qP5AKEKFPVAy/13v6tz2FdcBKQHq2QXHcN1SO6fJtFVlvCntn7s
kDFTlXs1wqlVK+0men0Y5aj3+NzzTM72W6UUGielgLsPBqB40rw9ZhJNkpvtIQIV
UIhX92COoBBaNstwceD17z0mtKUs8RM63RfASxJBQf/KKzpxNVrUaAyLu8cX9v6o
fQEIQDslJUhf7HNorAc23mAOr9RaRWd7Q5KbKZ8Gjxk2bvIiK9fnFJ6xISIkYPk5
NaCCOuJmcGMsbXHIKWgeQvXbDo7ULuP83pGRWnuxK7s4utSIRobchO3KE4bS+Uuj
4VXkqvxgKTKZazkvBB8NfKwkwuoG+hnB7O/LjFn2yUfHuwloabZWjeJrKp6klekl
PXT4ZApuu8UkhYkU4bM/GQ8T4iwEWSEmNhHwzvQ4urtrsKCDuCdGKXcX/vLZTgts
Zk6/2wRmjnoPMLcb3chzSaV1DN2fC7WNhV6dgCKZh42x90OV5sCpt7jYTmdAg/VO
/+R078rWUlUgzbk33O5tM/YF6MRuqJMeHa8OZJttA2QHmQ74v8ajlMXfeeUqUelX
We8Xnod/08MLTeMjztTe9HtmByZ1t9DZ76HuTbf4nSe+AN0Iusz2g5oxMbeZ6lr4
Qo7EysWWjcCSIUUSm5NsGzPXQ0NoOULh+IIH/oeqK5f9OO4wrh61rtWTIoYcIqNe
P32IXf5a4SNHDNTcoMSRxH43syAJw5gwK8y7S7CBsmvhQxiYXVuyeCSCRMSdjv//
F+jpttzYWNNPFWuLogxkz890QuTLpURsDrFAgmsGpI0I085R1GjkdV1MkNBC0Zye
OPAyzuwY6Qkb/qMCnRGdNjoJcUWyrNeWg9c1ezgDPBoLXxBeYor6nDV6xPazO+yP
cKDzJzAog4Flno41ADK8lVMkll7drmllRN8DByL1KgTJmi2NRuoMtOAV0dUkHaob
ivMc7XZqWfKMwANkB6kuvvr5nR8/KTPcS8XWNTTN9OP2N9Yi6BNgFwDU60pX7PDY
wN83EACZjTu9n95j6UPJWrh99RyKdNkxUi6PiA7nfOXNpCUV15jwhr/R1T48eziP
LuR9NFbgXVAZ7JO+47atnGk4kiXeszYEh2dnRaLi353tcEOl/r4b7oiUpivZWzmo
0ctqfP5SJ2wXfj7OuOMue4CwVpRVzLPdb15eHI6+RvCYETmdVh/gyzjHGT0oJUvn
pEjedpmSYrtY7ESmbNuxUo6tFknz+KdeqbD+a4V66OugNp4pbx5q5fo16gms64wH
t4kiYT3LtZmMjpTsaSbcXKh32pNvn2dZH+fGX6KZjqHRdWHTUx9k+0cc53RxAatC
DOknp9EzdGIlQwbcgSh5rMRk+XPnjswvvC6o0h8iVb3FzMnOzCceEtV4Ao++jtL7
cia6pAMecimor3OFXxDVgs6kgs0BNZC37oyHctl0EfZGFPM7lTSMRTpHTICfCqTw
r//2m7YRTM+CC+KZtnPDcqoaU8Ku22wC8gN+Eusyq6Aws1hcAAdvFCA+IxkTYcV/
dsIXtD3z0VrAsELLbo5hOzAOFLO6sBEiUK+0uMbU6zxRxz3kxxnpsZ4wZxHZ5+V/
io68FmvCQeGPsHq22VqWYkbbjtM5DDp1DAlZs3/o7djek1Tgpl17sfODDZD6vp68
17wKBe00Kb7rE+nCiSMlJTghYCCtRnPnkF9tfYfUYtTPx2LnLUZxHOrJEuwWe4Dg
dnaJbYE7wFfZYPgbIMwlNgrZapCDdcItp8oAg/UzgcodTOEkezHaLwVg1FyjBT1J
dL2zhMqhbvJ5riw2AWQJUAIWrNysgIBPrtPrxaj2+IMHye8LhE9c5XRsMg3fCVcH
vXoNFGCW5kKZWIDDDMRZMLOFlIxxOTRf8wzyD7w7XN+k1wHjlPk1Kz40qrAhItWi
VxZVRmR2oB5aXqa+wzYl26/+sRDcEnsskZHuicL0XqTlQqGzw7MseFqbHbipi5CR
zXsWAE1UGCZLsSwjz8wVhiDMyZHLGDF4WsxjSNa8NvP8ZLV6plIpAi+9kF59F4oB
2n2B9Ze5vftayfKkWwYrF7u+ITNmMdJYvZj8CY3KQHgK6QSFDVk70tKvIM9rfdkS
SKCl8ijeqoCbTs79uH/v2/PlFJOLCc4AjYwMZWGMRo4EPnnA9lMvuiV1BHlTwnrL
+QgE0NJuRVAZpRfYQl9AQ77DRpmU7w/wEUtZB9LFI8EEZTUMdyax7hsixckH8ONv
SWplFrsHF2YvBXyv56vgpouqoZQ/lNmSBwInlMQ8JNsl1JXllMoQf9nNDSIMIgU0
pIJOS+AGJ4fm2iBtqUd6AZ3hBxVsK8wmVWMqRL9eCBkhDwhTmE236yTuXXY11Ajb
ia/BuN+wQ1/g0ODe6MADfE6WGEhLQX4lY5YmVDLjyQUy77GJ+EcsNZdMZtfh+TlG
wIAJrPxRONxMDT2wEwyUeV1/lPrQ9mCYYO4ci3s1HXs4i548EgOKKHnPQQPqqEjH
idiFV21BeeDd5uZLyRbxRL3oKlxhqfEIX2ZqSQcF2ZtVJAOWH2JHup1ES7W6YsjK
fpZYW5IyebKO0rA80MsEFcTv0YMsaEsH9w+D4G0sn5J7NpvOCB89AoKYmajetgLB
JeXwZlfde/U8wHlhkAfQP2ZT36Dq9kFQ/Ds+uOuIRadSD/Dkb5iP5+0CZVJRb7Pb
neV8+cs5N9zm8v4LpyO2bwmRGnBx+Dzydx6fy7ItsrkfFHC2yQTzDOnkv6XRL7Qh
gy1iBLurlt8R+slgQhVv7UbDizs1xD9jQzIlkRTHHVkxnar1bqgoX2iWjdCSOO9D
0lTQxeFthG9AniQmfOkiB16DwnyfclyKcI/lD7nRRN7hHsJrlPVGMZaWN/zM+/Nj
OYcNxY1mlEo6E4OJYejkXhgEhrCLmJaTNFj4nlFwV9o8xs5ZNnx/+Q6LgbYCf7dt
axibDys8kMvpPEbPuoNfI5MddFtSqiK/9oweJiSmKmAC1hARYMZjorhzYxMkzxoC
3+IEMbRUOHQs2BxxhbTv+WcQPQRRXOjCc/JyelmJb9dbTiFWLTsCmZSlT1/C5Ogp
9U3l5MJ/a2QY7KtIMLwHtgIkPfPh17Zk6Qci/0vIGys80ap5LqM/hkMb6T51MYA/
aPwwNFrpkXFQHNECMR+D08nAhUs/1TCwUcjRGqWGxItraTrGRxNok+pX0RmdcWaN
4fU7x/j01x0fiiTYrU6ehYvZWO3M9nYB17vZY6uTxw29ChKuq4LAqs9i37bH7JFV
9lD7YWV1d9BaaeIhK5cxI/1H4oqGQX48w4oLvNnn8VJQEfaSy/tHqWXFChxvagHQ
7aq8IDtdwFuX89AH+xvv0hnsb8XtfGUbxH9IhLrCzxWmWb0yZWcqNDDujFOLG5W9
MdXY6k9W6zB1JdXSLOb1LYCWyYNVWiIHbYIv/bvDg71wfYzg3bT00p0UISJuK23l
m5xqAMq8Wj7EB0UqcgHo+1nSF+dsFHjZfGPqN+od7gDD/Yfxn6B+AkA+gjij7xd5
mwIFWSvZfAKvJ4u9QOYex6gjjwtRYw8JCy2geI3kedX9inQENu2cuW7ezyy3Wvj/
m5k5c4pfIKbrW3alibr21Wm2laEeVjC6bFQchswa7sb7kU4E39B/+AdruThOXoyc
sbGTGpSM3RK4UasY4Pq9soaUra6D6sxI+BfJmD2GAG2dkYFujz+ajAfaxq0bIzo9
jLnXah/ZoVxLhMJ3PO7+aDbuYZJXOYH5wzsHZh5soguHY8XMy5en7O2PcVLsyLFx
OnwduxUObVj1os+msTAqhHIBxW5nxk4z0TLTIqbd8ceQr/lQkI1nCqG1dQTI4v+e
ekpRr8pL1jpL+ae3N60mTDWrzc7JgbSRx3YzYDYbBOw1YkFc0vTnaAH/9axpg3LT
1fNABOk+8FwkB7HcUkM3xGCGozoupnPvIHRC79/nLEgAGVov+wvgZZF35sMBNDG5
c/mRPQrKJqFMiUEqDkCp573d4Mzla0/TRFFcp12Hv67XzKG1bnPNG9iFSJPo75vs
h137XOVRVIkhfAhh0r73WfyyJb2LoID/A9WksF4KSailw/i3lzM46uxXfC+Gz3/v
E2RhKMYIEzeBAmBzGRjYlrIpaaDxQqfqzT8toULjIlDbMJM7VWr4SMZGVQhVIvdq
ZxHO50N6bdhnBEc3hbmbcjHbYQrTdvo4XkiwVyUVyzx9ZaXirptTSzwbW4yzS8zB
HGoVvaBr8VjuDjkzyR/uDnQGlusQwNh44HJMMVRD7z0Tl49V5aEK70yeuBUg0WXt
o0FA0XzxyNhR8i6bHcxyUkC2lNXtaC2P6ecyvRNx+mHCbAwNBFXHnOzvTPVJ8udn
a5PmOBJjNlYmgww/HTys/NVPoOiPMRSycdWjryJLoVQhXIm0a0MXrmzWMuOy1vB1
gdOOkcsQ0IWGTB0hukIaPOA5hPhVGcy5heSAP8KdELWp0Gt1sb/MOHfx/1BGll+C
TpaGyp3FX1JsoT+U3lGjhV/wNyq39lEiYS283sFs9AqWw2tv4/HclIiQlDpYDMVl
f6DQfRu1b/ypnRS5LMhoNviCLwDBGyPk8ixAvY39v0u7cIS/yoPEnowKyYt4uLP6
csE1ASRgcL9RO2WIeQNwkN7uL3dNEjlm8kSHtT9Bur8Mda96l+1fk6kgR1LKymNo
gzncFzKqrD8SKPCADofsME+fAPtCGA/ZxY4jxBFxZfBD/OZ8AzrZ9nbG1r1fvL20
kaySTXACVvby/O5pskMMxm3gnNu8/hpM1Sqyh/9JBfk1IShvQ7X3UzQtZtv4sAuH
w/Z6SyN6RF8/1eQAncvOjZIOn83lQcLqHfEjdDpVxuAELxAOs7FMRDgpFAHy+Lqh
lCACJbyyadTXrvtQ17aCkTY2154RdV28rS+QDCPMJkTvIcNV5TbH5xjg2AoTFJz8
kXpbq045R7pnJmZnyuSMvVWkOyDx4VH2/o1xPrZ1BAHmkv0Ilrbc/3AvL9/JZ2R1
GhS60nyUa6D2aiGO6EUTYTyBJsl+Gb4Hki7YEDKiqj9qJeb0XwEVmSNxjzut7Pzh
b2WTOgf1ehK38cyuluxOK0Wnek8lq0Zc4Ie9YvSTiKRVD3uMLga8hjIHnCIEPI0q
DMZR/D8ga58nTH+BuMqoNu/hftcm+SAI0YjBCI4xdLKpMbjPmXu+WPxlvP05mVDO
wn6qeI9pd0ADHkvCaLkOfS1bYKSuh8BQhmzblmhoiSfufA8RIl2Jz9/Fb/867pTh
bT2KQPNSq49wH1bwUj/guBDhvdXQGvBa1AdUNeLDareb8fDgkcIYcEwCEeM583H8
pN9TQ5dPiKBj5YEPXIhKUbF0YbL2ejd8w4exy+QGbmy/dyDn33zHB+SAauk9x/9V
XYetnJUgd0rvsmwVEbpwXipkbtanXKMRD6ba+/Tnvf1UMcmy0B6LBc5IjfIjzTuD
2dlpRnxAdmjbLmbOHa+kLd5rfY0Wsi6vHDDXQSQeECYiSLk08GjfrI+VptIsyV5n
Miy8CTKTbrUxM1GX86SYzm6jF65cfUPXfGUXmQw+5rp140cu6baRr+TwVuWFo+IF
qHKtJE/0oyg1xZqNE8AjuS32sy7p5AH3heY6BqYA6v5rUK576A/asJhExO3YHidq
BGcTpouH1Sk+Cj+OxT8MLDuRDMARRVmJs2NdtKflhXBdi7X/ONZkXCJdYudTj76M
dW6ONcZmaxshazKCgEqWOvDf476h/JMQgbkjoQS36e3/yFZqapho0N7FwZ+ZqWJY
zVoKZ+2Dukt61ifVJ/kXXWB/tIWrSZjlJ61cwsj+G6SDG4g21hr4f+osjUJfZVTn
nS8cXyTqepr2m0KrKZmxpx4h3xsuyajLIDgo5ixZmqsS5M6l25gnT6qJkk0NSi6p
v/Ws0IR+Ya5wceVT3ATaUxADc/DAdrb6micmUlM0NmuWzYALF/Bmox7Bv4uie0pz
Zdu1CmQ0GzVZm54YNU+oafJOHuU1l/3nyhEkevpQZsGjkSc3TeSyKdxgu1mTcNsi
Qgv69muclqwKDfwWgmODqExtXxJBwHJOmYR3+uqEWauxwEdHHgVrjPlSenxeRzz7
5LNckOgH9aSMhIWoK+gISLkx2DqrzV4XHc6h8ZfEQx5VE5n1x7PaoMRzNUtYQ3uL
VVyk5HCC1PYqTDY3rltC4FLoW2VDBb+jjK8IadVmhSdpKCEz0R5nvRtqtObDjTDX
cRhasXtQCHv5n1IFecsi+bkqVkxHHeWz107mx+YxSxVy+dTmFQ62/EU//b4nPvIb
t8b1U546w72Cff1Vv6HZwAuxMf/D9sJOfEBhRfcBscpYaHUUYkNjdmdp2zbnGB4e
dWs0EVAlVk6brsf+DtwZnxIKbYpolCAhTpnh4mBCFEttMNIWZK4GyTHitUfIuHC+
LNe/6em5vgZU+LDkWPeM7+k8lFOEnzlSxFw49Z1jyxpKRA4pkcQe2QQM5q9RCWrt
uWlQfqcFhgHY8imUl1b6NhHQ2pd08X3h2eQVWf2dZQfTMgiw3mJvFg8QHKaw22KP
UX+K6pB3A418zbQEQXjkQ2OhH2dlqhjFdtIUShuUqLSUcDlrYf4rwA1aLM5loHwY
6/IuszSxWNBmieFLEheVUXX+h80eoAxoFh7r3R96CuFF1jJuitoXGb7hE+37JMjy
68pkXOe1ldeFm/PuJ40oRMf3l+hhiG6BNWvkN1LFmTPs/QpwoHDXGRtXpdjsKEol
Bky+z+P9ZB5MnZt1I0IJqVlo49z1OSTLqHZNxzOYfiWmYAj1J6gIjwMrDhrmbjxQ
UqKZ/UdXIKiqyLxjmmBUtr96bXL/bcHEwf15FK3iMyezHYKoowyoweFUGM3NnbsB
c6IZN57+kh5KzpcfSrx4EeWSXni77mw2y9noUKZC+MlOlWyB16t1oZFq771GAVpq
Cg+F1exaZ+m/CXULFDtFGRAHYO3bXMAn0qkM5uIpFfrLB/V0NDAw8kofu58dtknM
eNhox0UJwGFBbaRf6EtRJvspajnI2o4WBThMNsqQOOwpgnetL1jk2U/ytsPb4/cX
BRsBg/Z8dLhFCtkkmKAaJyXGTBuqs01L82WNbH2Qj8jIpubUT6+Nos1lP8a7TTdy
5nnTCDDNMPmkxjEscamS4+I5nl0ADFURIrxGDET4wl3AcwtvD8MyT6oYneRU2CRw
I2ZUBtHjU5Kb9yUZNIj5sOSJ4KUr85TozV8Rx4QX1GJbYjkqitPNpSsQI8ptCMs1
wry0GRU5XX4SvKyPDUiLzcutKHiSEwyz/wlGpQO9LT6A2YP7UpqQgDpFPrGFkuUZ
XHZ42dsgd2DAGnok6l9pKhkz1esTprYkpl2Uam1jdN8Ohq6/pyaIJ04IysUXUl3W
U8SATxwVzKzeSqKFbQmsgbA0ioa2iuPqxCPUoku7Xfr49QWXJ1VKwKi7gBsLgnxW
EN3dTYJoen+sz+XQP/yO7AagY5p0QAt90vSBhRoKJKJNM10DV7/N6eL+keaok0yG
58G1XD1IcRIfL56efyWxPWDvhkOw3xfHprBCUxKP0sX1dLthrQTx0jdu7Q+c/Fb0
pea6R7UTo/C24qF8OqAFMddbv9PPjTMvdAOjfCSy2CJHyVW4dUaexqLwir6lrkYH
N2TwqT5PkJ9/NXnZyRU07o5H/TJY+Juix4pDLw3M6pROjGu5lW2S22jXSO7HgzPO
2y5J/ZYodq74vL9yYfDjX7gSrEWaxgO/LJ/f+nuI9FSleAG6a8CV4N8eP5DZgazB
icY61s4aznUTdGYdv9xC1V3eQGUTw/8z+ULjj5zssSblDdAXtyiN+ytUVl8gtQbD
cbGEjfHsnt5U2MD73uoL4FLqLnu0CC5H64wxS0DGGCON1IygmcQMHzaC6EI3wL9l
iKxTvfIhyhCI42HKrKCuF9kwvT4mI8qjBih9rK2f3XXeBPoTmX363tISfWeRApx+
fQMKQKcHugSCJwMEFc2A/G3rbeHQAqViif/gPnJd6S5I4gIHzWy0fE6+LO43foWr
ahXZ1HqbIG+8D8ttIkJp9kNYXEXrrxZmcccsuhkpJVOEf3FXtUbT1/z6KK9E4CjD
euROhOw3/47VVytGeIVRJySP/UHd5mw+e997Y/oXCgJMqsoS9DLaPAxirsPXFW29
+PyyOWoapSdqtsZSJN/gU58AEhXSgKODbVGQEd0fa7DBUPqZPEL19T7TDHoAkm4K
iT99lF7AK4TIreqF+I8Fha9A1o65fDPCc2qWrcr9iy+BaZVEaIjsWCddUkNTeZ6I
spKhVcWFbraS17JYg8a+eDMz8VISiZT2gidrO4YId/I9HWlxqwExCL6UMFc5B1mS
Kk/XJkV+AtmhSDp7Rq1HCKBiOjqc0AVAUNGnwrshd/2+5MQV6gxVMqVeG801whDB
EEHfaL0BCvNKJCF6Oas7QdtFv+zxTqRsbIysmt6yKH8sajQETW2t6b7VM737Iy7y
QFvcumHTUYAvOsEG/vIWWaGa8rmN1wreGrPYHyI6e0x8vV+0gJcvCa4lBjpyu33m
X51fUZFO+oWXjRrLkvyRdarI48LCAu/mbigeXOUUqPIQUYO1GyKIgQ7cp+CgITmI
lIyBsOfqUyWztNyl1D7ftm64TsS2/dHQICQo4CPK1s6VueZWaeoNFhyYPQqwtA6T
N5f2890TAu9pNWSRzvvj1TWZzp/ruV6uVhNGQoCltwnbNc0bJpPd/jREoPBcjb1h
hxI4g5NLgT6CKpQ88JVXIfaZtio+0LnSJAo6ztUUKJtSNsh5u1WeJMSDS148FqHj
d46VfNxKsDPcfCPQKbdsSuuGH9bIg6OnUV9Qa2HEXqIFMe7i04qaWx+LGQtHyUIf
wvZuFDKoIN4Yv5ZiZ3TJKGkS1wR51pKc4gYnMdgv5fvkQRSd9G8NMm01PnNT6/Si
egme03YImPtXmnXWkeLurnU+3VVaoF6JQpcpynlg/Xl5ZzjUVmS6OEQo2r8BOwbO
rdwSQoJd6Dy9Kc9ym1x7UZBeszXYYnuY7ZsCJJb2qFyAZXBSMTkxkhyuY+fb3scm
vE6C1g52s9Kuxsy9i8cc6FWsLGBPCOaYOVSjbndgrpFBq65L/lR0WT8CoYR/ew4r
VbES1TMvZjzK5o7HyxR7dsGFZJqVVdosS6jtYIPoJsG24vy3LPCEHQO7miGH0rX7
aQB+4ARRLwPcPfiqcewpJqCwhcp2SFqD377GSD4wsVeK+yfZi1MQDRbrKp9sz8vE
yxCfovr8TI5P8HayzmjCulad6JRDi3V/y2BEQpKQEiDZV8kjqq0aS8+dbTmxOuF3
x+ojDqCZmsMbwI16dGVf8w40GSFL3NVapaSwX/baJcucmvrBQiXozYYOF/H/kLlx
na/lGnN2iXspEMcfkKjzrnN9Bii/2hqPUd01//nByJlsIx92+1KA4aKNCrGypw4O
r86yZwsfatw/Ymce2JLzSUGdzPyZiybRe7/QKui5BAs7pdaWCM3tSyc4FqeOYFj0
j8MG+kgzsx0yPMi1pit5k4t8CPAD0sZq2gpERSHNfB/sUXBp0eA7VVPf288GghAa
0TEY/40Kf4wxU7zbrr8TtbbY7K2m64ZDk6rtPA7kHt9Hna2Nv+j0V/x+Fs0WRTcp
Mxj7QjoNfsnjhdVw1t61xtxhzblySPsIYPz795EB7aMPE2QSBMxo1CR7i0+wLUlU
kE8XLQgBsEebLEMgaLnuT1yMkxrQ0v47qvYV0XukB6fCyllMfgdISP1psjcZZEd4
/dqlsVkUfZ+XoBNUVCV3DhgOlm6v+g+NiZojgE6HlgPd0B6cQKcmMnGg/bHFnOKh
dtH50uefqGcXPt+/ztWUS16dH07wDB4kBjqTOZFkkIlkWZKiQ8+pjNFKSL0fL9ED
aJHdf0kukSP3tbLgqrWtzbVYSDep7Pn3xEorI7zfRJyHoqyl0vKfTvXMPY42yrFP
BsxVcetdcNmJMD/QTZVMLvW1a6Wf9g8yxbwDloOjED+ae8YWR6cQf8LK4amYb26K
7Fu1Pu4o3JCi8t1LCEtjlEgqkVkjgDSHMIvUWU29sHRv77j2Hvm3r8illPnzCh3B
tuLx0Ipi/JsHotWgQRE+uNkOXpglIR1kJv9Jzt6q2XGo3/beDtXE4j2EnauKc9Oj
puitdryIgnpzs25b7Q0wj0erTmTwlvK2aG4ev8w68UbHo1RVjXEAcsjbN0gW2ryX
Ye/HIb8Tke1G612GtQJOEQz56fbeAH5B9Vmd6oe5poQv5PKA8vBqLrT+eWzpwY1s
WwRYc3RylLyqc1sVf76XpgBaEaacp5jtX6lH7B6ohxO2KiMctBjxObK8+q/UTuh+
EjPCH5xXAQF7vKd/aeRbPOa6zWt1JFHb9JJpdtt8QvurLBzm9vp5j9/J+NTTKheD
+XLgZxNOXFdqDfbxJFnRK4wGdEPU1P9P3RS/w4pyhUcLOWf5XhfVl3VR1Nsq+lAp
epmyvIXyhKY9kUhf+Hc4ZeuO35w9GFNssNTcDJtaKhz409iMHlDWLiAAo3EDClPR
zW1I9eVO4r/e9a/Tzx8q7xy57aQ4zQWBm/CkSVZBGkDMUX4iqHtnUPZxknNrzcxR
s7QSG2fZhS7FVa1Plx8ydDAckawEbActMyOWl2gZwW7fqP9Mo2uF2GHbenofL+FK
+qUroRTHDuEqF3cjoL8qMliyWCqI+in3b6gbZIuIOSfumCQ5M83irLAwP30aN9jq
gQ2hHeGBF1OBTo9XOmdzh9hsx+Gfdrdkdhr0fgzFYIrO/QWNjc8RIaONtVpS5b+O
6qPZpFi0iB6ecO5Fp79ZpwAtQtMy2u8/EyjIlRCOBT0Z+ur9nRJSVsmDMdEfalGc
2ljRdovZTtvdnosdAKKgnaY/SEY2+A4/+EWzQ5xcUuvVtm8uxyT9AM9A7GBQFJGP
oX8m8DSlIdwuKaEQYPI9+1O5+KnLMThSjfh2ACM/YL8dP8ErYCKuQKig4cZujgIx
meHwSrwIZCt+IqhNL661bbeVaT2aPsv2eKOV2ifsV+in1cMSVnXskWCncfhXQoBh
jsJFGupSzMtklTu6lvRGyOfuqs6Q8ZtkcUc699wtVrPRAt1nvIqa/fSjYIiLIOv/
323SS1E50TQe9t+4bmlpgHO855By4YmibWReeZ42PDHGDL7BrtOwmMYEdAA5/dSu
uYRnheFpbL2CLqYCqX38Tq2AW7Zin4rskr4V/fIuLv89VA1+TkgBRM91V2ge7ZJE
K2k2Mgmood8lO0jLSI/rJIU3PbYfcgzY+KVNaqtqj1Bymg9skmvIPITe3nDg19z7
25UMQfrIwxmRmVsoZ8Adl/9s3knARv54CdRQ6qgrlYPzv+nmDtee6R//Bh5Lchdq
Fzj89tPoq5EXPSz/nkBKEPmB8ji/YFvllBDaNeZ+duv1lXgnQI77GJMTYvI6GEwg
eXAcRuKGOmPnLveUt0eJo6Wv1t4rgJS/r8MWLQYBcpnuGNXmGHKYamKVaNEJ9scB
jfz1u4rouIpiy3G76SGvE2QCsgj0MKBTs+tfjziM6FPT2/O0QX1K6M9OqEGxrZ9F
4uX7ivvB4XkEgkpsaTpyNGfVh3AHi40HOeCsB32jPL6HZpiJHEvn6aNk9j5BwRl9
4hmGuHyj1wqjf+XER89UpF8p5qxxGh+ycVWrjOAL9bfLMHUllYAD7SkiQaFCU58v
62oiFnjx91jk92WiBI3jHITuzBBI7qzpAYCG9GmKRZJLHaVjrbxvz81KfdUhaJq1
wgGYSQwAXwQyG+dO95i5U3v1Xp92luy+I7X7nvdKl6qWQV1K95y3pRwXlaZxH361
DapqxzqhzWz59HtB2TBCwCIxUykEWubnPWFTsN5DICnwQ+6WqpzXs56lJehPU3DP
dUSQIz1spXBvt2/GPmL9ee/RMVOUj6gc/0IUBxx3WOZISozoaVmKBoxkIGUq7mz9
5YPEvamIHozhk4n47cTHTAfrCoDUpLtAnXkqwK+K55STeZdXzRsdARmnQNifNxr2
TbdK2StGQXwAv+GsABzsRZaq647avbOf6SZrL/BDRRCAimv8tSiHWIpNutfV6zjw
9EPWjSQO0pN0v6IE1rrAItJoCpmmN9oHSf6SalRMLAZQMOuM1iDXa5cw5+6YGYQs
35FUMF+QLw8owJB0l9Q3PSsoH53drfXbYsH3iC5YJhlHrvNMpjBU+lNqsv/Zl9le
HYxMIX08pC/iABX1rFiBCur4SJo/HeET+0MDW1uAmn0duDqL+8vbuI8y5v7UxSUr
hQyrDwoluw0i6DAbLQFFEfQG3+d4kgHkrJLXh/th9jSoIWzOuHgDLOqmaTUBZrMX
i5DMymFQkDbO0wkWgulnGu8/RF5Kk4AhANuzp/1cUqRtEYyjlv6+gQeG/K7mDFNZ
J5cziQDUnYSebPMmJhpOa0PUSpDuBy9okcZkkaCpKfiXELp8My6FPbQivP2XvZ5G
3WcFN22BIY3zf1T4ocetKJIYJuxerQ6ykgK8A4Rjyb+DSC+feNfZWeBZzh83PWLs
wPXEvTka5Po3ZmB4gyhaJwXJTs7WCGnBiDj5kQIGU2zzsDcl8rWHNmu1YNRmFnK8
1Gr2Hx4d3VGnKOa+tQDSpqdDksJfgyxY88elQg308jv7+/S8ppKdUb/m+EnNiVjO
QDMIRkrjk9CPCmMPlxRkL5Y7t4g8EIg167T2gMeIZCBeI11tnQ8mciDbN0BQlsFI
YgikyQA7brNcozu4WVU/IPW8hg3KqChhQwfIZcoOzxxbIHGOTDvVqlI82+hFR24a
Zab4W/agFeDkMTYER98POLKHb/7GprKlUk5Yn1TGzEbLfoHBIQ5n6BXZ2Kmfndz1
/A60+j2v3CuA3wMwBd26wYw6UzxwsXI6Myfmk/YkKAz1KtXn5uZq7cb6gVhWdzvr
9dYiWPmrE6QCZGGAhTJVuPrrYUP27TyLCGMEY2qaoCiJWpowcf6jp4hc4bmws0HM
RGQBEr5NbMTBN5Gbp4J0pRokPEW+SCZ1o4ndJI93I/RLuVB8izfT7++p3fN/LCIc
wnkF+autnwbimEf5mgTYqukR0RRuNMRXtp15IaP6iXY694j4cRGDTSN4Y5qzbedq
bNK8hrx4GzRPPXCwEzDuU5Yfkvk0easoOacDZYcSJvCaEv7u90o2zWA56QWs0YC5
Zg2D6n72arBbU1F6Ulybxb9ZW7xlwh5QtcoEm3km+l2ymEJJ5SsaLOfbXA+MeNvh
Yfs6nANVKqqeh7ZUeXrKFvRJIZ1jXVWV+AWxeWw0WkGMJfJt76rG0IG8xPIj7rKn
BUnfQMdd7vwXtUSWP1oSGgN/VfXTd7y0XfsbKn/JeHsbTbd2VoH7KIfLZSiER1rf
q6Dchk8Jxo/4II79Oy5/zvtDtXZF3WmAZoTgaNNNAxMiHvQGoGBkIfuCeliQqST7
8KrpV+L1LWGYE33kP/8joyQgneeyTGRREJ1oZ6nFsfrcYb5bqUSbfeFLJAoqEeFZ
Rf0vAG5ktoDyyMTKGx3k/paBCIxuOsL9xBneXf86fo96ySFMiJqftPYevcx+JB4v
VPhIZzQxDdsYmBaRGy8cfmoGAizTllZ6SdD3Kz4x1cXeluEjm2y31qA5wUuHXgJO
/0ZQoXgr1jMCw2DqJJ8M1icImzu7RMSMwtoO6igP7mUUHqJdlUEsC7uNiYpByjqb
Hlhh9Z2tk1HX0uXTgCVivlzgw4Dxl1W3mOyyG4y/STgVRYCQcXfDy8xvBrX1Gieu
p4asabkDKm2bBpF9ciKDXYwmhB5zjEQY47LuP7rTLgOb7iAGSvbxCWH+ea4zVfkR
+WLZJ+f/C17QmGqQDdUDGuhBzAr3u3kS1ezfQ8pHAIlfUBUuBDZg0X/ZkUj20PpN
PabnvVpLzqOYJRlPA6wkiCbW9u/LzBHIWPey6In0z9E3d+oeoOs4QWTQION6hXiW
sKAjcnZOgHOvQi7mc5R0rq0/ZPRH1JHfIt56L1SSdXkOCR6VmSM/z/81C4HbliW5
9ts6+RwRMgL89AYwlj+4+31Vcjt7E3Z+ZYrToOpGQOKTn+iTzrcYz9FgQU/Eek9k
tpf+SSZl7ygzGn+aRGe0Vjs28Ianb7XnlLRBOYan3nVRJp62HPuWrGu28iyvuSb7
pKawY6/4MefV+V4rca1RDfGPzWoKJoDrq2M0dtUDI4y8QXBLDD5P4pZz9OGbrbH7
GZHl/uEteXpUnvbZS+7kN3VAOZFVtfYontNlVFfR4jUs3skdJRbqXsfLkJ/5C/Re
7ESLtg/N1b5SBvrhodaUkK4s3Vjf8T0k4K4sAplsKkmOy4jsnxVX8owUK2HPIhTl
HQlZd3rfVykZRR2jFS2J8APoTp1rPEPB2IuAyQ842XxRvyneu+YtAQAcO9M9P4rS
HYWZdG3gwyEwPcHkLUwbtUXF86NhUqv3uj0UWUDRL/JnMRMJ9SzOz78gQ6NsrtGH
rQJqJkNOpQIo0aFHo4D6YaCXMJi113rcDce8gfTa9yPc1lpA6IAAtHeIYfK8zWO1
5usRa4EkqlgZy2MW8O04GMkw1MzHkCXqc4UjEPeOJ6FIHpx3o6ID+WMmglSfr6ek
BDWddZ1moPuwS+EVDq9X2u8pd3T7gCCvz/3fKWdOTYU/nYOZe4BQ6yNMZyOaqZwF
V7MK/5P27tcNRP55L/Rl0wwlDDC/YNQJldq2m3fanMLz6YDgn+tbZv101nN75y6c
ab9ae0B+jJECtPiLnAv0IjkxG3ruwD7ibJzbp/KEQbsxGn6R09Y+k4KjIRqrGujp
UxzyX/jUSKLTQNknPVJFQrU4w+4WYBoNVMtJnVWgQhrQ/e0HcmY03wkRYBs6Rx9Z
R/AnnFJX6jfMGSdOxz/jXTZhsNMBhjcjsd73CiPTSMvOgx/BeM+pouPUy8synWDX
gvFfZ3ZISmqRWQRA2NCLlGi+i8i7DIZJ2OpnI1Fe7yoPym2dv1dwycoebuNOGjic
Vy+GJwq78lTsJl+G09YvKOVJmvxulP4WMYZxhysjyaorCIuiCUT3Fo8/Er5WyyNG
gGofBxNJS3EIJu353ZNl/1dzBEBwotwCDk0Yy9bXbBIc00pC8oLEI0p2968/F90H
rg4jIxIvs409zJFOmZc9ToTN2/Ej6Ut1dQAVCPRDTj5fpe8sySNmf8ktXjEIbN9O
VYMqSPfT0AaC4DuPjck4z9GQLwazd80LtQfl5JSwKyHMLTVDK0Ffo6JmjS6QFly6
DySj/o91crdVgoYvD/Flw2x4SmCsU0ijej/K86R0I93AsXFXhEfHjtjd9nAKH8mf
zXlBQ2XnjpFjw5AAYInYpGHWDt1nU0bXSgsubjTIS/N61+mld/RvfQSZHdkfbppc
ihBIftUa7iBJuDcLHGzrnl6t6nZfP9CgN3z1GcZ7bCY6Rt5uzkN0aZK2LGTXcjjo
LopfwguSeQJWHeeCqHb7RhCcermKC/I1bWqic4AUftCAL6+w4SPcP6Qi4YqViJRd
TGfM6xyWXpCAZONtwgq92wYsjfR4QdiY+h9P+IWIuXV0qmXkwCrie5ovy17iio3X
OFR8/kU0EYi36C5t9iJO5nEmYsg7L+ZQ42ckyvnJggAZhzf0/SzMM5Av0fOo7Ers
/fQfLLWibIHmfYvBNUfKrcrJB3yplbU2zzhYWx1VZaM2l2n+vyl/Dnrad1ZYXc24
fRkte36YaS17CK8x9qS33t6whz9daKvPF6M/fRgE6SVWzxvTEl5ZS+dEr2r9Y47d
mo143CkTQW+cOedB0rP5Cv/nuCG3lCY0lDBLnyeZDNwy5pUO2LO467DBRielOGP7
0JaCysWNONj3DBM59VJtQ7hMVQ5jlmLcvUUwqkhBV5gMgMlY0Lf039otwdCl96YJ
9vzWVV/lul4YXlNolniPNLYiZS9mNmCsyaTMZB9XDCty70nxbIUoPdGlsCkci8z2
mnGjeUcNxYuqB6E6onTCISsGuHENSCtCskmvpSuoYURiepHCf4HcbaWrARZUOxFq
VpM1zAoQkiHVO21fcObEv3K6YnkLAA6qxZ1EIMAK8Bq1ADlOsHGTaaSMhtWfqfG2
w9kb5HVXH9d13/JooDplaHqDd889hS/wps9x9d3Wf6iYaHbJWmswEQW6BkMM+0lJ
t3gVPm8a5U4jrmGw4u7qiKV/c4CJVBtPWPBC3JtFfKKweDrtC0Qlzjw/wJE38/GN
BudvbvRR0efsVg17d8L3WhgipCBgcVGKBgbtstMg3ogdyr1HvXFpywdg17boWXv8
fhkdhDN+skf0BAzIeWWhnksPFIe+iA6j2zlV0Q+JffpoVSMd1+rIWG1smoP+H6ta
NJL5/piUBa4Il8iHXBzR2BWG6xqsMH5R+Z/2M+RfpGbl+LR7O2uU/CaEb+lqgW1S
48zSElqo8ystluHknHqCrJRnt9BJzOcX7KN23/Nb/Ma4JCZMXXwMdbgo48c6Aze6
fDlxQM9t4rkjvxYRmwwNrVwi3/Cm4YXaPD8JP45dqobtWaJBuOsMvlAOoirvS5W1
QZFoqL2ftBZEegaXJF0X8Bj3RjH23i1SHd5PfPw16iBiUkugqfvvdtDlo+C4AsGU
WMMmVCuBIcxS1P7J63JkIUP+Cg0TWJyQCacy8/bAsCwL0skqfF6ddcAkHtA9q6bU
2sC5qeqgB1JjmYrkEEtpRE7rWWP5sOfWCncUJUeDaGoGYtGPyRnSkbr7acZWhYRU
18bhCU8UMDAJqa7wjKqTCIMuKHLiwDBArXnKrHUfCntzYZz3NOdXc5hJnxZqIxHh
Ryg2m8TV6D/BLG6KbybvQyo+3FZq/OL04JLs4wdPAHN3W1Y5ABm30xFdo8jQNLWq
sS79yyZxjrHtsVc8vI9aJd+ogDkpcikj0GZIEIR0CgCcCEzvBJMaiRt4eoMTOIHs
/4BZffVys1B+ENDF8/QgJPUZMG038Fkk6zUDSXlmMeiqRRgsXX/LMHit1VwiLpjB
twXyLJ/8556z8wV9zKgr6KBb3T4R5nGkQ+/ZrD0DK8zvX6Y07nrZSi86gYJadBL7
nrA7QAb/eZi+Btk5G24lWi2+hmMAVunQ4xhKkuIi1LGjJBFcvF+EKR0UA/jIswqf
5V0ElIpJMWnlalz/8jWnAuRlAJKvWnXuTueGbdXtBgHNJlS2IdS1/BZIyiPvwMGM
JasnzvDtfF590WB7jds8V8uiFXyfPtc864RnKRYGN77obQA2kq5Ttt/S9aSVvx6H
I20NGnZI7ZXCphPNIV2Gw1WAaWTcNHGIrir+BIXFi9i7BwXaCBTzftIm/4mGiVf1
S2P2YGTQ17NGaJLslV8KvmWKg/KxFtAFBp5/oa6JN8Dp54yEN0xSMhS+ucqzEvWu
tSsKmxODv5i38E14nAv2Z8S1ezlQdmV8CDFjplEU4KSpdz8S9szrTXFkgOef1Ll2
4Wa0dnk19SmWBM66HQDPCFJ2pDJqeNkIcdiGfS8/xWcoMTWRzlPK5HaU4SezE5j0
6QPP0no9QbAN9iXekAlc3DAGmS3gHXkWlOqvkz+k3MLlBUMp9LNyLVM4z15pQzij
uCaryySM2RPTn2RsdcytOyCEGisMxyFsEexaCeHj1GlpMpKwD3a7zxL4k7gkKAhx
UMNclam+vSjGZji3rDbUGmiCwarDSZJQNNuRPYk3raaUNu30MyaZzf5QT1nIChCG
JqTVMDZndzPYdDYomp/PIBmWp3UzwtjkeH91by38NJeBVf1OVU58Kb3/zXRZK+K7
xYSUBZIlJKIurpG+T/lSat8TGnxikr9k1N7cpiHXlact7+fuMXlJebwdtwWT3vgT
ZKMYuMhL6Rf0fQBKPOTxbOkKDk+pk2FSTxk4qV1esoPgK9swkkcnsv/hQFhaW3b7
ZYUcNGC1ltlS/1dAgsdw76jLOKof6WjlbtrFgQfJKV71P0i8ugPY/U/mMXrL+7QE
NlRTPsmbij4ZxjRQn84liOSUqXLwesGQaUY7ATcL8GLfGJ9WZW5z1xuNFp1WRa3n
8aBAKu1g9DmXQJmn/tMIjYZe7PubMNc103ycIfiPK79u1bmu67yBS+cNkykGvHMR
8dm9qWylQFaXeSVQW68eJp8ofXjb8dpuvUc1XB40N9T6W+CkZ86niTQj0T8ZtGP2
hOzFoBODg1vZ/kiFUaxz2dwRaoUyyHF90De+hbno9+jaZZgn9akaMaLauTSW9x9U
LvRvq2kNxNoYOPZanli1N3tCex9fxZLdTWPkx2QUrceZ93ur+BaVIdRk6C1gSXIM
YOTNQesf5czfH2GUlZ0Ariu16HShF0fPGqvf2ik4uGDQXCL15O15ocDJH2Sp9MKh
JgUVi+GSlcpMyOL9m/FynNEdv+wL4pqA48+Pg/u9aDIXI4euhlg4RkJLfCBXxfqQ
h7mQQSFQkAqBwUPf8DGPKFs8Xo1WxZb6encqVjXNM0PhHtWJK2nbkaa1ZqzEXuaR
JQ6+O3CNeg/g/XPwHx4M4EiyXVxcUowCKDpWuqsG4jKmhqc9X78drsi4oCFjHoWQ
73klK57wEAhXjCBTTY5L1c6Ah7iKaY8IhNE8ct2c7Ozj4I5FXulngXKbLQvuHiHL
NVbrG3OnbQG4Bsy3KQqoM7Lwcxm0THN2aTaKbFQ0HQ90Dp36ls9DEupObN6QwS+r
LGQbz9fN80WaslyjvJdXCsGCyusj4BCTmgV0P6KrbEAclajJXpXkgR4/WBFStTTG
AiiKhgZw0LhqO8Ohjo2zbp/pd9/w52r4mNkB8uLW5YQoJL4F0Ge3YO7wnMZ+R5r+
3xma8QE5rRFV6rCBzmr0V0wi51XVJxAh7h2Co3oQNuEfAHselyXgNezrJBbfxDw3
GVGgsvLeDp8iaWs1mnomXthbtfAKLcq2Hwy40iZjevqJGUJ7cRw8lJe5zaoEXsQk
q25zMU1gwRG1ZmWkdy4m9D4tCZnUt+TbwqrocXKBYdYR74Ie0rVTKu4ltDX2s0xx
0lEHXkz8sxMbzxdQG3Hp7QhEqPV1ca30/gNPMqREs+ibdcwec1O/g8vs5HhD5DRm
ohj41ghBjpoio8AN/llDlYjnlh5zh92bHqCjg1ujQ10/ETxvv2007Cvo2U0hVxJd
xqlSDkRuU/YK5L1w6n8ZaDpK1ge2JDWLCPdmzsIoaR+aEYdccFKr0MTBre63DYGr
gQJatiUA1z+umr2KjSXSopcgFTQtthQJ4Q9Jds8w17R5U9muH2I/3Dr2VAaOFAix
AZ111h3wZBM96iaVQ2CcOHuA2z3VJkUp+ADXnlC1zXdiUvLa2tRdRAJNeqIEGn74
PiT882ygNu7AtW9TC1aXYNL6CnMbucuyeSruOaiQaw3q4XA8/ES2MlXiZsj6dUD1
3z0MCmtGyUyKGgDKwMs/bIlZ6yT93Imi/QbafJfTaz2NgZW4Up6umcGscdQhtNb/
jTpYI7EyaaJdh1OywpBcM/S0JFbBru+1JKBUHDXNHGkuVWu3RbqzW8s+rQ4uP3Qf
y9LyRPAUZI5uuAe+bpRe+0ev6Ntg110XOiLMfcDx+qy1NyMSumKJDF5f+pEuQOJJ
DJfUQLda/rjgWHGV+opQGKvDTG6fXSwh7fUXT33Kzp7L+dSz8tSVdY4JbAUfKNpW
5jO1C3C6a4/+72/VhrIzqkn0Mr5f75Hhd5zE7VuB30Dt5JXtyS8rulSenECXumGx
zRJr/2TBXsDIBJvV6m9AOZUtj2bw3wzQaa3GHb93th1VH4WMKr3hBHCDFntCornG
vQTgVqJ5NcHegadrkGZ4giJ7jqhsiSSM4FhtD/UAXfZjDVeA1g4aSXm+NKzeQ1g4
mCUnmcFx2gGH6kF+3Lg0s3o99NeFrrbk2YImiB4bK/mkF9Sa1Mh/0NjCpVjUhUMJ
NHgdbyCSOJflYPNEdFQMCtVAYWIq6qztFLW1QxZXBNAFTV83tIkmaz0Ffv2w9X/3
+ep9fqRY5yO2oXefsXnXl9L5a8N8E3MjUMGX28KIK92qXJQWc2QDnLcSZiJ+j62S
OZKRxSL4SRlecNBtQPuok0w45aKzOVnn6ypNX0DWqPJ87avUJI3zgP1HuDcZ73Vg
6y+MUBDXdCOBDzmDotkyyRJRSOicMTeIbJfo3/hm8JdpOumlQbrnSlzUhh5L7fh2
jdqKfSDTg64MxH7nviuys/G/el3IZim/HNTqoWcw1bZduBPh6+o7ubabLTKK4yTO
pWyTn/6/3P4Ju0nnS6mguXkyafTHj7oSuDBcEsSlp5phlt1JbRVaDKjxB5yAvt6B
ukX+X1a4llOvOOkuzEu2c4vjTrLeM6nETNe2m7zRWsiU8T6Jr3sbo+EkZyILiR7T
0TvTB5Lp62orNuqVwhlOjKnqv+6+HsVDiNAnFytqq0+udEVTB1maMfoeIUScjzlw
cJuA96+kPHK+z2ZSXCtEUtjmFHYJWANTbducqxxuAE9YyqJOawtTVER34dQ2/oXk
zVfzGAppB8gDE0cJsEEwhtf3XSAr4+J3lDEUyZCA3RPASkMSMKjWpL1OwSLJ+oj8
RvgRDjuS7tOY1JwVC5WN+HWbQt4NyxdbFiBhFklO0d4zA23mCID6+P3PXtb9NTKk
nBx1NHLYxfGQOeHIO209WLxCeQDcSrT4qzh/1U7IQqPH+QIGEvkAk56Gvu59qbSu
xQutxl91Tqu5H+UlpTkEmyNk1ggnjXPj9aXh9/X29GBdMwXOmuhL16qbQ5jkF0iP
nx1TLrqaOdPcfGj2ln3WwEZwr+ciSkzDabsu/i+gpSgrCVK7cQ2hsBFmVqC+AHCU
jo9rjFjVn0wBiKAOOwGGq7gZxhbxoL1C+Ns7nqoSZ54U0iqZrCXUjgzT34BIukKF
qezCus1ptNxehIW8rjzjKlFWaHcUzR7JBBP4q5GgOPecnguU8Ps9tbV31E8QAR/K
Hu0jE9trjvcB2ZmmNwzGPGOE30c0HCTMLDWFHHt9uLWYcp6cuVJFJdpAIgkm5k6+
7GrDQ+nify34Le3sRespyMeWRcrkhxyCLerVheP8f3rYUg2uGW1jLxI3LTqf3O+i
UJaq+KninkM0JHSrnDnGYinlEA24kFTfm1NbkVOowB8CfS5HkEMguAYCudaRmmYo
+2Z3BqsKCZSwxYlbpB1kpKWMtTLvYYW2lBaPjaZPnEYieziYY5/4x+KMf8+19+b6
c4hFedpVIq+9yfY0B1vOYC4K1YnXrVrPbJFYCljoM4nvL3NXYBRcXHjOmb2W+KOd
Fp84ctu+x32sUWmLBaA8FaRQol85YLOs5ZetWNe3uE2KWxBUVhKilwqxjMF2MqtE
MVgeFWjkJ3bHYsCz1Tv5VlVDoc3UXCEGwyO7upv+xGNHRNI8HDzvy+3EI+Snf0iS
BG28tPgYcXkMnPgHyn2bC0FwnjF2eFOyK3E0znTtKqdKs3+h1jq8/etaOcZbIE0l
T48dDKBMTYMZh+dgwlmZU7e2CzypW0a5/0bPlcw34ivFhle7pdYrX7BrQjsOGsG6
Tn29PAAGvQwnpziRDzo11gAZANeh208zyysqcYAuVDzBw0VHhoX31L3Fy5Oa7Mhq
tI5/M6cDMRih5LPUtUPIpSIjTAKcl6MHYQbIOVdgxUxf3UE0LzWEQ9VjzhUtnDrz
cN2AEcBfY8AxAjCGS2tknVWa5X2F3ZW0ybQUvxncjvcZ0qs2OfSxtCxxG2IhdyGV
rJ/JT9jHYg0TyAJbXTWcBzLRRLJE0InNbJJfXJtOhRatseQ3DPjxuijmQub1Hwb7
EG4hdzfDhf3hs99jOTNgS1RP9znH+NnsGOdUJwRJll2Rn8RMsmM2uTOBb+hu7lD7
zrNASWJOydCxfT72oNRvW8mP7M5F5Bv8Vnlr3QwJsGvFVyGZl8/4QpmWe7Y8dAGi
XQbCLdI0F+Rir+9HPO4Vf7GPW7H2rrt1nVR5MEACqlC1Geo1if1If9IUyzgb2Ev2
qxMPUpdVp5Q/iVf4NVUlye1y6jgpgdh2DaN6F1VBbUu3sA9prD1uwFC9/I81A3IZ
9pWE/cMlSAKvehg05aBWr3+KcULcowTq683yzQ7K2zJHM5zF6dOd5lLGdITmJyVs
2l7LipPaSzkCKUgXbg4efxu4OMIxn4ZmQDR4FR4uLE2dVrERMkuWVFJEegp5ZDEm
OazXDC8LwHAC8jMcyXghKA4oIddkCcoVvt9SRJfluVNGYj16KlnMhXhJ5g+0oGfL
jPh0TU6maL09gfFzByridOl0UyrCnpQEpCTRivVLWLV7zwOK0hVf7I/gXmpIHdcn
cZgt8272GX4hJEh88USiNmp/6yGjrag9YCgOGbtiaCOaN1QJcwnzF+raIdIthVG2
hQrZdzI7tFgZ0Zp3ffNElhVTJFcosahbE7T0X4LNQGBSjHBM+aU6kZJb+45qVJx9
BF/mJbbu8VaUp+vXHm3LoVrYAjrxaOtZKgCq95cFYdftdXhXvwI3LplW57hOhNSW
EWOOEfOKvS+TpDCgKPpw2us5tzWwIubZHGPTWjI5kfSX3/Uo+JqwSRnMH1ypVpXq
H51/nkhyZZuDJYSvx9hTR0vdwKEA4h4qLtibRXO7W4AsUEr7KBYtg7awBjvTQpCe
FVefd/EWxLL2Wyfv0XZUoajL1wxIlW569Od/y8tWLcZqbQ2EJYNbwuIsIQGAwNOC
SjqrjCE3kF5a6EPlCeqRdpTPe4PL4R5+LekBzVRmOTMsQQcZjtYiKwKvi/NJcRI3
o0oFn4j37txvlSEHdNtC3W+0F5kmqXrFx8GbVPeI6sj4d3qW5VinW9rt2bCbRnX2
tEX3lqDgVkO6HqyCMS2ZY9VwJiV2+W8oqGqyYOm5Mp9ttsfA5uy8Zl7Az28+Thcx
/WDliaQsikqCQjw4A033f4a8QX0RNrIhuSrbOYI58VrnlYUqOEbE22xQkJpzS+95
/H1uMbwuMDorYOhRKYuz9cZ5PZNwJL9Ibn5DYJEkR2WWCZejG6npFP8aNel+fqcm
ARYoqkTNdtkZFqM+MkRrKnOy6dD/D4B/Ju+NgIqiw+s7ORP+sARr+3U+K7IuRcHD
izw0DgacbahCeQstX+sGkQiU9Vee+1Mmm5SI1LEwC+kWohxEQRPUFX/RNL6CJ2QI
Cxz332WdTqSGK3tW6sKyLOc9JcdQ71GlbvhpxvY1FEfHfVh2KWRACk005h4MkMMp
+lqP+3iCo98sZvZhre+PM0Z4IOkkLzBuYUbxpsdcOZ1Ve/+UvbN4gRN04vV2XpAb
R0ze9WbK4rR7z/VBj7Xj3vbWhDmSr0GaLUNtgMnu3vus4BF5li3Aed0a2Y5DRTjE
pti6PeaER+FvY/h9T76J85OQe09A91YhsXrQktqpLsyXPNguUyQ1zSHPJuD0Iin6
IqrYYQ1noWLY1sihptYWwCH+vQMHE/KTC1WKRCk+mTWTjCPppqdWw5CiM1xHUQ7m
Kv38LsISqEeOS+iOPSZXCQG6luOrdFGWS+6C8JVzBkwzqHp91+HMokNzCIKm1/Mm
63tehYhcIHZDSz1DOqPj64SQrN9NyZPp3Iqp6zOjxWSA8zhe3Udr0Y1kaJWfCcRE
Thsd42/3naFht8u8wPrrNb/kECfVNqYHrl8kOYJajLIlHPQNCLCSa/y4xJS0f26Q
pE8NIMPAIqpSo7YsTwOQyl8P/WbmyXD2cP9tMQTog3Na8CS6CEnKXUhv3XokmJrS
kE9ErMBJmEh1Dgi097SANCTonOm3nsA2RnKl/ELL1JFUXh65WmNkjdzgpOFBYYu6
bFINYPMcgIalSBjs3GopwfOisWZPfpZSNxkwzKbUXVMQvnfnthsce7AyiPvY5QOn
Us9Q8ghdZkcR+US1omPDgXQswMX0Cjh6GhLPvwvgMgBqNJgcJTkKs/3YWs2WA7bA
C1pZnfo54ngQfOQhAF1XawaY6mV25XoukZkjLb9hTCLi7/1y10aVDA9FDY+f8uN1
dTA2SBF4gGRMM7CRlFSwRl9t9EWAHzQZy2lfLIG0m2r1di+l0Gr3IDofqiqjlJQw
RD8oyfh9qMB8FlIdOzcjLqLaDJM79Wpm/tIhZQwwOMuVVxmfcxpnqvjYhuCcrO3P
TM+ZclTDpUTPsHKvquCnCjeLcTlnT4SdJcwatErF3lUDyBtLG+1pBKUGEPsy7etN
cCHDpk+h9U8L2c/j2F9N55D8SuMAksvtKh4MzWhPyzvPlKwWpRl8FYUMwsMJeQT7
u/RQ7350e91tw6jpOb8cpk4nuIhspp8J2DiXAqpD9tyDqYZEN0JcNdWsqSxC0eos
H5OVYIX2nPTR4kzN2w4+rWQ6zK5auwdpUG9SA7MupRF0Sx/yupQXtx6qBavfD1HZ
KtzSWATrvTpLvdX+FDdhI14KcQcqSOsLep10bSBMh0Q3BdgTzYlnXgOGmRmATexF
l+0lhyqjzYJbLkR/SBu4uqkTCz+3yNL1v3aUlBK91EJDbWItuTAUxuD7Vmg+zord
xG1okkFczccR8Zepx5v4bVB4/pTN5hwHYWjKki2g3FkvGXZgwz4f8xe3CjxoB+HG
9rnqbZ6SRdamq5+O3kTmDF3u9pmpSwT7WJDJ68W0M8EGbU5vE4hTang75h6vKqcP
R5tsf5w9hz+B3nil1SVHypj2Mf3gSUyeiTrQFt2QREaSMeT+Khm9DYvYD1r+J7Du
K8XBo2aAc0cGfALz509zZUYnDabU5YLjlLFB/S4hTcX2zEEMyBR3NHjAyuU/R9D8
mqtBFA0jfOpk0BdP+lg2tpo94ovuYth0ikVtEF7QTm2tx5Odxw727NUFjT7pMcFh
VruVBmLbjw56L6WLwSqXQ82+dpcwfD4B+VFIcFnIcY9pC+4WqkSLusjD2Rsuv1xf
Ra8yVze86KUa6MszY0TT2yV6EteWIuoG8ByPUOWAvpGNcyWXFFYTDiddpqvrw9Z8
g+6g4HUTb82ABAYtTw3f4TWjOUY5vgHA7ELVheiQYkRxoNGGmRrPZpTtR9V0JGin
m6Xjpdl9xtVZvwip57Pxc/URJ9Sju/3cZrVIvnzb/VB8yMXF9VDmm7TCl2442Fgh
wQ3wX7ymdED+nn7Fq2YQfdanemfau2mh+pJeVNX+vRwFAWzjK1J1ToSDLYT//1sR
YU3WlxdMCYrymfVV3zquGI8h4oV5HBJw3oSCWo9LZR3jiURuPFC7bloUrR4CgSqw
F+2FMrhElMzoyySAPzOekLo4z1KrYVUhlUVDYESEYOR029qya3thxk9jehFjCcuE
kdftsEeOfzufrDUJ2z9P7bDeuMQzAnv1lgOF7Bgv26woCIKjp3nc3U3++p82dBPz
9rWTjuU5pT/8gwv+hUbliP93f71QU1ruXy0LIkY7q+ng1tXsXvyFe/InbbA95t2M
Rc5S9rC9b9tMnhhyvEEboo90T7fy/JhHG4PgR6HIqXXBYWePeRnzXyZG63iWAESe
Hw8ypoikEiXYJboqNa69jVn5PIEXnBE1xOT36qRMqot6TaHidZJMb7Ag33dlDenn
+jWrgPtVp6VgWpLFr7imcYI/hNzY2PpGN45UEXtnfdBSXfyjkG4s7jvTahgOPmjq
YBCsYcfkrp/Ux3dxqtUytRm3X1NgCVHYodvTEY3Ol2UigYeLAp8b5bmzSd/UENjs
3cwoW0ikxSrfFfUVUeqTl6ToJkmaVDM3u4pEGpJk+w200K6PBMOqpsSj4G2265QE
wQKYCm6wFa8brPpbjlwUVT5oNyNNixTpszNrhLOT1XwHaMfDk3QLtbF23OnzY4ZW
A+RVE8idK7tObGL6o5sW/sH1absUKrxII3gi5yy8pbCdIgAt1VeD2nPR16QhK64Y
8bRsrByphBqpxWwubMXHSGm7BwMpbKVjY7fuivZAKnSx+zZMaYGozut0LTDV1/Ll
xpL7UMepse9gSdGTwMliyMMFep9UrD1rdv27QAZqnreTa/fiTiYUklwlF2UnkZUN
AktAsRsH6dJGbw9tpLhh7r5N/mSim6CUiQ5FAiZ96paZbMPTCLzLTP1gpWlIi9PE
vO0l7FtcpoQt1TLDPrJeLOByNGUpkuv1EN2VZ+SJK0H5xm0+lk7vzfIMRmH4Ezvc
+XzQm+XNbTVwT0tmOiayo2VXW8i6nHo8gNgjDOMHzHUXMu94zNq5bQCUynVRPidH
KrnbOdd1RhBdnueFz6lAaO+eaA6TlobKAMnGGWdrPjc6RRQHhUpjWdKAZJTX3y/j
sRXh1rs5N4iPuhjU9Es1jY0d/CWJiv1RqV/+c/ni60RNQoonIemr/FJXY/7T/MiY
hOFGfS5N9KeOpKv+4PW0hNmCgFAHdxxpmr6JwZv/ChxbhocF+38pyOpK3UV+rRZJ
8RQv/Bt/eFcDge0KkZUdoLKIiAl+ozDVwWNnaNUK2H/WxoLIU5F9JvH6ks6oYJAu
hn5i6HIY224REg2KvPE+ZQPOp02aKSK3qhw7IHI5IMppQereo5Ubp1L9w9SHhyP7
tQG5Dc/61mz9NFui5MbCgIKQU0JWBqgatwK7XWD8ylutX1S2rLu8E1SuqbRhLmqi
23KLTAmgu+h+X4ogeOI/A9DlVGvmOT8X96utOvW+xJdxmb3quvCM2YmP9xsrIZ2y
EFlaUgvQ41SLjATRG0fFSlbikfc2H/yyQvxAD+Y3OmWOIaFHYKj3tUqlv5eD05RG
EEgmUBf9oBTDOkCtryGzl3Z3ChGrU5u6c9xKYxIKUsVd1zLBKiuJ5WlV3seL57IB
pCCiuGXC7YpbVBp6pa96tpkTXxZtSbbSnx29kScc9u6iijI/Y6F+4LaAoiVaHEFd
advZTBn49aaWgnaflQUG7dxq4LI27V17YcVmctm76SJL0MxN4WznA1twAvTwYswW
fXZK4yiGd3Nc59VLdpHo0X0u0OsRzQaUEvfz7zZ+ALKFvAHOVW8m1wzIB3xqye0J
GSBawR9NjdZXVlcHQEOlWaEkObCJgjvpX8i/PPFxUXWG36Vml8hLruTrATPb2E1o
jGIZSNzEiOSJPVy0xbCOgksbCEhZGRGSKN3HUct7aqeJdHUW3RTGyfhKQAhHcYzU
auyb7/f7fhVtNxYqOcAopYt2lSX/uFwXRfze1BBQKIgLVyCJ7Kf66JznNaa+Ycjx
/F6yGZEAaGYr0X8G9jTRzYWBvTXIdoWiZYawHiIuhBQDUDSyUvrwdFZsC0RDd9vn
ZSSL4QUdNDyEwlceYpkjVbv3LqyWJoDxVzgE6UR8Nh+R79Ee4CJinGGtv+wE2X7/
pT2bDRZzI41iXHD2dct/TrAFksQKpkwOXkrE4o0yP/ybP4urTu5lZe0f6KOQg7X1
OJaZydZAg3xhQxBH/1gnXJfYyy5TgMr6vgZ8+h1ZGub1e5RRhzxNKrfXX791cTXV
9ICndp4BXjpj2Dm1zbMIBMFPq7dqekCFYCN6crFMDj8EDZIKiftsLHehrj0wDlvZ
O72eoU6uIkWggZXuK7jvX6sNYnQ/5L7ofgOy04RMTJjIViKyZqyeYQ2vqU5kpfuk
XsiPFW2Nn9HN7aNmCRIljIm3ec6LZ3h9MPqTFKmw6FYUcjl2KQUCyI1wOzO/9/LL
R3Miil3SsGEcp9F65NnuMBV4FP+9zp+oxTFIETlX2JJcYbAxQT1mIYpJdoaTgAsm
Ra26kRRMfmA7p7h1EVOzTWjqP98e3wtlct9rSnhb9wupCFW7cCytmgyXumX2fQsP
Kb+flaFCXz6q4gMk6s34hagKQ8uCuQkOm/p2wn3h3fXBibSycXgnQMjOcS7BXYll
9bmNBqE74Akb1fgjVvlMU3/zAELg1XVRr6bfRdqlC3Sf8ilGC7/klQ/15gG40MDw
q4DuBE3RmdcQjlckvqd/3Fg/ujt0cvi9/nIthPMcnDZaUh5y8imWc6XSTeIgIIGC
qUdOfvDJZj9FG3ci4t9OGKgysVU5MmWi+dXSj5Hi1PWwxeVEgBpoo3HSvsnq4WDl
BZvekrTlVpRt+vItfnpwVgK2CE9g0OhoKHb0+IpEccZfCSQDqbnx/KoLcjC0f8Xy
X0WeSLl5nzYVyOYPHdoeMewbVnyqkLVQivJUktnRmDSxMVhCjlKzQlAaRUhdhFf7
j17AI4NBIxV143o02+cEFb+g3OPklE5YbPW6j+iga7d90QzV4vY+odEyAehJ3ZxO
FaXwU6CEB7xRJeqULnwdXvLhSx3X5EnUvv/ZeKXJhgbQF+kgwCPT84emiL3yPBfF
3oAECxaT5tZ5bU7fGJYZDArmBN1us6Z3aeoqazZ6RjLtcQqTfb9/NOKmpTYhiZk6
1b4lMZP/M3WuM81A3WprM4HNvSywZgC3rIEPi4HDIhEJLEMPsBGGAeM93KpL+nVL
37+xovtEuRiCbifiMPd9rBEsBKNlGgc3dY98GT6mLmrDmq9FfbiW18elffX0VP18
+5BkvSaGQQgeeo+0vmxcBgj0RqUKt9hmGciByNaXmU5iACvn4BQ00uvwhbOHs+8b
k9HZbDozaGJnODGjzCwQO5JWZeS05Ky4Eqjb07RfrugMZZzAs5OixjJMxDXbnL2W
MV+E0xhpt5cVszvjE70TZC591RWPkwea/9J6XAMovJz9LD5dfAakmsjGqGdXJpNM
LMuOeYsVuENZY/h6TKzessRotnl7+xFqANkRi0RZEv0aJNr0JH+6pJ27LFu8GKjl
YQnIDBAgkRpEQ6lHo1qdXLuUG/KsH3knvKlouWoclrIgeRoTJ0dokhe5wrRRrOPT
B5ud9SbPTSmVHjHhfKofBE9TOdf8MLRJzVdjM7pVpIpSq4U1aT2JEyqr9lcLxiIP
oDv9VvJxgODhYvavfBPHmBcBI10gtKie7K6r7QimKlktwfFD4/v8owIExMn/Wxyn
SuLAszlpVjH7tgBh1flJGrma4KX0Jz6T2z+HYQxc2PnB6W0GWuWvqsWAUp7fEpRo
uJyqhsbjTj850ULccaIqtshmThzv2OenUU70nwjFRKLquSEEps4Cw5rWKaVc76yy
lqD9RPn4To0zJr0kmPmiT7HjgVF4qE4amfAZL5VZiZaMEjX6iBnFaQCPMT9pGkt8
Hdlytmmkcm9HMl4O0QeHchf1C5KwSvGBfHQHIzXPb//BKiU60rKAOfw3sUlvwfNY
0emENPjRsIhP5D3owInWkF/V/8/GL4JGkWbknQRtCVCJiAjJqxiReXs3B/JJOQOh
hqmyD4OS5mvTl6O8Wcz/8vcCK70rFEks4D8Cm+2H13kmxWMYGFuN2qSKQMp6Dm/9
05RWsXf2aLkGl4jg0SCq118fy4tfLirabaZ7TbnNBQWOoIUxEzyKYAYE0PpzU7Cz
0ILgw1BJepktyQRpcgrlLw08Gk7JWo4jHh4YmIyjt4//vhoXc8D0No5jKCw9am1d
iRKc607Ps3kjvi4FRWvxhGRzrm0nm83A4ZjZT1/9RzuSqbItdGHWw7nuF59YbxZQ
4FbwXQ8Gy1WagvIaiPzqRMe2JQRWNyQTuFPoDiTWd2n/NOc40kIqM5mueHllRStT
WJeaS48LRTRDLHy1iIGjOnJVi003Dc4j4gjSC8Ko37TI5zcFF4vdnVTguGMT8BX8
3E/wr/OtQyJ6N7L0RSR6hypXYorUsOxkFjupkp3uEHJSWj1d/T9OYCGo9bKw0SXK
1MCw+xp5/e/hpQPhQPvDf+Bk43uWRUI7G5270LJ9W89vLuLRD9nbb5+pLH7Y76nz
aIA0vb9XpG/i8Lx+CUUpPWwg/YRX28VZhqVy7/AR0t5EPbBv2ITB2LazFs9TFSSm
L1gLhkomBBNlRpdQkMPrhHIT8a4l6twdK/7AZUs1x6pHaywquYIfZL9XePFj6cVj
XnxSNQrU0g8m7BnoBV+5OkAH6NNktOW8FFecDmNh8QiesRYUjloCrqP9H6eBU6zn
A9SBBfbFNxTbgN3R5n6x+0jk9gb3vm2wbU1Di0WF0XwW2srvYke+glmo1GHTduGu
0rqhJVrYa1op8ZPQ4985iTRKD/2NoHb9Zo+tgLYXUv39vlrSl/1uF8jqXSR+YKT8
op+xv7f8IiFeEuimxNQuBtKjbuUc6iDS/tapyMu3Nif+B0JLlqg24J8o38Nr3kLR
I9Yjo99AlfMaomnkGcGZACflpB4P2oa6yG1i8qvjbNg1kaswiKtiDIo/Dsna5ph+
44aypCzdJl8KNOTTJwYvbXPNJAhYBmII/doKwJiKDq9EtzUZdqnapFdpZfw9u1I8
Nlma8RBIoIpMyVvQBR66KkeII60yiIjKj1NWxEOnm++UENM9tSlWwAS99dM2WXls
S4MuPKT9fgF069yQVwFt1TCUnRNkRi5Qx1+E2kBvQccgWyF3K6xgocQvuOxEh7GU
cq/Zdcqg1ANxFzgVSvk9jByK+9YYJjx+poPZbjbrf7wkMVxGTzYTdauRun0v180y
dmgOUoR21B/3RTaNdTnhGiuEsb1Yaf1WV3fUVJKEa8a4nYs82VCNwzi3pj052vhA
fgaODH8s7FLNWN/YFDvQFxGi1s5FDMQUvDq1shIAOmYMEnb7xsTXv21kxgGZpg4K
DNzdkzhX98Ddul9jUiHT1bQ4VJC/eWVLIAeJT/+r1zKblX2j5roHHfmf5JX1Epxm
7WlebeclPBfYwzjKlcaM980R7m7w0aTvRL0J0UzRVe26JctnCfeJAjtgyKkLCc8M
cOg8XLO5fy9AGyApXagt62rWKhf+2LMrJ2PAu60m+oiWM4ssS9cmFWnKQTgblSPP
B2pppl6OPYVGrN5mHD333tAjGUXUryR89GTBtOGmOt1VUiKEOOmNvOBZFZArSCxJ
uVzYUi1k43mRS4yFXCPJWyUHqq6Z4FhPHvaBuIQYxWE2YnwNVmRg/Yx12b4rohr4
kqz4HTCZzsAjd4YxGIRAFfgbu+9uP3UH4bhTSbBe5Ypj+HhMszTr8ocGzy+y+CD4
wXEkmYUR4HmM1s2cl13CUbd+ndSwZnt0XZeUhOxIfCGGNm879+Q3l/TVjaJk6RA2
dkfVKTMNZhFm1sEZNMN/DNqz72LTDksau9EqTME4i9KlL1dLWuh+JKDmqqnewAhE
AnhEsna2n9+0TOpdxCuSGafBy559tKzyfde/hWTWeZkoftOikaC0WQA9+ri7zqOl
SuHDmyFNh10FNb0eNzclE63SAO8cP7AX4eBJrsnl4P9yjuYNwhm75OnQvh6r24sX
e207UrZGy+XI6Oj4QPTSTX4GVRrErbOHItsIsWTHupWNyqDbc38aVicb+A5/R8TI
dOQEvzLdLpnCXtPIvBoP9dS2lWSP4tF1Ahc91kxvlABEUfuchC+b7l+9ZkyNPpyE
glta6SFPfQuuoVoTR+ngKkQiAd9ar13nO/qhfldSvRczoY2/4NiQK73coZaLDiKU
0B/6EJx+S0C0Sda98PEFW6Yn6Tw4hfjReIYdBnLihrKEMw1jk08kvWZvvN6vlqyA
9qBO6hChi7zu4pkS9Q2yIwpLX8J/wPLl7soDHzAGrXrqx4XwLIKzQoCJmLPXL32P
6hXO4kf95B8HLlZRwD1BXtJ1Y3kIEoKatE7j8tiVIyklkxXJ7IylUKEwu0JVoVZR
8AeD4gYFyDFFlk+tqKdy6QyEUqDgwuiXnZ+20CFJJRqyndmY4gtrw8TNmSpUbJYt
MNguR/HIIo4G+EhCkgiqp4ya87EZqzX9wsr+VgxCuiD/ve5vx7jpVoPS1pLyUQnJ
xs9gb1PfyND0zJDtDugM38SIYIUvT+V+2zuQO04Y20ZiaxmFrf2zb+ot1m+NwRy3
zbN3L/0BaAKuoMMHtgMoBcpjrMvCTRXYY1uzKDYGrFHH3Wgz5ALTM5FMr0uMmYtK
kUf/ha6KGCyqR1TuELW/vCLLWbXmrGhlHzzISqlupzbxE1SxsLxLqf8O+qVYUqGR
DcTkbrf2JAv76FebaiN1bqCRyDd0kKxNu94nWuA5Qs13XxsPqLJfOOulLBG4zIZQ
tHI318LAhzcBpmaBdrVNjoLN1YDsTOuPuJeF7CwFpTNSga1+ddV4IQVbAYq5f/zu
b8CeW4YaQkDgFF99m76z5HWk3V62N/7iZckhyzF+h2LURgQ1HYsSRDeULzOcSe6C
idFm+Qnx7ZPrRkPF0kJQuC+p0hHMSlUTDAKVSuFJ9K2TSXF7miaIiSCjjRaHKTeT
/WchVbKQyxzPKvu3vCh25VYn4QVS1BZOGqpx547sB5pe7Bhpw5GHYicURjbBVgfr
P5t51TcwcGTmPX8pfXKD+DN3g6ehiIYavxzDbyIE7/7BSwHZ7dUFTB5oj6QJ92ki
wI2P/22KnF2fuzO7N7JotcFx/bHSVeWhqv9BMfILCYW8Nt6FzkYCsGT8cUSISXNV
GDVyAiP+z23HDs+6yx8arGnYt4rvhd0w96VqcKB5YUsL3oXsGHFR9SLqb5lo3i5u
qOskSQx2e31WrqULQKPIjQAcU5uqmT1Qc4F1QGuVpUzQP7hTRLVhsPPeJmNSBl8G
tGzGLphLeIvxocez9txv39n/hOke3mqaE4pc9rJS99QRJLNWlbxXFxBhtpG0+9Fa
cvC9YRlQ1hWlUEel3CvP51TWt0vWAMsxEEcRvi1flxRK19OX3uxEWVyL+2oet87e
qtoxTaTuSyKHZlyfge+y4zFp6f3A4NJ/+a6++fjvFF1/bAZCc3QJKe5Q3pF6911A
oEzcQQBvtj7UI3DijborysJBcVGpor0La1qWl1DtU0pz2GOGtVsvrkXr7ERmaQLx
Bkeswd6jhVMype4qwfVazc0EuIr8Zemu2rgW4DsZCaSNT6ybi3emYFfIepnEupKF
hNym9MY0G9/4z2SvjppV4s0PDysQwX1ucU4GaUJCviSNEPXIjckmlQ1gmpO+Zyw4
JPixVAYV3ECVQExtWp/owHisv0qU3GrREsat3byAkCjHMkuHaKp/J6gKku+efr+r
zcODhrEJX2k8P9uCYj/EqBG42TOgrH7av2o+xwrItA5Y8PhUiS6FwklPlXhy14T2
7+68GlIrCefsnyNv4/BvGEXrg6FNf+P5hAB1EYbm8B+CCljDlN81EjdQ/SrL0yMR
yFl18XD/L0JQgEDYasNxSMxwKOCXW3TF/kc9DxmI5fEluiHVrijHdNfUhhBY5X3R
lRf5E0YTmsIudrD1mV6nXfAAEVhi4/k+3DqeQtDafIsGaMradm/YOGIa7iqZn+va
N+/PHN1W4XKE21BeVhc3rrOgGkF6AtPn7S33xMUKQtFKeeskPckrP08qclspUMDL
aHT/xqE5L/KAQ9m10woka2ZgMVqsmOZ/jl7I64MeOXeUHkFbNjKlX/PLe194s59D
+i7AWJRDav5/Y/kaXN4EIUWgSzxOjBub3aE6wMcYYbV6N3L8eLgT6mFlUWXF7IjT
FfWOZSkq7rXR9/GV9LETqMWHl8XnngwopBzqTF9tqLoszjiuz6wwCpxOKv3dvgTy
T9sMzxmHWjX6M/LcVGnm8h0WCP77nougIW9vI7I0HKZb87FphtxlkUxIFljGD6sn
gFzgIJ/Ino2X0s4jETh1RIeDI6d+u4iXalUU1RbPBL4OADjf/7t4YYg8Ku/8GQg5
46gGb5jimdJvbiJ4PK5Co4zbwfAuRWIUEKVU40x9VgZy8KCj8fu2nrnUTjhmq1fQ
aFiwKaK6cMQ+vhpL2NEIiW+TJol+fcbGsTMcPyPN8Mwk+hdfr4UFtr/wvsQm4dA+
i1c98gW3mzarjduSxpfiVnXcA5Sh3JoHW+JjNJD+HPxP51+sHNfZ+46AR6ZHvvY7
AER938SOpdDEWSeM+ZzS+VwKY4iSEHkEJ4ZyEeWhCv35bO8L3aAl3xOD+TnBFcqN
g55eFIU6Sqb2hH6WNhrEbWoZYANzGQbSp/e0Wjz2AUOs7XYXnqoL9aBFOJpWA6Ct
zTAzO+Sp9/1rwaqtORCquyeJpue7fxToR6ci0+lwTjPdWXm3EylZusUo7zig64XL
jlUfEltrgjBcOkWQhTPfHLFW8Uuglv0nJYJfL3ugKsusv9AXYZSsFdP39kVKkpM6
BWnrKOM3K9NH/MJ7IjkmfNiseMDD+qhNzFCz9OKv1K+siIT5DRnXlXtWCaABpat4
iP0lYzZN74keOk3Ti9kh6+8iSDJ6tIaULOxnjcefAjr2R5v0D/vA4Qh3JUm9PRVY
JpBPDw3rnRDx4jK9X1C4mllkfi0M8XyPpHVHr1/hQbMmdqSKo5viTa73bUUNOjJp
mcmQ53dkWKCQog5SGGm+u4mCEybhkYBmC2OnxWcndLVCpdU2Jvq0nHHSgZDAPEYY
ZeWHvcbhdDey96O86/VzMOSdKxn/btJeG/vY2SXvmwLBqsrwzSRzax2VDwSpWx54
xebWrr/6WZPVehbJlV14iqx/d4/D05hJU3j9lDJYYurcaw9N55D04Lk0Hvm+oQ1Q
0O9WKn+cpMneVc8MCUg9CxupstfHcj6UwLZjmT9voQLvB+Hqybp+cZNW0xDsYAf6
lI3Lkq5EDcxbTVUuL/DuRRYdztidxPAVjuVg93C0zls3Rv+lJDP7muug0vu4nDNk
0zxhWziQIkDJiT+Ac4ZoE1jr0AzWVnqIqUTqyM224FABXaTh5R4vAi/OAR1O5lRh
XLZhCJQ7J07vKYkMcp/ZDDyfEU6bWN7dOQ5zc9WR/gyGPtDLflBOnDGZu/f0lUUM
1LDVS9GmXsVcw311WD3lvmaLu976t8advlH86Tsjpmrbxg5lXX4sAd56qxKenvyk
B2YdLxDrNKdHFAdXST7R1fZeiMWOXuoDOOqb5qE6FX/iQKScA+2c3UgxjUQTUFG/
qLscvTterPGnJQfOfI4O3/DqPRMgP2f7DkFLvjzzZ5mM6IHHiZMhPWCE5iNXGsBp
x6+WhofX/tESWHfsUHSYyA==
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFVGNCX9S4gRX97OUBq9MdTEViimPh+SKl9k7nMK2QZIg
2I4LJKoPvB1+RT11CuG45kLIOn1JOdbM8QksCAA0ad9D2Y1lXiP1zj0kbr4KBpI3
niwF65/3RG/GEEN5BXX9JzZsVb3Lth+hY0wg7mBiQ4lZ9E10DgZ6YL4u180NSqLe
fjQWOHdoZcEwzdDOhn9SDubvqsr649TgoD1PdRabXv1X+ltq3v9LpM3v+Hcs2PqX
6byxqcVp0ux7njzkwAqNaqJliMA3rPlw6xdQOjY7y1070O77e9210CZAMOmXH9a+
9NphXd9V7Z1JVV88K7o82BEMQqcOZQ3W7492LWSqxzTTQIf1oX2btMpGtB0dm7Ug
WQCZEE+qwHW9Cx+ZQNMMxFOlJ9dIl3jLOgfcqGuK0FiJ4gGO3ioSx0J3w5SFzM1J
s2DBKRL1Me9VhNO5fMNBPmJMiOH+GkznQGRqFSsCdwQ/FQaueRtfX05Qe3Hr26vc
1njEqKzVBP68/JLzj0L5F2fSPOJWiwfBQ6UXaG+L1HnTSp7lEmDIkhs3sydG17yv
TnJonHaDYhyXJDkukfcJZyRzYJnNoxwxrVXK0VI/h2nM2B6E2BeYnYpwFaFNg57K
LTTp9RsPeZfeTVMsdDwa/HhTB7BodteHDShBCDVPU66X6yTDtxvd6xKTsQmVYr88
kZQUKfYx54RSgu8Xg6+feVHgCYXejQ4dJQw15YYcvy2xP8GXlZlYxamJt+9r+9Ps
cqZmE6wizrumm6W0j1PK8cTsh3yEUbmGVzvrqHulBL+GBzb6+vfIIXIdk7Rbigis
JtIsvGR6FEoowilxW24k5j2mgQDFaJLngXtQBPAg1dDJwqOKhnKZxq/Rzy3yVzFa
Ov3EhI8Yg8/RhEP1cHeOWXNNEodNilbpAySdMgNMNhKV9zoLUtqxEhW62giTFn0g
l9aK95TTMp1JTZ0Jd/RAm0pnSwsPMiQddXJjhhlNODzzZGS7gEIdGzqITcYrtWMw
nhbPcVzK9YpkARQ4kAgMnndX7aO4dcrXsqEw2IFBgPdFe4sLEcGxWA75HaVnOJE6
HnFOUwEmS79PGlvnEx0FaeMf6Goh3qP/MRuFij8cWDJk3FTJquPs7GCu74mJXCpM
JuFq7Xoyw/vCnOOFbdhnrlys2ARqczPYu/Z7yrrxpEUzSMAul4+xaOo9g8YUGucn
bkkWmtoyk6o+dvwI+k7c8BQ1u0cQRF9Dd0aAsJBYeR+xXdWDwBGhzxubeI0L1ZiD
EVTnJDCAmynX4eG4qQF1DEMkduJ1QaFOyfL4O0wxHE5k3xRfoNOQJmdNu0I0vVuw
DxyQLvQyOGgcHa3vMDlRKiL5TqHjggzvbDZ4oas8sy65UrL1LVVWG8Mh7UKoj4VX
isMmdjRvAowUJwPJO6vzxpux7gEXyxc8ajqMrDUGkjkI7nWwcquJukaLcVfAhT3F
wFz9LnCU60r2aBZnohsIArSPkoBY0LnFK/MJO8nB4daL3lmZf9L0ZZIJE3yxIf80
mcfWkgcx2Ls9nb8/DDcq/aHiWQ/InyZdDE0aVMvzGNgmlrDtej4oQld3/hVn6Ovc
Pj17SFSTKdZnZ0Jg9+lrnXzKVRmjSJgmNA3utRzXjQ8cPwYElVxMie76UFOpEAST
Rx4wB4iu+iKX7C8zHLTZw6i697drzot0x4sqQS01Z0yE2+3Uyp07FpOx22J8phHv
vXXIiaZIXbBoJdCpogUkKTwZUW7jFocK03SwVcbNBc80LfVE99DZVWsIEjPG3B/g
ZMe/Cq+W7L4H4vZYymKvrdsi+YRKYYgeBCH3Wv9yYHQLDVwXZuGMHSh2DqHBFPte
A6GmbH3wgPJ0ZMMKWtj5IGlRCJMKCn1yAqKQlF/kwI4BhPfy3hiuXrPa/JVNS9np
Dhsx3i/+Nnn0VdOkmIIUbwe4vwJf/XDxzyyqvM/HACgrCVrXfDDq6a5ULZHBW8tC
VSkIQgnnvrOLlf6klgMNtEsMqj8DCp2aZhXeGVd+ac27tZVM8rVTsWf7oPVVefWU
d0UXPNiiLTnI6EAxlbCIxDVTX0fLT8s+pJu2T7O/aIfUI+YSpFzf2T0PmHpo9fFV
uz/ldA+s0qZ7/REKUWTGZoqNE43NLxUbJACspqCAqrCHJUJs+4mzdnAzFqdLNYfE
SqXemIJFLuld2w4KdW64+noSu11YrsyRzsIxD6mqYyIh+6OAtJlFnXfudet/BsKj
4vP8wgL7VcEc0Vu6gCG1i6VPpGMbq0YZEQ35LAY0Jpp5DjfPQQZqPXDblidOSPym
z6g+SoLQ90iYlQxWSNwnUDtk5vYE8Rux58J2Dz1YHoLOzr2AI5ksxvBLhHalvlEC
un2lU5L9y5OsYrEJiE3PfsW64yWDGtFMWJBorqZQmxASTDUFPXESQhy+hkaMEC51
g8aEh8FZa99YE168C/7pX+Ul3EXGugc5Gu+J2nPVXiawELvzeZAWGTkKItPxlSwu
BlRxUTocabQaQoZn3se2YT+tSHSVq1T53aZCuaf7jXIH24erGIk3Ou9YPQasOpAh
YyaB3UnRa1QAKCzKDmHpCWuEgKiBHBWQy0QlDYjHY1vkSVauWTYszKqch7yk3KDi
BsFBOsKp9QiZr4JKV7pBfQeNfA587bus8ysIqdGyvIsUZw8t+1hHn6pAiF+jVEZz
SP74GKxYGv0vM9fFqpJS4PLrqgKQrYFTbx9JIt8lJGgAvsD1uvwr3Xsd5LezXgXO
YnfjMCBoOE9K7MQoOUWL9UqSKN1g0FbwQvLsj+390Jy+G2zFgzROtUjoUyB1C8F7
B9luiwQAD5zlzveZelJKU8A9G6Y8tsb2SnWXvVzdkRsVY5GQ4Ln/gpnwIujKnBZ7
YYk2SA91NK6JS+HytJRrXJFN+OwHc5lO5BynPqg5G76YmOY557z3gSSQI8sd40FJ
9Q4b+IExEZEJ1SETc8mAi8IAZI3O2acecfYQurtk4cZG8/CLr1hXgYrknFKlgRoW
Dthzs4ETv3EZ4sSyosW3bL9i28M5CxQQGjDhiLgWHneyUoH819/fYmXoapG7U6m9
Rl5ZLAmCzDNHtQ4Q2JGz/R620NKyt6WxaVfNoWOWJMv2DDLuEmnT2d34nYaVxEhk
DTpA3agyUyIQGMhqiNFNk8RPUe5o0zM5S7gQvP8PEYS0OzrOqXBnpQrS0e1W5r8K
Af+vC4u/m3UJaHjpbOhq8PPbcqxOq9a9Z2Xhv7VKOkqTCokhmh6axcBXFekS02Ab
TtpgzIRibepx4umBlwlwv8HWJxMklqqW1o9euc3dLzW5R6+6z/du11zGuQkfFTFn
VmWGGWjZMYalCOQ5ihKrYbSip4z6qUhVDHk57M17E4rD4hkFmtuyaImXpQswHjH0
dIAf71IuGawz/7nP8XLfjJt0mMgB3JRAAuHK1CgYB1NM0KCgavQmHk4aFexWuEcN
WXGnV2Mqs4K5M1pNKtH7+cwm1jBU48/FUgFo2gotjTAscAGRiFVrE2QEEbKFF2yR
h5+WKnYJpOlohMyeD7c/lRSmEFy9K+zR8wFow+adZtTblRCVBjgHYilc463FI7ph
KQSH56J4am1eolnP+YCpH7MG8r7o/agLoKInWWHfmVi2SUX7XWEeL650xE2K58/N
cchg57tvunkN2YwUynpynPCyk4i4cANDbzCxTIilHJ2ePuQdDwZam3XS0JI8V8jv
UImU1gc5w96SjFykxkPvQrymY7sPDJHKZdffzaL1qnSd1KKlks+LItzIGcIXV+qd
qYOe4brRQOES+MFa9/rPW3aMN/mZOSAmByJ9srAiAiWf5bxYUNX3UktqghuwrQnB
A4Rp4GrJvoAdQQgNnuIGoqsx4j7qE5jdwhcEqwezkpebFKHKLtdeEmXXH0CuF8IH
IW0aTePP0pKB50pp6MwkI1N9BWEwK4PUfeJGCRCQ/ZBt0pCncpAc5AinkUJkHl6e
nAtoHJ7YG3B/kjQtXEAwWkFAzD8bqBKcMGHuDXlmsTP7orTwiFMbj6NHTx5ilYJW
M50jnj9pHXWfIngEFVuHhoe/JiXtTu+bgVfGUAsb5itcs2huaUhXVzD7BxkBHREl
KZ4TJDFTwS6whJpElBfEetEIaVLh4B+K2lnVDdrsUrhdTkIh/yrOfl0lJCBeSgfi
0DaAe8pyTz1K2Y+021+QdXN+4VDbnYeTuFVCEQldt+7139WZt1VVfO1EF9mW91Uy
S30aW+tJPgJiYRzJmQromyj955Tb9a5ss6dtuOpaQCeydJAdTTlMfWXazqUh2nTK
wE0RhMP34XWbnSE988K54l2TfLInHFlsOU+D1t/pX7U4LK0KD9pLkxBjLERSTOh4
DAgcFdyzRIyMBCvLjoyAZOV/21bhDl+ePVwblwrXBbFzV+MM/1SNUCcTOTz3fIlY
ED7jnZJxKV39/1r2TA5YLftUIJW2zBclEwa21gPZLvVSLctBk7/O8Mz6jKQK+ZYh
dwereMtaSEGOhztu3lb8yutBtNbsODXqoDO/uF+/H1DhTQfH8szmInzwB10BO5uR
eup9GVrNdSDsHuMI6ZBFHddPj47O4wCWwiGL8SqGpz1rRYZcbO/pKG5f2hbTRBEP
X69UiR7iW3UjLbDfPnSk4wUF0sF//ETLDjLtvbeTA7mvPO6OtQ8yZNl2ygQvoktm
zHKaB5NimfegAYkRnyLBNsyT5TT2EeG2fk+lIoDi7dXLuAmc4mT9FllgI2To2dy+
nfzHWWKCLqir/sQlfWH3J7IxP8t+dQFQdnzj75GoQKnSOsMcELzxwHENoNiSasfD
drC42pxaa4zD3loqNATsBU6Ki8rHPcadxUxOTRyRLxUHoL0rQTSyiACsBPUlUU/Y
sKAZqnwKMbaUdl5APHKNyZ/gdRyn3keihPjY7co5I5fu330ptDaU36C+cyu8eRzc
nMe9frYIG2DSyIIVJ5BsIwq/9xjP2PEeU1quDX3H/luDMGXn8aPVF37eixb+tz50
Sm4RnQE+V7LkRrHAhFcPz/MlnYOSN1RaOyr//nj/B8y8W00Su1ElOlZOmC3sh98O
MjtpT7Bp0gmQgP54eoodysh23CQxMk9G94yN6Wp6AhEFQBoc8qZm2I4MHGDzCg8N
pRB2K2yO9YAGAD0xhZIYZd0aDo/V1c1u3eS1ea0QktvyJBBfy3b2iQI1BBiLTDRw
5dEU3XwUVk8MyREmYbG2RpGGcif4o+9x6HASUL832E+fAn4WEDKA4RTi8w0st8Wq
deenTAl/R7zA5zvsFBRKvFpSHAazx3dT48lkGLDtSGNqcc2jtNNGp+pagg5OtBua
4QdBdGCsyUcFXaYFPNO2B+g/Di2ohVFFl5I/cnDJdsjrdOnbJrjxii5iIsHIbFHP
iAQQeIeQORCq8Hgqdlcncdit07k4qik/O2ckLR5wxf8hw07rKVTcdBBrZqgy60Nr
vxDKdq1X0Ph0fngwS5m6IZHbTMtqAQoPUgPb4n8qPLSvoLNBeQrqY8NEZdPucgM1
QGqjn+A2DBwdnwlDMwea4+IsvANyY3xNJz+W1IsbxY7hx6i1itG0eDGwarOZTJVM
C+1brsD9amxFQisB18h1JCSg2qwCQ5Yr1tUHd9mTZvIWmJ9WakeWvdFKIFEkm4ea
FGI1VrqwGIFeocwM+Fyjqs+ekT1U7BKn2GYNPNUAYH4ygQK4aYYFLqoPpeUG9ozl
1ZUSoWVYmbXIDbfwIcDa/Z00jnuGdW7R4thAe8Yzr0N6HCW6H6iYREuT/XTUsjfM
ljMHVMC42GLXbeTAjIm2xhLh0aAnIFcqxmnwnVoES2p7hc0PaL9lJIAnWDNYkUfv
o7LCsUd/bPK3swq3gU99UZvNlazjsiJzmt3RkNsoWo8y9kJma2ftFbL/nFvjjsWa
gZT/bBxazbsTBiWVxr0hkN1jmiSHffz4bg3HiHNXYVv25F+ARaxExhwONOceOYNY
j65328JjUgL8djizHalvbosuIUnUSoQHObiwoUjlz2dyO/xTXp3SQ2npUk24H34R
OW+hjUyFO+RpIyuGz80r3dFCW6TGP2OUGfQfw7Bkp2VpamTwDkGiPLBdSQ3NP1ny
X8DE80+SumAHn0dTh/m3LP+Ga0lb4Kx/AJgiVu/jWpXDLVuAiERA2XLNrW9GAltz
hrCIRRCvWlJ+9gvAQsVmhd9vN/pYJs9Vh5/cU/E0TeHYad9IlOtbd9A22Qw/vj27
5v+CyA+EvqTez0HzJQ4fwzgZfh1HHym9/Z+wZgL9rhNjOAIY+L3TLBbgMqyvQgVO
IBgWRjsvcppLwe1Seq8kcc7Ot8a5lhfAWC9xrjJ45Tvy1taQQ6shHoMgX5VBf52n
1fcHk3pcR2xRgautTUamqOSLIKwx4FqR8tUGEC42RKxqmfhkuemcR6Cj+nXARlY7
5Iieivf/xwAX/CDNYwE1m+6d3gLenVrLrs57Q6S42t7mG/U+Aq2A8pTvJh4tAnv5
Edt1O5Z+SZVoZjWBxkpf/0KiWtXGHvoMtncWDm3rTebk8mW9bPGa9LNjrEWk9RfD
AUXGDXTVcg/e6QxK0TqZx0sOZe8W1BXysYfSbBsBu/v8WdLPr/Rg+xj4lhJoBBuo
ofiYhjhV4d+p0u9hZlXjzOTmNXOyALFIXLaeV3xM+pKwSNo4sZK1bgggOn1VWM9f
Z9BX0E0RFJxnJk6fhUKGALyAtU9fKtHZqop4fA0hUeLpS1ta3+uMdsr6iYidKhhR
eRgV4vZMRQRGkdkN5HpNvuO0FmK2XbUkC6iKPx3G1tf8zwM++fccDRytN6NaZ5xt
ojhTMGyJ03OKnCf4t6ohokdoym8vV/QhJfnNBRGdcoI7Xp9MWFy+GIj85tQMADaa
PeW8YDJbmV/HJwJJOWLx/VXNrFxfZE6zTjY4IbxnfzIMTZLyGsG6uiKbS8xTVQB8
GYGlRodVUHFnqC7QBTeUfVUEcj4PxjODMpfTkFKmft4S+C6ZX5PH01cY8JZ10lQo
hGBMv7jqLxaLJJJEIr9sfOkyAzUYqfwkTaj+8E2yIXzsO/CwcodzxnP2fH1lXXxc
pEjby7VzmxmrF88x1d4g6MVN9ssd5DSz1eNNp9gf3hBGCIuK2uV50R2nOMRRizqP
3w2OSq795jDq5clL7klGPqxnkmYP5nxnTccw1CE82X+0ftXDi2NoVzjRMX29WaEq
H35+3wzuFMR+2R+KcNc75YZ3BPrMBLYzWRMzoGvZtnerOJnzBte8E7yEw5KAtdCG
Np9x0qQV47V+B0J6it2EOS5UdRagh/ICCAH5CwUGLfSOwG0QxQ/3thx2jcGbV0Na
xdrQtxDSHB2yywrg4xD2DwnduGM0bYhXpvgCD+pQ0Kr+sj5cbMEFuVJ02xn6lKWB
0uF7dvZ9/Zdh9hiX1JDXQj+z6ezBm+/lISktlhPwezcbq5T9h5DJV4Lnv9cyNck1
cN3BCfoSOluLNglMLfeU7fEOumhzo799BBdnE0ZIPh01ZsGLRGb+lizdBj56J29z
fi2mxqEG1kT6/Oywp5XvmD4Q6Z55Ch8veh6t4E/sWQUrL2fWwmxfyu3/BmhbgEhw
RTQ4y2OikeYlNy/eIwgi4Own+BSlnu+AJtjCqL5ZJDo2qNW3Gr5EAkWsWRYdJRmF
mdjAP9XnnlNquBfM7ll/YIbqVvkgCDwXIqOw4TBsT3px/tFqiWkhnoKO7NEnBUYt
Z4jHQcC4+bFqZwYIJ01DChmUvOrht1yx4YOyOFpLz+gAs9g27EQK11Vj0yoeg0mP
tzKAy3xjt2CCipPDDcE1XSN/2oZpneN58JDm0XSi1ahoPARsBFjtP5fhzWQ7AL5N
l0qG2NaLaDbVu3Q6A9MR2ckwcvFq4MXYcLgmX7kzl0OFF0sFpJU+vCVnr+u5g2i5
x5Niw1lUwGi/iJp0Z9PuVuX+pTkMhH0hPdXcY1A40/dQZrVTtN/4k20Gwe7dyIZg
La613Nn+qnubKBzllNGrqOIE57zZtStiWESK3r1UOFRslag1IJLwGfeoiO/uqDlA
fCZOkeYSgHjDHRoAb1JnDmhgV/aOuAVEff8H0SO8C+qLLuv7ZbkD7V5cm/EbWcxX
lsAnO3eCC55bhRHGQVbD7JI9Y5gqbZXu4IwTHN2vYb7dAkkqefMZsfRLwtIfpvfd
Fa0QulXkJ4/jUXc70XHHnwvatd1pKJT1BYK8xwLU/3Yti9CH8U3Jh/O8He4tMVcT
8D8ouJzw3GwKeYsR0dPzWDTDEF9E1p5X29ipKohgu/cpu4OS8akwdaQWmr1gxD5i
9gXk/k60+R5UYEF/rQf5QiVKhmMCzdCap9wWqW60ibsPrwAeuT8xKk7TGAn+ZCbc
rwfyoLrw+JKB9lYKk1dJUlx3AY75HOHSTCpjl4bVHkMjT2UP4hhu0wRJTeqkrn0j
pX3eYw2ejua/p1s4+mCxhWPk0RtBEaNiLxBec2eTim1MNDpEXiuDc/U/6zmEIdE8
oC1SiGLDuyRlfsoTcTNY1dx71EBsEy5WwS1cwxNq5D79drPKtzNN3DCycY0VsTrM
3bS3xRudSiEM2Qyjj0bN+cs5h0jyT20MH3GfL0vbFhm2mIESWMqfaG26Xw5hsQJO
768S8P5OUz4HHraBdGOFAEXyDXvlaUvBIQQVO4pBf14tzrRbQIXmfm3ZolAgq9oa
nudB4kHzmBcOJdevQvph2QClsWV2kzuwBBhUsMLfG/ki13UbxjH1w6JBh2pp+Djo
RPNGGhz+cSiPZO2mOd4520gOZu6qg0Ss968YnUMzcPiwEHSlHIPq61Q4PMZo824a
WLXAzSty8q61e9gRAQhntvSqa2aXAtGRhgTiTK9jSNtpscRt6yTCnG6Y7ANf1y6h
tjWfTud0u1GlEt0udBaqxSzhaypZMF0IVKryZeXBP7rW7bL55k1CLLI1M612MLE5
dSd6/CcLCF7whWQriu30Bqb7xGBSGIW/0O5iTOXt8qqhBFCxNNuBb1tvL2MlxgJX
iAnGvt02TYVx2zLzILJvJw5YaKg54u+Wf1UTxlsqI8RBqthT68zryuGwTN08Q2hP
xJ0uUsZwFWi//SmuZBYk6JWoVV0bESCNTowFKmqfL9p0Dz7VNOQ+Q2um6ilPl+u/
nOvUC5jJ5a1yd3jUJ7TN18/2KIbEQeyMHRgT4EiAXVg1R+SDAF4dA84xsJzNXPup
GOZE9hxUVQLSa4KhhR9OoovPVC34WgC+JZU8vaEqM9VmZHhzh1K31XLRC/IXi3lx
2JqDEdW0qK5t8DBjHVi6+e20prsSome6UbHW/HqiJzbirUNWzT4Bpe3L2zzaE9qR
W8gWbrCZDSRDLVNaLEzZT/zq0JoOl8sK+W32E21Ne6WCyH/IQoEUZbNgvo7jtiYF
pBeaMc+TdbrSAvo8+q86zN/m49/iTA7N5fXn+6UkSIwhOv0E6MDprrUpOvWOrV8P
YeoVYHUcD03eZWrlOMKrrLDxcvdb8fDn0lTEbab7uCH7QWUsq+wq3DWStQoDycdo
lvqgEvRoEUQ7VrSo5Yve5Glst1FytpTiUK13fS4n8vdHT+IPAPiKe0t1Hdh4GG3r
uYqr44ScFw++u8fYc1XuaQ5mK8ZtxahG4IpWHf3noQw6vGXlWmQF1eWXkAoIK1Rz
+Bti/fKq/0IgY2y4NwsBdxYmP3WTfBVcfcwYnbAfFkWPVrwUwKfGaH5JUA/l0RdS
OxTVauEI4u95ExK01IAJJTFWJ9rt4P8GqXIvMTiLbRDWbz6xGFFtRJcQOCvQUVje
QOdg8D5rqv5fVi7oSOytvJfCKBoyZkpRVHeh9FRaMpFcREUPGaNqBNgqzZ5htviC
qCeA5djhJrUwF0o/tDz253bOcx6MRFuPXb5RTdbq+2CMNs27aiKE0mr46pTFNnv+
A7PUrbrfEIG1hfnDoVgPnK/0vWitBZuBqXHOg62J2Jr3z0UnJEbehBopAs1L53Gq
0B27jtdgznGG/SqXLZ1V+qng8dXInYRQj3JfIin6wjDNqWgV20ivxmzCZBco6W0S
Sp9b70wCbsK92NFlUAh58LUyeOJf7FQDTlIdBX4/vBM6YhIhcVC0DW9AHwM99OCT
t8+BDUMIuGQJETYolJHDFFMRwaNaAR3q2iKpV0ayEfq12E6BrefKX5TTmQymLhCr
XZAIOpmOvMBWsn4SD9BQ1sJkPvKiUsWOYAxp4Gx4ShnR+r7MewHb8xc6uukxEyJg
2hRJh8OzrsI3bEOGu5nqjdK+DUn2ldAg8S8NVl2slCPo6jxo8lJYs9TKJTxbsK5+
zcfrdLcinxqO+SO9Whl3TpWGs9BEtKCY/uDAf0ykcht34iNq5pPs4gp1+oo88Tyy
0dL6bC1O2qIZKeZ4f01gQSp0KkUKg52zE/Clh5rNvgFrR5uEd4AhRSExr7fskDN2
ARqZeCn6GLVTr3Qrr380yyExI8k/05TBhvyfMMVkZzxEpLXpKe/Q0uR/e4UoUhfx
6YRecp/k39WaUUoBUBDIYmFIW8ifWgXOm3bL6292EQFxoco0wTUTRozj6esWuChD
qKXkNdOPQDVhxsA6wYfUttFc4isPxDiffWcWW3714gkfpiP0kouIJRCVQaqEYa5J
2t4hh4rxYEMIjQhcCnqBVBYLRUUG6w8KReKkv8VB4iRxgchzPJD81DRuH9VwM+xB
lsGbDPTTzdaQeWZWTNG+je5/Tt9uJD1r8Ms2O1unseJQcQbHQuFi3TYDTPE2P4qS
Bq4p4re1f5Sfn7/+vehD5OGjYjqX8APprD3WdBmTnQuC3UCektF1PRDg57AkBfjp
w8IZqnG2cMg7UMEz/mE2BmJn0kFzfxdyHjqXg8xm7v4b/LbdTZKp6kJUO7ZxeMGV
2bac9lkK/5sQAo8j+iQrn25WHi8ZUKm3xi5OhKG5ukVU30IGXAYGZK3dqGpzKXdz
q1GeM460mRhW9a/+wkIla9tU8e4RdrmC2xk7X9UAL2m1O9Z0zZk7qzBLCR/E6Z3I
Rxsg963ataN//xWkbE58JoC4ZsWTXBxiFare/yGxfnEnJnhXcFAlyyXKicrianoH
dd9K04cOvvJjFRZeQ3cItn+KbWZW+ruLRtm5ZfTxbyjMwSXSG9mFih5PdBeauK5j
G1Pzzt4Z36z3QvOlgTMlqs0/u8Dj6khHf84oiarytyAxF38BtoomyKYaR99R9Rms
cHFIBlEmJZxPEHCQzBlqv8mAxMcDUp/pObKvYiv5ruiV5us/wN5dYASYSq7WQ+mm
NCaasV2dhTi8/kfR9p2UF5SwWoiIM9BHY1zDz2cEQiVwjuLm/fkCl7sAl9quQO84
JB21JPQ/VB3UPWL6X6M3uOeKvw7LkUh4UzuILLDhS0SzVdpO2qdKb/u7JCS6jtNA
igpHgAf3A3G0l86NtS5FSb4awxRvotqo/6cT4ogLlE0dwW/HofEh9vR+eLBkPTuU
akN1JzPbH+uNWXOPs1XkazHIvoIaZpm6eTD8tvXrise6d8veF98QmznRc23qOmzl
ZYzRs8NnOxcGr8AASqiOwGMEUmxOm8O5t8YSLC91OLH9uxrmS+wQkFy2aqOzpJJv
qgDZqohwKVwDQp9pSHKFMBhZj8tkaHALXLYs7BwiMXaWH2fB6ZbxWNmpAcXLeSLq
T1E/hbB5ubMOLSc/4wtSfH7i90y+u16TZ0jAP6u/pZKi8xCmfwt88BJnrKKvEkqN
WhY80Mu0tq9o4xMkFhjkqx70q0Vpg4twrY/WZAeyGGMCnlabtYqZ1eE+X6b9tX2N
Q+OOMaGgcretBSne7iYJx6kcByyVfFLMrt2g6H6CdnoJsJzom9MGgE7XmBESS2ys
3msaR7OZx7RFfFOI3/3G7amDubQvv1alSNCRAAAcbpMMmHWIfdJEmTHSeqEl206Q
W2PR1/NdyltY5FwQi8VPus7XCTGEaTbuc9DbiMBcmRsmbJrs8dANexuKFur0Wz/g
3spRPrknBnKBsKli9O6yb5KGodqnlMUmxInDei1VnmAveEsS65dm91xljmjsCrKF
K0N93AKtofihJY8ZlK9n3wULpY6Jp1uGStM9Mwu7ASYC0mMnkD3ECmHf4l5afq0R
7f1wWcY9nUStrwt0R+sQvJ8sg97YONWbAa1D8MMKxY+AITvlF6hG/Y509a2jWqJU
B52ecCrjRqO8LZd37Q62ByUHU+M680m6qVP3qsC3DcOE+aqjkLL60lxAyNbQ02QF
W0Of7AJn32CdTb5HrC6Gvcu9GtNeF04IWEZrUVXrziGBFsIupK7Wxf1Fb/Mvt8AA
cWomz3STnQ9+Dt+T/3Iwz98qmPgQIQQMcKPEiaJMh/EcuO/6UvOIvGO1f5v9mxvb
2Lyxz4uiPm96qMA+4wrCLTSu3NxBJLBRnxRkwTXMKl5KhU3uk+g0b7gjOqRb96B4
gEi9qZ5pixc4juVJFXUH+oI+XJok8aPoQEKXcHGRG2PGlw1ZlKrtCl7F/Dwn6O6w
zqfHbWCncv9QinH9/GcGX7Z2EGtD60QLkU4Psx9w2ljxS9LBqat00RejyNCL0KiJ
e1UBhAbNekktimkuBGQGqinYDNzLmOf6jP6VlVhF5/xAXw2KVxHcvJBAPF2wNwEo
KV0qn3kfHMkcFz+R7J8JKw8tRhRn41JeJ+4uI6kvm/1D666qQQh5REk6y7L4FlfV
//Ux/JG6GKyggZVUoIa1dN3J78ot4CRqkKb/DLk9QUAwDp6JprKoFFNOtLZPO+KL
pbFSZVIQSvSXg+gf8KFdxF0va0frKREbFq1r/IGSngTu1lC1WBg/HesTWAkQVAeR
gDd3v9yEHHHpyv+EtnF3mH6t2JagVCwydDGkv0EDNlRFFp+y8xP4+ElvcYlmdXLA
sK5W6tkNv07fec8Nj2IigthrGV5kEimPDZ+CIZmN4FgwillawDkhQhxqNr4IOu+J
JWvlMBDjinzaZhKcCJFG8M3qX6Na+/le3KT/vT4+Mev/oRpsCBFa/FlnCs5OrTAj
KRyYAS0942EVUTch1M8d9ICu4/f1eK/nFTLI5IKvRC66CnYEI781F90pyr4h1qGY
VVyIwASqw6knMPXnWh/SiNFeelHGE6c8a2FqX8M6VDQgIOyPTq3wWPZRmfhdcGoJ
pdw8jkLNrIxrVFOPkLZ7eJsdF7r4KQDuCK74kQx8qVFYdq55ELHhI/giSdBCtFca
/no7rtmZEDEGblPOINWSWJ2nyD99+PYEg42qH5MvPgd4ZL95fCU2YcQgZR9hO/m4
eU9L1qRahriS1x55ooS0wYwRSxf3kuFOthrj1OdmD0DP1dcU/TJdfUscWmYzOyTe
pu2MVNbX4Lv7xTHvKTstYPsESNEAhFFAfyR0fvlCxJMc7/E9spLbx5HMi8HWOF5f
LJj9N2aXLLoIieIV1JdU2BYqCNw+8DrfS5o0gb8zMm9oIZbvTR3CoYPuh//pevXy
3Xo4WvRC+3CQEklx3W5EdzZH2Ws4qEe4xlW9hM83SXsX5uTvhm5xQwVugAtiecFI
DZB194JYFoGAIw2KZx8BmSuzs3V2glGz/Ow6E6zHiI/Vq3qhmhBr2wt2wyjo3icA
vCghYCuIoZXXS4NU26i6BF5EJxu0QxAG+2gchnXrKBIaZKon5Mucrt/8eFWpHl0W
0lmXYqFt0gSfmsL4Vq6SXVCyNbyy8XL7envjkjwrd9G9zgGaVivhgBxJ47YiGOiN
VRSFldB7KCYNm/wWp2Yg0CH/Mm8vNNL25KEpOfq0LZdGphhSpRAu+vgOGdP0PAwE
xFhoa4OXrLMN+Pj5hX/7HsHudHDKzMcXea7FQcE75wbUoRLosu2UMY/x97QOqKmM
yv3vsueOsiXzDsoDBYD/sjPZpU/CFH0s+dHc4PYTvrNrIybjb30+q/xmU05GUE+7
rpR+mmjI7VWyYEbMVo4P14+SB2QyEw2JYqdGRML6FJvTa+YvoyshoasCz3UknBh2
iHPwpTxrtnufkFribptVslb6+uFvUV4IDVyhesDuZ6KIv3QI9J4392lf3cllzAhZ
Rr4Eco981GGI6EJP40WQopPZnk5JNuhYD/qNNWHcCFzo28yQHmoG2USSbgXkVLcG
xvdtDhgGlG6HqwsSRdHt936/dKSqIU+IMW2xwk0ervtQL6ehREb4pjIM51eLOwwZ
c2CJefAUuxhFZgkuuc/EGyhCdoO7kXxjhRYFx4yWR130rk6rp5/BU08Io42n/fsY
APbsadRqjlxRz/b3ZEMGE9EweO3FBEb9pmpLrNcNuhKjNTGxEN3strInwIBGbZ1x
jm2fcjc9ZbI4EMJvMNFcTytyyMdcNUHPMikshwJ5tqs0TWyyl65R5eZGQeq+m3fN
gMgydI+vcgRJff/8HoF0wsPsDYmhXMWWa9uACsNPsInIybJRlrK7Qhu/xnCI+vBT
b8f59lim0PqcTJzrL0TsosrKQIs4URt+661Qfh35nADdUqNkKf5Xi+YIQYbGJdiS
ph2CrVDeI8geY5PxGt/aRElhWP3XkCpmJ/rrZAUJeEzQ/qHk5Ziak9re7suQiypH
UOwOs1gX0ohCeTczUAMQ6Lc/r2OCK02r7KWDoDURhwRcA9SWAwyDBzz+1DWM9gN+
1VzucnDB6gTEe9WmTsQ5DhvtXRKTSt4uvYGt14HrESGDV32YWh7zlBTusbzr59f6
zT6fl8CSoohfGw/xruE+u8dKUvufD0vp09ztFvgNrVykDqxfJOm1pc0+DS5mKtzv
uVUMR+Zd/UmpxV5fB6msjimpsR+xZ0bEeu6UdM2Wboa4bStpxIgk/gup0OdCpr5/
9Za79vNGYXotbgMYbgrIryn+9+qc6fvhTRu3iepL2SzkdlX+9ceIsG9PZVwbGL0i
Hgjwauso+Scw4k1s252WYcJdOp4jv7PT1phyVVhftLPRVrtnUfZTlZUR0SG6uVD7
L6x+jLpjnm1V4a+UyoCDBItr/0/fnDYyZaz9gckajc2LHpoL3ZgHOICq+dMnWoA0
icN3PtcGf2sXuBL/aLPsLQh4BJQ62jaXtU1lCOj7t1IjWbGN0lGZuAeh9QUQX6va
vz0H8Rf4FWCuEDap2HbPARur/9OWJRzb5inGA4vuXvLQFqdA6yz/103knDuC71Ik
24N8vIxK0yvWjBE5B4RxOiRznIRwU5my5Fr92ZgW0omIJwjl7g03q/6ixn/rLUTZ
NIsMWWU4U1fkmIQXxRt3UOjdWPmaMTtiTk6TryIjDonLEILZ//DgNqgvW7IxjoeZ
mBUeaL0JYv7uYazKA0jxhTp2/BZyYYv9hofCNTrISUhDM6WPw4ofIdo36cWDCkvN
mgwQnJLBGNiGHTPlSNBp/hWD5bcFezolTAwkyncPHN0RIznr8do79fcUW+tvGWNn
wueDEcl1kBE2GW2/3z5QuZrYukc9BwIM550xgZjkRuO6/Es6yXk0elvbUeYCJaFd
WebrUCnG8Mi0wWWcM48yyvqPgbzjj0Pw1X3A44/PMj0J9vBIEtkh8p1gOCqFOiCb
p5SGpGStyLBqH3e9H5im88L2KY9FmwtzedZZZzZGKIxOcNJAiq0QPUC7S3oDjhSE
lm9gpBVbtuA1UQWTI6hhuGXMfmM/KzL7J2ghxqpjswhNaLtVOF20FsATCrPEMb+u
82j4xAyR0ZRYHUoGhv00JmHq5uK8cZ6jsUH/PRMdWuIvCGbt8PVmd8x75rcB5BeA
rvDeQjOB+RHlikuYhbIA1CmhQck5IwNXY6vSZ0Y7Vusp7pxYKsjzRQzj+hACmpz7
MpkexZ6gnbK4lG+fSZoJM00ClJOY3l7zbVf4Lq7OSxwoL5ryNnfs/2YuYLhLI3Sw
5I6RKeC8AYEBuifxohx6TMES8k6yOQaQ4MiTcKPhQxWpjtMwEojbuc8DdvrMLKCy
+Pe5qf0fcYLqgRRmEdqbr3tNpbh4JuT2AZd9AaJVFXsAaE/n9fEGSIn8AnX3MSL/
IwYFa8nqhwnmEpwA+dEEgBAQx4Kz21vCT2KfIhX4V8Wp83NUJK0O40SHtzQ8kuZv
Z9x8wVxLzOvmJAhFN6J1visnI5qnjS66CpR1cHW5GYtcDsMLsMvOVgoHi5sF+w/T
nPz9TlXvhPae3McCXlvfJl+JCWcHWK3z9i5FYak5ZOJEamMSpLFSbauUUM5HVuBt
qFvHfsQ453H96XmYAJ3k1VhWR/dVrWFYoKdyBxhib+iSxJg6FzAD1dNY8BdlXlZ/
Lw4BJFI3zeDwg4tVsLBxP3SG7eKh9/BNZIXxOBowpaUobA2FMjdSyOsw1ADb7Ho7
R+XsHsY1z8hLH3TTV0H3/4/lEr6ea5UbyUUrxvj+GxySN9K8mnE4/TcReq83y0Ys
OS4ALtVb+o40qO19cRXF7/QHABp0pD5RXzUhXX09TThzM8In8WCWOYQ9Vd1IujNP
5olp5znwQwzrajmYUR+Uu2BuT/9Wew1YfstCL20BGTpnFiC0DzvsBAfOgr9ejMlW
SWZWGBR1oxdiiMeTcJd+2hHEVXn2qI8QxoLEJzUgjW7SDTHghNjFfuXJ4VkAGTRt
0VXTb1nW+SSyjNogaj1h1aMHIqjIa5ATiRCbR6csOFnlslxLOZqE0DbKONTgF/SD
2CxJZJ7P2eDEeNaHhaPe76UOgeUSOynRCLsC4XIPQeGagbB3nq85IClIfAIiLzZ+
8auGKNDPR9mtQhvyYQkNE/u9bbIcKIpJnXydXr2tjsiNWG995MrNbvjMpav2R2In
Hd8b1A5R7ztoRC/IRMCCb+qDbaKahx6MQjFvFR567AmkDlie6IBot2A1OY+ADAxB
qCHvnlpBM4WxQGOEm36/198tEkT1VvBgmYKlm21P0FUKLx3692nNDy9DOJ+3pu0I
H3MRiRBBJg5VoyNyMruf3ilyyd8+N9QUswnQ7lR0I8hCYxoWK7ZIcM5PMSWxQPg7
j9gkNQrJzgVLlZ4EKve/131bmXGPjX0am4IGuk3bDyvgzFRLJ27tEfeBPptRlEkd
SrjV6ZPAdt6UZVpMc0KgTd7udFlzoDtAXvHw8U/ojqIsKaUEdabjzc6jTZjyMClS
EByTbomipSHfjfaVsRBps55xl3ZEo26WcdwAYTr2nwKG7o/QLmAlACcVffgcs2pR
WCO8N4aBY/k+shl3MfLYQ4Kw6808drOLVf+TyqHD5J8gmKkxTtQUeqncQNeRWxG4
9hyQFHjqXJHefGpprcFkjaokbYWmn7qtZ3BFEnBUOMZm4r+5AdSowB4b3lRXIiC9
3bVQtLeCb3d46ujG46NOJoLSxKxiEyIrGl/TWaZTrRQRd0JLugI8gS0bA6KCdtB7
Gtrd1dRAstD5pxRc4TrTPrpuveRDSkwBGTTSTSRDxACt7ZbrjPW+xp4IuVoeQ+r1
9jEeM43PAvhNT5QKndwm+xHLwY5ZJknVyvMjsf70lksc5ASJrrsBr2TIReH4NKIP
MOhA+bexUs3qWSjnI1gCy4hkzrah85CQHo37RARas/hU0q/OGWx58lB6Ll3NWmK6
w92R42Qcehp1RBpulRrStC36/tq0HPlyLV5d8TNxR9f1hyeZjM9hKbXeFZKaXCRP
LLBCg03opDtP4oIHsA3VvSSQ1d7jMzQCWDK+9tfN/+TO4FwYj2grQUPGOOM9gN+0
7ZTgHZT2GCTnP2JwoSHjQA2fuDmXjKG80/PeJU7PpkfYjWdHhVKlgFajEVNJoTL5
i8wNtMy+LtEXM5QPs1LhgV6xHAQnOVQZw/gr+zl4ndUF5LGFNX6CgrrQ2MVv61sR
jAX0C1Ol693FM/QbXP1FxALXhVaf9KkTYcyApY7RXOwWIWUl0MoLiYSJ1svg/Z66
CAWkKxQF1AGQOH0L4NiRsEWXrmeoa1rYmROTNikV4K6bvHzOiPuKUfYxgU6sZQbZ
O62g0FA9HKXxN0lAqgdSY0zld4aHBkvMHj5nAQhlWJqqPWGP6IQmCHdu4mz63fSD
TUgF4ia5HO95H+VD8HaBKjG4r0B9owmzN3Z1pJg64iZuOMyIRyq1Vhigvv15bOSR
j8jJXwsAQlghsj6aiskt0JNE3L2KYlg0XLpbE+mYuGOnJ4vLq2dekOcLx0bsM/ZB
EQv3hmFjNa0CgCwleiRAfGz9Nz/F7rnkT/3Tu5pH8hyYGf9eRW57HtR8hXavYwCG
AJBf8lFQZMsIb9jtASiMy0PXwOUbbH25VxTj0IvFwkeZE/Nfiye6E5z2Ag1i8+fZ
fwTxlqtkqGMsFGXH4dYaorNIQx19QOrREY6iqy9LMfK8OiH7n3hopCxhzrY5Dnlz
ysoj8Acbc5t32NaDle4fRjrDq8L2f3VAqYRny2j9Cpzm59ITIEnnhjqWF0m4tNRt
vj3hFbiN2UIhqzgsKs2qZwsO6YIRx/w3RLm2Cr/A+hGY+MtpEaEt4tyW3w4ckRSW
jVXpeMSbL5HqZKyVVxK+6D1E5HuWGdOb9iKf2xmnMzpUj90FdIPsqwlLVa0J+jQW
MHy3YlGzFdv6ENK3s1UC6zdZKCr/aoXSRulNqwj0CgAfixN67Vv9/CIkh7ZPvYwn
MJ0M/cfnyC2dLrx5h6sff5FOZfub0plpFbhm9eBdrfOBddn1AXWRRmaPob1MPRQz
u8+JtZd2pD22jKbtNcnTeFHph+JBnWiuh4A8BcVyNFr7LPDx2gdyakyMuvi//Mz8
32LSoxXDTjpw6qrWIduRGSM7OpegG41VZB0LhG6UnWNYFa43YWT0WQjNSGJQ0LsR
sLAJYm1C2/DhhN7pJXlVwFgupH6Ipmv72uSnqbxBpZ0qxpDG2/GsnBbJHNyvVhHH
Akw4qOkkWtGE4XvC99uBuHFQ7BYBwcbmUnAFiDVM0jfmPbf26rc7zzotdwpnIwh2
LZr6D7hw65P0+l9KQBQPYqINdpDz9H+G3ZufizoqtiTOQezFgmSbN+9yltwalDDc
5eKpVXamJacK55koTRmANIEuXdRxDm9f6LNS9Wj3fJfMSNsUVfHhugw4qHtGiLHB
MiwPUGDEMm+mkP953aQVlGwVtaLaxtsMupM5Rt0+kMBIsIXNbl1pz43qUP6WMxOc
C3w1KOxdi+l9g50Oj4rw2Zx0NgY4HHS9FUWTf2gwGOIwcKi4UT9FeoK3OB71rqjj
RAEwzLDd9NsnRAZQfuJw9NwxPtTNqdexo1oSelRlC0jmFS6cscUTn2BXEolXt3Vr
bNOrMfnUYGmUf8AahxYkYEV4zZXWgE5/R3zwl+bNOGHuYtp5/zxvLjgV/VN5HZbD
lKYOp7t6uY0Sw4BooPm7uZuFwUT7sDVDYJ9hAjLSsteou7nkOb57vzoAUsKDFCmS
piQLrBiYiV+pcE5X8ZqIrXYwkci1XLxR5qfMKOgdzTY4W+R1Gk9Wo+OnnuhSwLTO
X6Gwpm/5RDR+EMJb0w+hq2Mrg1i3bD+noiWAzHVhuekOQ0TYyHl4j3roZusxEOAU
yvOUE7JSA7Ta2bCE8C99FbdzvNg0yDy/Zjbonrw54R8M5CpTGUOIYOk1Sj+Z89zT
knEtpMtADqOaCl/CaHsZlhRp3oYoYsO7nZnDFLMMlgEpHLTcCnaW72H9unrhQgpC
nuHR38P2cbiSvEJ5LCGzqdPcdISF40ltObSBf9F97HEHOCpUS01/fLjrL8BYRxqO
MC9SEn6YBfY1SaEIEXeoQ2wJj093/yZQIk74qEjQumRETJUzCO+3eVsXOgW1NuqZ
FREnBOVVBbnS/wGUJFfuKCH+RlkfOeZYKOcRw/OfGaw0HTOjD42RmcPlOhctsSzM
5O0NzZq1OqQFnqnzUjJLTWS9R7CICTHMV6yH4lipurJqv0JKBu0qOpuPkCEdpZ9f
LgtWr+Jh4jjVaEpu1EUDDBd1Nz2UK5iRKYopFx2ff1IaEXQfOWQTw7aDOi8PN4Ic
DnDj4cRoxoiT8buDrNQvJNYVL1aAJNWsEYhXYAeZzN7M5lmTGBK8co3DXz/3uSen
hiqR0ghShNb+DNT01+hT8w4seBY9gfII2WqPNYzIHjOghjmi8wviXhwgkED39iEx
l2pq4jCdgwDwi75dZvdXrpmyA2Higtr+jnklbHOGzNDYxMkansehHoef9JHuQRqB
UZcp0l0CRxOK+MfN58DJgCUXIVHGYjDl0nJBMR5QAbASCDUJPzU9zbdrSY79bdTg
BLhcSU4F9/wpzpiLGCCQzYaNdIy9VNWGCg97L6shwVYM3yM5ok00a+8gmXZALATu
6+lpdUoBQ7PhSrYUDvN/8DtdFx1yNIJotH4oLJa+tl1MstCzgHmQDP+kEqoS/uQO
pnscuJq0UOHaWGG8g5HahU46jxP+FYQgyaHtdvHSeCRKiZovcz3Y0+0LG0orE8T/
Muls4p/RmCk2MkGLoQJ8Sbwsv4I8WLgIJOxXByZd9g5/eTZlhFJ9fo/w904RRX89
AmHJvbwftFdK9MgASA0otZz28V+qu+BiT98q+/chV5Y1NUH44o1sP/LO+2z9kY2K
91FmKB7+/4HgJn2a1UsudQ+nTyY6sDspnA0yjZm/MgoEIJPo3GGteua+OUMj6Djr
brvNG4gDPKGQZkKbYvTQohMI+BQl3dMOSlgzixslbO4FUR9RH/2kJbvvq+sZd6So
w5rJu8hVIbbhHbxJ5gcR/irhOdHLjGDygYaAjEsE6CMazZV22NaEKaBQev8iGd0g
IHMyuqrOsSZHGnnA1MbEtxP0mk3XkZaHsgrwTz15aqjDUW0Zdv6+lIXdEcdMJo9P
yiaA14NTV+F4PdF0QyfchBAkJwZK3mvGJyNSLsX3pO+/Zq5UEgHb1iFw0uGjMfPA
EryH14idLpMVZ/PoBGWQ363LjdkzS1t7lq/vYD/1jD1K5qWE6Wc78K+c51LMoXjk
v4j6Q+z+WjWJ0lcanejiKeq2WG8+FtNVgHADkYiCBU7T5EVU0Sxw/kBXJTrC1zgo
vDI3061jo8MpuqJYqBvDPdq4BFHArLX0G6YQFFk4nZr6XnjEe5Nx7ByNGp/xeOaN
zbIJ9Wk3a84JCGRQrmQD+YMPw1rfgmmq4xoGuv1/RdvllLEDfFJerG5XAPhnYJ0L
2bTamsEoieby6lsHLLq9Tj5EeSg6KQ5kdrTJ/pmORtG7kTZMMlY+KlqW4YMj7cFi
eFdIqsGqS4Lc619jreeIErKgxtdMIs8eFX72EUyrCrL5CH9lH+TmPs3b761TEXIg
S084kj3HzIGTaF9FnoSwoP/J6nu28z+rKSY9OAYDfxpMBnJa/mQLo0AnRNVsKNn0
nU42UpR7E2T+yMXPqCt8+0/nBiSM5KUKH6vvNU0RhW3yRFNAdiTtbB1huhQI2qCS
sXpgyRSq1I/X2wbCfJpCUQlN9jWh5CvyAhJYDEgyE//P5g1nxxlZo2LszhrZvUfS
qXahhCc04/KskJZWJdGXnArbISXGaNgNNqfu6AmC2JJHbVqQ11U1xjzwizEAovba
qkoIdxjMOGj6XiAZ6lQIWILw9VhO2dfYNITbN6N+fXVzP/EVeVu4tRwcJbw5ZjYh
o0J4rjCeNVdWiZJTZwDNRZcwL0U2Y9wIlnmTxuh3M84aQtGA9Git4Ej9JbZUyRzC
vxQM53Am8FVczud1tm/3d6pBhTLz+YMxKVC3ZNQdxlJ5iGM9hpUXG+FfmbiLQBoo
F7eGG/28hqkLgCZPxTWQIuum99x3qdUA2au/r3PDI8UdayLfQmi58EymEOSNONFt
/M8zXyQLE4WfxM9L1Yjpw5jWSZYv6S+HdKVLjoPcrEmhphjAlKcKxdVJaJkhVHHi
r/YitdIGjusPHKtbqfKZUVl3RG6DlRGRS1c47WqnHmBYn9jPkbTueJJHC6LKsyRs
+Dd7pwwmr0fRt7oxDqkCb3VYu8QVxqVKFCe2C0Rg2TlTRxSfrix4ydh3tpr/SlXo
3ia5Bay5UwvIQDR65oVgV9cEX0SvT/N44MzPbDlHNLib+gRyZBGThmLYpTSM3D4o
B1VC4ROhWt0ez9coXDwCGrFPTsd/K/3iJAz2pW0dkzaAnHFwc6NNpEyxBh6UUujn
37mwNBzsu/Ay/Wj4XeaTg8mrM0LL2JP+cPHqlQPWTXna+O0uzFln3kHmG9IXf9+C
NiJyYpJKbckN4WvxUviFxU+bbzEfYsYhjCKCPcJeP3hLivpM4IDrbqXxFLPBpBxR
/IoopteiZTUC+zEmFbsyQFZdKm09vjwf4rBYFMgDKbi74mOFcahFj1jZ0wTpy1Ps
Slr74Gcqqhu7EarEha63YVQ6c/AhEBO9Hxe3/mGcNVGCqR/3bSPK8tpW2XcyiOJc
MnYpZATWsFxLDabwtbYqpfwcmsoGHWD4a//1YSk4JiKIyuurSaQVHZN5Sf4CHuK/
11SJeKcQNiYkNho/bBeA9S8zgJ0alE0ApYXrfldAqp49aWumlSkKqlD4q26KE52p
FKn+vR0WgETmOMSRXgkTYNxhNIIf7XA+7zxG4DHnUAO3WDoVDO94YbHV2CFM83oe
cpnWOHoH0sjFAc3DqcBYfPz9cLIIEU8RbzkIgV/SostM6pBfXSnkdp1nZDIEZKnG
Jg+gQ6K8ucMqNg88XcH/3iVmSXtB15Pi9YYmP6vFqFbYdA2I8rlJsVDZ16DPUiGp
u+YaHnAlU/FjYlDntgfD8UOnlKDnDVyqAC2BNBJCjHDJxtD3NRbncf9OMxfNJBPO
nFo4wOudWF4RA4O2BWp/1HTq6JsM6SGgSpnWkCwGZufAGGu/hZkj1QInNvqD/RqM
cGAxuYGporN84rmLpr5WCFjaib5/Fv/IgKkGwkh79bVMysFVbCxPpKGCAF1Ar2J1
vfYht6YOPVcroN4Yu5MgB1MgqFQuPvDPL+qwJ7I6xxgH29eI7uIh+I7NbEJPEGOm
9dzm1y/tuH02hFsoSxz4vlWTgXFxB9z/83K/76HyWcwTp7uGnEPqzwvk255MBoid
eufS3BAsYItyb+wTTMrhlhoItSbIRJqqv+Ia4743PcGB8aVwEZ49i9p3srTl9wCV
KFV1Dw4+VrLjAcDELfU1442MfHdvxoNOJdFdgVLSEh9OZ/zcA1agYt8I1HaaedjX
faiu7N5T08pnkZXe6z3wr+UzZywHFHfnV8rQgjQ+oIsMgvr38qczucgCiJRgLYYf
ZLHORZhSQr+Dwya3d1uOpwvHKhI2drGggmMyq+sI6fJvgE3P5Qg6mYBIfJCkkNep
sMTNqggM2SaZdq5kv9KEqnPaUh8HBeSZjl05QW5wnlS5+dfc3zMDsLSRMvhB0rn7
MG+pvirivpajt9WnWqVBsM5X/4KkOZ/kTAwfliByo5eL+YlW1L3US+5bh0SA6AdH
RFja4Uu/LYiogZlvkC5ByRfCLb3fUDcDzm5enLU78rI2ewCK+zkyg5GNG5BUFJ71
jhuWyV541tvq7z01ISCJi7S/nvBYLYxeANJIrgcKPnhSrBLauceVWZn8csY5Cuha
j7wtUJX2jioxAjrrdOFwfoTls1PXHc9EreAmx1/8mrjTu9XqjkjNXUZ2gLTqRW2B
y+isvzTs78CtdiiHUTWkd5JcH8n+o5/HZk0I6UVguQ6z8PaCQlUbtd7KPrO2ynrg
pUzJbsQQH2ksc0KZS+OudrvSohWU/12t09vbvAHrcI5vrqmlcPvfcN1CaI987oOb
glRJWuXqEvhJ2jFWzAQXzIW0sFJxqAd23EmHg37rtaZ9nLKMKuU/wecw66lydcCo
jlsbymEV81mB5UAx/fC/AC74v2ljGu2GF2p9nM9axNXhm8RneNZDVzOcKVVeFoAO
dx/wDYbayhVdC3t3+86WrZQhmN1SPQ8utlccafliXsHjjBj2LgPKvUWHhu2J7ZJ3
ZQXOOA+yllOJZMNvVL9l7fpG1LQIyhNaRe+t2vfnDJWGM8YpmSddLW7bs33Ogt1y
VhumE8e4flMo3xtYpaJj5ABehNe3AIJ2TPUL0nvgPtH9mdGeuSITczYfX+vaj2n1
p+MYFEFrwnthmhrvLxSUSCzl7xWPXXmbWnKoJZ8kl+hqT/5yT7fnDldy9hlITK9O
mWHByNrnPxC/tIXyw4oQ0fzXOkuwLMS/BrPTYIk/XgU8243DERCyE17+hlMBmur3
UyohzzaGtVO4p3X6R0MU2YucczieVvhUpm8AOyrZwHxH3TPEQrJgYKyQt6pKKUiO
/GfsNj8qeo7Aa0sxAd4xC3udIinfP4Q7Ad5YolMpWkxlhCfLnfKKLh51DuUYcWMZ
zBK/TayfreEtU2EnL8dv761FwH3sz0IAu2PF+gLIfZU5GxHC7JOCt7l5/JAMTVPO
EgAGWb186w3HBnmSTfoF4GrrXVZFSkTJ+XDTePoudatVK1XqYkIuR/KX4Rp+fMVg
PHymZMN4Eogy63Tve99nhYjlOTbkoBita05vdRjfjHzjh2qxrGNG/Z3IC6ey8Mre
OmlaoNOmvON4vIho3+nKe4tdw55H3DY60yEZpxpccbMq2FAFVo+7YDpK0tosrtoR
uDvgVgW+9lRG/inPDyyoQjupuWV/PmqFwxaoIP0DMXTaaY4cB3azsmv79zI/26av
GXd8Toc343WLLj83JCE4sqfi7KT9/X2MLr6zLzNgnXyF/KY7zvD5nu3r5suV/dZw
bJB73Ed4s/b73ETWukeN9nLJROUDKm1d1et3dUfaWMIohj6M2zChFM22HJ3Nx4p9
1sdk5H4wmvdMeDvbBW+O7u5/AvZOXUWifwPyQDG0H8eaoTOYZde9qzzgJpnKL2NY
w0S9jmXWIW9WSUte7ttUuVidWMPjvPeF8seRCVW+eFGEKziWjQNqzkH2Wes0U4sl
Be8GeJCN3nGgiOckxmMRx7Tt3kwarYbv+DiDemSygVW9nWd6MNYG5uKJMTkgk/ev
vXWCr30j2cFphqvgx/h8VFL4Vyas6+nVEi+zqLN+fFO8pqzBYFA/lEWapZCq638T
QnqIplLUXb7EUc3o/TqEpnHDrPlC2X4bjZel7vbk8ZmIpwXqgSehoOC4oqrEPPET
fB0IZtngp2t1/6UWAZqnCXBFfUmcUhm4pNo8YjcuJ03JBUUz2cUhlqjq5/oOLM/h
/MicI4UTifOJuCZxcWze3ufJb/RqVTbDqfT26aDuMVQZibCoNzs+AdwfHEzo/wMC
ZfHjhhoingbLRjjnhbyezEdP4Cph99cQR6oqCYQpH4lEVvjdcJLThXHdXqEnwGjP
VznDWVYiA6BnhFN3uuwndOkOwfQ5b4RSUAC4YYQKyMKXx4LY+7Ln//ly/+AIJSHY
GpLUoct1YZEgfWqctXOiwJhF13JVlKbzV9SUOiUA6OKQ8IlcdIgUdNizS16tJBkP
Vd1pfH2wTAe/9rzJblFMmL7JNHVRnw+gd40iUo/iD5aDicFELHC1EykiSh+0eBRr
Ux8BvLtg7jJ3WSB7iKso6LBTKlmo4DlCuFZKH6IbH2PG4grOfseT/AYsXkTgOx0y
uWjjZYiZ8pQtvdzbUb4gBnIRD5BttEFRDLx61GlV2tM2eDFWxge1kYQ65TgzjgA+
lUcPCVH2PPswfJqWyXUKzIZLU24d5vbbBkAMbOIJQwPImMELLe1hjzZiRDdCO7D/
8c+R6mjTigLC46BrWXdr8eVTNxLSdfQ/wAcYMsDz8MPE/AN/nzEBpYbbRrxM71tU
/XapSDdU6JCWEXQ87732JY4ljtG7Bh08yMxGF6rOsp1umOdpcMokxrrlkL+m1EMz
29v4U7o1EEX5lXjhe0lpTK5/NKi6ErapC+WLshlIfVPNGQbwJA/cAEAb+oFJjVm2
JlIhw89NhuMcgxd0EDa0nEiKbYr1YTsZlIpMnZpf3D9r2bSZgL4STnlpTmANhFzz
uwR9mz84TlLgYUeqEDGz6QxvkbA9X1DsS14y6cX4BKrGqZrkUxhfO0Sufv2niK8E
Y4p8CC4MHcMjcLH2ec6gTzHvJdqdHBV5jm0LKsteFAXYaSD1UpMpUvEDIF0P/Qz6
sOgBi9JldYHVmI/ZSv7nW4vGDBDisreLDF6PXGQ/y0tWC7NOSHQm/g26DSS16Llh
aYG1CH8Td9CIftjWECkA/VvIOl0lY+D0f9VtsiYXXe1ILFIqKC+upgcX9sAZMNGp
m+JjiHUvkqbXv2jfVjkNdWrSpqHrgEboETmDSZrfov8cdiFIpyzbiCl75g+12bQh
iEPlAzYvLhIh7VWAbd9SDwoX4S2PbO3ALW6y/YUffwgzI7ZGqMFw4yo+53EQsFB5
vFpbyBDtNTkK4Heo98dCnXDa+mvidWonslYEe1aDwRe4qmIf5jApzSJWl33Gcke3
X2i0dEbVSltBt2Y+7Rgc4OX20N2ZGrN5tfRiUcT7aRLFKxqjBltK8EI6dmoa7MvC
sHuAuqrEkhXwqZT6kB3N3OBFf9BnC4uTOAjLCnQ5t4y3js7hP5j1ogffRm+okYyM
W6D5hg5tM8gfGkeCQ54k043nzhjINqPrek5EEpGyh462taZFBuEQyqKNre6AU7Lo
z5QCY+qLvbNlvVtzA44YMPPIt/bHwsv4xBo1dgTBMNzh00SkS2loZCFyZA/+qdCH
gf9rA3QCfHNARYDGdolYinGZD47TNFlUZNSvXafMKaiX/gsgbaviK2Qlk6vpALLU
ewvqJOIpQ4Z/h73wO0GzSosXtE2Y/5oBHUjmxaFjkaLhex2dRHEcb9+UNquhEgLL
IvX0YJcTyOJ30g4MpY/2uFOXfmrjRrxqLpaEb+00oyVjrByDn6/GxLq3RDgr0h03
oQLxIkS23zUOAuXcWp9oVHrr89YVh007E3yQgqEzUmALtDG6jCOFFmY4wumrlQgE
NKAsOCl2u7X9kKY3VuGhrW5+WoEXf4l7cqNhh1MH6h/DbGRhDDOsRvDfD2/3Y1w7
KnxpEwqGsVNT7lVRkSftJxCt7YghpS089lHE+Ql4wDoGFV3IHHvGk6S2QZlHNDmf
ddhRM1I4T1W9fqLIeC4RWEziuyKu8t09+PCkmTC6CcVNT32z461PqB7pLTk6vOic
jTYC+2lC5jQudBkqlutvufOWEzI0wTmSvtIoTsz4i0mmT5l4mwdM0m+rn7E+TGpm
2vy+hzF9S0VRPLd3jw4UDpwE/YZ9JHq+Y+c8qZpu4VPyNJEBVx/h5H7ySOLnGAAN
Jc0/CVl1cqeAfHCR3gsV/b+BhMZrNelUWktTmWhwjbhV+gF5joulki0USD6F7tiR
sbXwnuJB64qktzi/okAJ2y6NvSKBaugqvkAdMdyS1b25DU5ZZmhNDfCU2s8PRQwc
yzJoCJKDqRtydkzlMUKS81Wx9Z1ppsq6nhrmDC/iYit9MyTGsazbk5rAaOH1jy2J
Yn3qSVYnr/96qrwZ5mgM9zV8rgZGiE8gNbAl/kW7iqeIws4BuFNIx+3LUXs0kBUQ
RNa7MndIGG8X2WW2SOhY96s+DID/Bmc2y8qVSA8EADI5SJX3DTuPP/A0q8W+mnIc
a5vHWmZGqswwh99mWJO/WrRS2C0Jx0RQB7Whb2bq/pGUgu0lWj2PnO7sJXvkEX4e
nn0bHXLbpA8qxaSfAtyCBV6K4r1XJa/X1T0tliWcx7XGeZYGAmhGVkm+atwP6uDP
APxQi1VDyYuZkHj9atJAWTPyIWFyatKCeR+LXw9T5n0DBFTsvIVsHWZu53wFSeGY
MMRh8XoU3a1SuFZTy42ew0lREaisOWSKiex+GaXnXlciw5/Uz+CzTmqys4rGXvDX
KVNKsEpJze/GAYEjX3laxOpDO+dphCK42aTE0Qi/8qvtWMwdt4hj7xoALXdeqFHq
cMlxGsfaLkGydV9vHAUli7x6mRgjJIA96Y35ZmuvS2fvWvIX8V4l5i8UPfexZ8o9
xjaHNBROabkip5Hw9AvcKOXoH0lu1zNx14j8Wkd6OfOgJCh/27TYjxWZEW6fFi1q
e0MOfH975ggu2FYtrj3tg7kDen2zC9om3F2RJWbRLRI+1qDYNPBEz9IWVa+xmqNI
ZOmjE0G7axEXM9ppFtNWvY5GJpxqp8q4aZn13F9/tnzuUlazNiwNxK3cIX/uOCpX
UJSv6FqCLU7/hQIgRtnLDoGD1VoaUBHOngU+M/NHRwkMqtLSS/qkgX2EAR0891DB
kl640M9tzNXhkFSIZRz5b7jnty+qqhHvHH/LyYs4xlx/HRW1RJ+hbf9xPmJ4o20s
xbpz9RtVoi9ACxGsmpFWmI3S66gg8cEHFDtiLWKFNSIUfq+Iz46BVjc0BbWtAmNq
tveumFF5GVfhNYeslcsZ4MZsrpyKmjllfUHfwAwhGNQQFWtploECi2+STAX0C9Ou
VbNwZvcSjesFA73iC4bNZBck/83oxOlMIuFfjVERDMBd2FgvBT3Pq7EfsgCi5L2f
SjcBAU/BybYewvdrbkdRVh4hZNCp/ey3Q21MPiKxHU32oIBEy+ZbVSxpHkr4pBdL
z2IE3al6bu/Ru3C58BP0DSbklcFDMLl7CiRzQ3ZpHW8TXYkxB+o4jR2qhoITmC/8
Guq2YZRNu+vzIo/Kbfq9w0oTzfR6hsjRHnL8CcLMGFXJmnQTvg2JHfMWtavKTmVZ
v0VnIruz8z8+QIquob6fAEbnCMKP+bWHvKyvwZD3znsY7dRHEtL/QXgrDTGlxypT
6EWrk6/wkH4Z02GJDJt4Uo6jwY9EGh0nYhGEo2D2fwnESLFgjPp52/UotcieCg2X
+ua1XCvAI411wLXwwAs5+eBeq64Ctoavji9OcrW4EbOPbtQwx5ovEsZqPLqdN6o0
gZbNgvd0K0htBvNAFodfsVXkCCRkNR9C6UoVY8Keftq6q35yawhxNkwOjE+0zzB9
H8bBFn52JXd+ydiEpkYSNxa/Zg1ok3m04ijnnYHkhpP/tPQxl5b3CGM91WQKsa4P
5B6Aka/9SiQlaT63ppj6YuABMob8CSixh5txJFCkSZNShj9HBsCtb89HYR5ILd9v
7kX3x6xpqxtYGDGtyXRgPclnOmtEdAT6S4tXYBqFDkyRQKZOLI1HshIBD5O10Yqh
QjA+OvDpqhllQp2J3o4QOfbVGvFmvTRsOJ1lUI9bq+bM/V5Y6rMifmdlHX7Ar6Nh
nWbZv2cXgc/6ga5Is/a02fOaK0nOHKHvIv1oFK2GdNxy4iY3SczJS9H8GPtmE6v/
VeNBzr/Z8tr4mkFYXY33/BUi+k1UhWNwC8F+p9n9xoQNmcqxpT89uEdCNQk/mww6
MMBVhl/WchzX6cjVv3VreHBUh95+VgorQqIEI2+ZaEWfMmY4SrGdyyoZfxxNe2Eo
9RWfD0N74i4cGXPem9kYkHNk7FCBnu+clF9i1M54ANfMK1RkobZ0qsy3ByIXy9/1
CcsTlsRPq9r2IxBGdRdUduCd6Hx0UwKyDEUfwlx3aO6Y/RuG33R7vA+VH7UxHMg/
b2TXsxiwvemKsoU9CZiICrcL5DreQP841JB42IMYeENqOv3O6yf9RB2jp3XK5g/M
gdVyaXPY2NAxtZ0n5GSQvFwYQRoOq7HFOEODQvlb+oMG0sre3vyu+5pE17tOGXC5
iank1Y63hwU9MWSspkvi/+zLl1qdxVU2H1zBxMTipnsfBkXDUHFYWjYXDMOTSY3N
jXdQ9wpMejMEPTiuw61NjJS0R/0Y5ntBET6den8NOMyp7uyX5QKmmjhCIJUUxogy
K5K3x+oEGMVITicGaRE2iZD7FWmySvMCqmSn68ZTpfbyxJWgBsM0XPKxpZU1mOmG
QdO2hhcfukfEuJqj6U5Rc7rTCFGS2CM6fwine+G6lbYw8Jb3oODov4kepFq4c9ex
N6BNLjsFT5AidqPpP3pvTYgRuk15HTA9sPGLAhDalzHsepPRuGg6/Q5eMa4MbAYz
MvJH16uzyJnGRMzrAACG/KA/ccdI4aR9Q6SZivlweC2gFyzR2zDoRsyMBJYICaeH
MIEGoOp03/BTivafoMA0yW267fXSZGdJ6EqFChxaU3yTqk3mFt1yHHM+KkxYA4VM
rcd9rHCf4p3wYoijvBGGOhXRHtDMssUIZr9WtVOl/WPA5dFdbOj4uv5RhRUSuR0F
LiJ6RtM9VxvSDxw6TIA+w6tiIdnEkbXWgK0JaRHXT7xUwrKKwRQ8S+glJHTW6k6H
wOFCSTfyEf3hMExoXoP6YnG/2yGL7wlliZ4Af/FSmmwdwBZw7sCFmXtVIlE8IQPD
o8M/YMG1q7koevAH1BVDT1cDl9ckN/Q5LS9T5n8iVS9XQwUSMDXMbOfoDrUS6cGs
6gf6BWcR7t+MF9tGLH1/oufhjQeymB+8xuVLD4lerkxlIGn1cpE4ckJibIqViGb8
jVYKGZc/Ym04SC2ee7ha4oXP2qwbUoSpNdbEP9W84DXqX0XjvWso6GMqeO2IeyTA
v7XsDD1npSEIKtf3W4qS0yn8UE02aPLV5qE9dXVhhrnLtBwLVUF8dxsw/jdxWEe/
Z5No5RuxYP4JOxHVA1M7fXDbLuJz0dHpgF/dlU8c8ObB/+pH9Qbh5VFQ2qJyVM0G
NZ5Nei1N2ccYeB3NUT9wV+H44sCOaih04aA91No0jCoBOc0D/IFyNtvqaIpvYBhc
hvbck8Tg1dCHncAohPqGyNkKJa/Kf6d+K5O4YnFCKib4yn5xGSQnfKKakertBdyn
t0GC7L6MnoiNT30rrDtBkfPVPY4vqyFSmaByF2d3c9JZOG7NVXE1fF3/0fa65mgC
yofzLnFaYTgkXkRjzAetv+uaG5DQb4lSc37ntaX3L+iaYXpmSVygAc9gADyKFtdx
Cs53M5EOQsec44gzwPuMFPh3MgDfA0xcrpcZi+MeDRanA5Z5JPtV5x1Ozkne1QIW
VOu7d58Yum727l+m2si9xYdWMx0Fahup1Qo0BSBsWt5LzlYP/+R0BC2tPO9xnslm
TiwNQyzWgKMTSr4MtCBjHOGX5wv9PBUrlL7/K1Q7PgX34FK4w5kdoaBqHQuQu9LU
prHBQOlx6GzEjeDeJtpVFprK6Cs07OUY1qlj8k4thGsm3yIJvsvoiZNahhPaDDaa
vmcQE4tRAD+C5YOFsdpolWbW9On3b+90RZbejmxi/B/0hue0vAB14y4Fy8/YW0Bk
Wb6gKGjhXvciHa+ae/ODG3NKfQarQ88WQBXfgsjuDq72yFae2MrPNTdZ0bKFRWwt
eAB4mUi9Vpf4mWPtoBDWO6dPR4fGqzek3eERBO2efSuazl3dNSTLOB+DYI79JgXi
40lCXkwtAjZXJpElI4PenPuB8ZREQiacmlfjQt0IkgLhVbYyE8VsGgSvW1n+ZckL
RT5dyRHV6JaaJGOmFssUAgzrIj+XcdWigZSw9J6albNAgUr+G+2zS/g7WhLBhd6v
G1WG+WzlmCTyRxf9aNt+lKHZS0D2h3O4+YgY2zBQX+o4OXhdq5vnZwHQe+PWJXoh
cOpYhCg9RvXN/vcsw3VOtYdfSeJ8F7a8z9o1rWhJhlspz8cCoak6Tn2ZQIrEb6a9
os7Z1tgY6MNl9syCFLkyf4WyQHi/5CTBnJEzDCdL8AV2KmavA46XLs9SFmcF+rFs
eX0uA1rfcSmdStvtNb0agFQxiGGj1FPHtEy1soyzKBLkpgFmRSOeFW4VkGu0BzU9
qovauQFkV9zxxveY3z0vTtFsdjwISBa4BvoMCRBE0N4cCsBeizhotQAfVjAfjbZz
pcg7/SXhlYufh07M9cJPmKjYJADDHRfujVKapDkJ3+ggzf3g+i2zVIVNPFI05Xhf
FxW/HSDHeHplRsqRoP8nvc05M46B8Gm+TzIF/6Pyv61ZeDkpYTOYNmDcbS5Wg5Fd
k2OkjRBb7GuhMpugtFtF42a1OcE+/BVUFo1UmqG/fmXtLPykqcVu6I7ELGlrpLNI
hloE37doKUsxRBUczpt8l1w6rgQMii/qfdjmYkyguIMllp66Q8JvDpPL1n0qjVnC
CFmafihR/RsvmXmpQeJS110MN4my91hgAl258E9RjLCUcWO+t5MYKHBfpLQgd8mx
NAMftN0tekgHkWGBov2Riqj5LV3htNOVP0jHqHxufFskYwCrj4rZtbjpMUGSKgje
6DaIPjVajxOM1MOL5Af85y99gE7u3qJrS5jneSj1N2IYylrAZa0nCda36NLMgVN2
ghMJHf+X6sRYMqM6abp+tfk9ODd1IC5T181CFuNOPG5OcCIGXe4JdFyyrwIzHXhf
xITqxA0VZm/J/+eoknzAT3aLcuZmvoUhaudjYGWh6N5HLaVvcz/9faO8nF4PHSD7
pr9E7UzP9ke/zjzbfEf2HSeAgoB3DQM3YxdqMbFiOUKS9sRs3BaKSn0/dxs0lUjD
ss2z7CNZHDW940TuzztzWqAEzQ0clCd2aC2x60FodmZbLihOKEZshWR3H7peIspv
v8OO7cJxc0adLrtDgzf2pSJ5lLcMlt5AkGeh+lPdFR49aezXVg+ZbFvRExzuMg9b
O77xGDz+dMIHf46jnzZ6uN7f8K8roYwh4W/QpBRpOKEg1ig3L52c5p2KsAm/KBB2
JR4MTLV6J5e5+Vi25OfmwQ1HCIdiBVilgtRIWjEmWRO2bkZYa86uUa8+vSmjDj/v
XBmLMpPDMGLO+fjLsB0U+zR7jjZFSKAC5l68w+EjrVheJsmvCB2XrS+ReurErrUH
HSQGuBLb19FfWsg4tWYvwElbmuLp/DPwLSn3C+BEiDIDHC0PuxsLizr+YZ6XvtM+
VD392k6pSiZq4aDeJiBzU8+B48998hmCWESF+eVelFVRYHtu+QRdfz5uiDai7R48
EpON1iykD1NXMzH1DiEqrCF1Cm9jcL4V59zkXBO5M0XrijD9I21/YREgkyaaQeh0
E3QgH6OKI25n0hnzIiy8YIa7NZdkj2jGqO+bwJQbJOt8hteB4Lck/XqpG5xFWV2U
5i+heZ9wpohwffYi3FdGYULtOT5jRkqOE+ZfDb1SJdPKh5f1HxgoKduvQZ/s1x8t
pxoq7+e9V5HNB2rnADt9b2cbueC/vpaW/xiJNRlrTyVMkbr4aZeD12JxaWWCCg+H
c5DeD/T1xFWqkyHnX/OSegTjciR9pU44y02mkCOBZ+DuqFYJ4HDjwqbhCNMF+xwB
AuLTWMfps1/gw7Q/Y+62/YkjrK0UpD3M6LN66cEa/y4Bpi9uHNJ08A9eo0jS2NkB
SfPJI9utnz1zSzFhXlF91HoOzDoW4cTDh9BL0M0eO5rjxaJ38LL/Ew4/Z+9dcyAq
ahCSW6HrwAGx8Qc4NSaOv+kWzoCVKbOfLJW8FbwM/MTtdB2PTGVTMP9meRF5BkHx
ecoE05WI27oI0rlpEdSzGtHkvZsdJIsqs18VvEhkkTGA53hx9P1cbnKfqsdCUOyr
y9MdOWOxbleExBTjewHtDPsMVt22QVZfnYMrKFXqWKTqO7J8pB/ApGr/U1MWPcsz
SQyLYZhBRT1T1kAuEXRU7y09j175GfcsiuA0n8D+2RcHPKIekVlmOjX9AH5zycIb
6mgOY3En28jVoRzsgHHP+xEE3hi/HJilL9eZJd6zJwSf67b35GrJBvx1eT/ZiZKK
n0dxWGsJwkM763cU46KVBMsizn9MWQp48HKIyNXBAxxjlejwl/EJfteoN3OqqqL4
GSQa3S8Et1HziBd1upH9izN3lrbeGHwSDlIWS59nLbyh4/nUNUqc12eohO//kxiO
MU3tjuLsuucmqddg0lWrvQuLEHQo/26QTWETAbHm0ocF5BC3GjH5tEKPOwjgHpaT
YCp95lMPIhHYMoKbyUZgqYv+zzR1KCPz9Z97EHDP72v9VsPyDxov3C7URD2D8yCj
N09So+rU21LIhslbRdNr4c8zSxShRggAHN/qgS0BP2av3EYRL41AXUumzqfeAHaP
KJNuoGBZewM1JX0LcSYXM+bldBUIDnt4X5EK9zG1VvjMienlcd/qm4NI2jLFFl65
70U8UFZVrnHEfe1TCXCuvB2v+i6N8AVspPZ1ngJarfBPhufu+PVGw+CgAO6YVwo6
v2YJCEtUjb1/EuHXA4K8XIaAyXFl8o0cQtzoe3XI1fHJXA1d98mh1VuCb7tdod4h
WZEoVsaRkkzbdSGrrQEdLSVTDDaArZloAI4JOAFyva4TIDHNkkQvfuFRzHdK2oMv
nG+BHo1xxz3i/0aqQlJayJZaYWu12WPSR26lEg1D9UIaN2OXscqL/UGwj/3sALJd
3As5s3KW176y/o0kiIjmS3Pug1DYWSuFo4xykCr0BOBQuJcY9OKuYwzGWbA2f69R
wlZqKvhiqgaCeRPVcmoMobz7/gYkcXH4QT15ReohNiinMrABsbjhwL7Vr+2ZK8l6
t6UmRq5m5J6s5lP/w4bMwGiic9kLwDlQV7N06Ak6Pl2O3lB3Kz4N7qOmIMrn9lSD
rH2uy4WRlQnRenCx9lYBnvWPKKQqOzcwByvz+SAOyfSoOGICbpcwBRgkzh2xPqUF
SYaimqABmuNGPkMxs+CnKVVDOyfHOowua/kLOf86CK0q1b4EhLKNhr1hmyyOtrb2
qDvijjh4veeSKjIPSbNUF350eyKhptoOHG1b7uMJm12SrhZ9AT0Qadu2Rn5J1/IP
inxRXbkIJwuISidkkfcj+kF9CloPGs0XPaYyXQlzsaObu+BjrpeevqovW21GYu2+
dmrakZ7N0yM9300aWAgLCE25SYz7JRnMErfvG5ed7HHfl4RrDeuhNBJj31Hyr4zG
ON3YkXM1wa3P6YnFS6bmTPTXH9X6C6PjL1i2GXb1NahRnRgzA+PptHZ5DZVxo8V3
vkwVSp2I5kQR3/dAb6StI8gNVOtfInbfJsfjKtOu+mJOs6nTfiuGqB+r31JH2Abl
GWDx2F8xsYZFu0eyjMOZzbJwBwHpsi4i+wliyUEVqpJp6OSAIicXYR3uDUVGQDMO
vcVMO6PTp31Ydls7mr03bynhU9tPguQoHWPHzzMmfXbpNCEDj9c7BjUIzsgvGFde
lrWFtW1hyZy4RskW+Gk8Gmj6NCeBLDG9s8E1/r7grc2XKtmgZPM9daG91XPseyuM
3x3sCzGl9WPbdMbj+quxGY4L0WQ631tjpb/oc1ux/Ei9RdIHZ0kRdBgT+KxNpM3E
yAbgHfADo7piNP5HCNLRgAbS2tx7VIwBta0M7txzRQHNl5W8HisBdBdFuYnvRFWO
r0+ZvBlKetxMFAAMcz5kar3vUAcQfNc7+lrOHyd5KFGNtwusb96Iq7IwJWQqD4Sm
9XOkNR3+zP4W8gQ7tD8RPi7Esmc5qlyZqL5Rs+hvRGvSUOIYmjSAmOso/8RdnJSx
GVQhOdW7odsODJKZS+kSXnfb8DBEvD9UFrxeQA9xVh9Tu4k2ZWR3/ufBNKnNP67t
fp579oGrDNHvlX8MJumT5/gDTTr6rsr0Kqk39frFII691gxO9pyZiP+5FjsJMtql
xb47sd1sZ0nl7QXYtSsGG6ls+bI1Ezj5RMwnbdS2Bg1UILrgIpUU+g1Hl4mlgrjR
IpqfCMUA74IuRJWQiTDZTrKgK9BA5ryE/xoA+DsSjjPGfBOZ+iU7dkEHzrnNmLFe
RRYnyFbRmfdmcmjnsk5H0FcMhA2pwMFysosH9VmJW5pGYu6Sj8CU/+UWQ9cBXxoc
MP5NHyJF956IHwjtptuBRTvAXM4mBCQ+Aoo30kAOHvezaMa/nEks5lfMbLYhGysN
euCax2ErPuBnN3qOV2zBZuoLIvwh39mK+NeWLMdijp+28Iapzrc8nonavgtNd7Iu
F/lfyBOwk9mGjYwZjLWKfSfwsS92zNpF1c1BpjVoqQ950uUJk/997ctoLtoezoir
/hzHUP5ZNm5/dOER7s/YZFcXJZrFcil5sv4Cfnok4CvyO0qt8yOGcWGF2KowXuk9
aIWwgBU+gUA4SrB+Ei0Hd9fE+ceehH+YIRO7oQcMz7Lx5JtQ6jvSVh05hpt+msQJ
Mpgbp+WuljacSNsv8RoBXb0MxNLaoQfVI0EImWkbJo09wkYQ8rqCzkPyBLS9zZhT
N04M1A4CX+hHeXv0iy4aronxd0tLQOq1S1sEjhfloWhsIg9xA8eLz4HGpmO0QL6p
z53yMiU+sm4dk0YA4jrkAFOql+5Ejzl6uQc0SQ5h1VRbd0Vxsiatw6AvmyoHIw93
/BauouU1BcCV/SlRFS4dstEj6vGzR2PTijlqQO2dMW+7edYGXEB7pZSiZ5RsiJb2
tzGKFh1Sgk6ee2ytcm4hVrhOVgCu7hssujc7rbEg8j/sq9ZodYPvrf4Iq41bQLcJ
mnIcktO9GCCkXhFCTpHFxfLscdAOURKglv2zMg5ANNqxAQK5aXII5Z71r7ewov57
jSWBzrDsAIrhmFgH8+62gqXDph4eQ3L8Rk8oSb51/CdzAan9D47J1YnqQBI0Zroo
vsP1sr3tzdKSNBgCqWAwYc7yO+jdIs4eezn4Z9OIwUStqobXMOxJW60RxOzf7ksF
+8j33z4nIlwFa02JtSv/NAj6RwcfpUFhnSAmn9H7OIUhDp2/MkV0KWDzUchtEf9T
sTmLHWtPgg+IBO9eRM9pNWzQ0vAP8ny5HFBIdc5J5tmXO0ofaEWDGW1/4CBcmx1d
mxjrEpgYvJtLcwViRgIgzP3voCcAL0THfd1JMm0id1qfyzT9LBj3cxq4E6FEiM4i
iJnsdbApqDlmC+7Dph711azitTb2l84ZTa1sClvJ1MCQBGHDNGXKvd89fGlgeIzC
IZUTp87h6ww8Bv2qBPSXCh0veUjxwfSkUE78KXmAsdwbZ1aV9xBJ3cU/BcyqkdtS
CCMdZ8tRJiLkrbcM71Jwu5ryDFcNePdhbod7OugfU1FKg8S7Kx8I1aNDJdtJe6jT
3Po6lN3G6BvdN1x9nFi7c12TyTCJwZVB3NOiHen9FsoLaSYFFCBkC51ghugQs6tu
/eH1FrJ4Z5Rpw4PypeMKLyRpOw6jDEtfEbADcD5KLI+dVyCMkllcP7odw5J2wxuk
Atp+khPyyeprs7bhltr7KalI8j/+i/DeAZ8qlGBZSVeeh7ClEHqd9+2jmKr9NaVo
DvnBiQBRgKaRMsOXDxm2Js0itP9M3RF7iEXcYKAP3xJiq40VYYYE4wF7PXbeUiE+
ySBYt82nD4zvvDXB0lr2IuU6oDtrK0VahBUWEQrlVESIbfdc+EVNpIku+4ZFUm0i
mbgTO6zOa1/kPR1UPIp/WOpYo0/0bK0eoxNuX41BBD+GU+saipXcy1EyV0eZW1MC
pKEmYyt+ahkZ3WxSpCXFjxSFwBMN5lUJUr4Xtzq32pOKiZAc3VAPgfeeGKAvfQMg
9/E43VXpaGmGlf3w9EqP5a3+gqZSP2fhxIw0cA7/Vdy1+DYWTRTFlgOJHHieNZQz
aqSOj/hyzVE8pIHuBNd19NcKnr1Ic4TGfFUnRF7rZeXpXkrb8BaTBlvnX2Z5W8iV
dzm06Dq+gti2BrA/qWFQG6MqKQiLHYw6AvoQ2UowwdxikyU6Dl1POp1Z58jqS12Z
hz6JFZAWgA0FrnE+sFJ7W+notrUf8HSwdV0rMWZthp3pyrOrkMl94ZzH8ti87JBB
Gk9nJGRjGpTic6sbDvDaR4FMitdERqdSvuueuETjWoKllxChSrAmf88RK0y+oWAl
WrXiqEBQnZoeRUSyDYq9D5rlzS5ZxMJc0y3IlRxgbP+HYs5X5f75VpxM+xbWo6nm
azRJJJbzdzEo3IkaiM025oPwI850iicN9s8qMrC6x1fG7CDC7V+yrk7wH/RdHCby
2jSmm1Wv8qkRx3vbqKorDz8nOUg4DSvEpzQq/oWkg9oumMWy1n9++jCS1Wl7Dv8J
775ofh/uSG6/KodGqe7ordr04CX0RXsjyPN5nqrI86P1Pc1m+h2ic+4RB9Nh9W7j
UpA+aPRcdAeFwNIqrnYJsUv0fNPF60WPfqXfSzQEPJYE3lE6lq+sluOWqnYi8sbM
BqwOCaIlQkm2qwe/AbB3XmHMThpYv4h9hz1+Hy53mYYt+2jNn7FS4FcfSyfG7//o
qDfRWTtXopAgubabiq8koWkBVo6+QBiuEValVsgLNQ5QIEKN+qFzSCi+d1g8LvrZ
62Y2g52BF3PsqSGT/Wo0ZSziambv1N6VJg8+3qjq7R4hugR8zkwhBhexWrml7tcw
yyIePoR7jaAW9jzJRDi2Bq5aoG/RgC9JabWL0Wq83tnyppGaHquCr/C02uelL5wQ
zqFyx9aJDruiT7sQLgN/04HCz/irpMmV/0bCIdLnZT95wuyrPOdcfM9CVx8S7yYH
F7rNwNMX14pYR6ROfmCrc/5O3Q8HYbz8aPN06BVZnDi79gh56/mb5pPzIV5D+XK0
zost+FWUA5eVsgpoH7l+mGTxAj9seuuobfE9cRhL1ueG9gee3Rzfb53KVpXEu/yZ
7N9PtrpzULpWF9FBBbzl56hwoiwIYJ3RztHINOAwKYalpjw5yYZnt7gG8o76EZ/3
GltjGZ4SRrkXSXqhrGHIdACXUxpCwpku4U+1s1jzoaPJx1XAQB0DlkvfRZU7PxNt
F32l/mmti9Vhr+BWnDzNI7uXUM5Do1MAsRVt8oPliK8IlxoGgdqrcafxZbJiECp6
UuYIzjm47XSGKFtPZrtzjJ72CTqS9fvlZhjnV9bA3ynQCtcDqvsUYTTqwgAzdFI8
ZxTJwK7hsR6AVUaS7CUA+ha0Q8TqGgjlGpbYioUq5uSPiDXBeidFGCS1YJlLBAhJ
l9inCxO/2BwNJhsIZs5JlwPJm/QUfLc/+myOBvmREHveRcnj6R4ny8EYDI3PUStC
Q5/VcQ+OFkXzEzfifmZaVL2uQ6ftC3IXpWF7O9oFL320uxD3McvGNPd1RCnzjgV+
1Lb6Ll0YpkdKorGXrdvujQkPdYYG6p8Vmo2y0uWkQp/cjCUFgauE1LSjGmFhFeOn
WiCNQHV/SUsNbMv6nzaQfyweBX0LKyjjaS227x6nUqhrYFV3kpkajoSqmrVN3Kqk
93pb11mGzQUe4/+YCQtsuWSu/cycnCXHqP2rOGOqSTXXZA2/99PqztmQlmJvknJ2
92exjHiEIbmhCX0sx+NP8WK/kZJ30FWIeiO4+kZ9SGcRi5fdfI3T/KDw7y1eaLh1
UdkPUH62t181eXIWGolcvx9CFwI0gSeKAvviWJYRT7q9AHSjVfK29s0QYUlK/JA7
jgUavnDL6Otina5+ZxPuM60myz0+XJSCeljflO3ZBijiBGwmzVFMUrrMw6vxqZ7V
nAL4UDL7y8lV2Wa9QG9J1GDIFuifIKet2Z51ZR37MLg9sXXGNrDqx1RcdAkZszWZ
TRh4QuPge1eMib4tx5dz6P225SLrd1RCYI8Vu38UrW5whQXemr9qJVckOz4heqGY
DTqJ2XQQGkBhGjlsWyQgYYTzZGGVO4hJgxuuxOJ8k5f/mJ6/BVXJxd5kWCAE+2vs
ngjtCFnPbhfPkpLrBuXZhnD4Lil9yGrvrO75vZuepMj2fNYrLpz6M5ZLzTJn5kPP
IleLpvtXKakRmd51EanIhNaJ5K+ptIEkPDSTalonewOeL+YuAGxAYR6E+Li+HQ3l
JkH0xz8xhaTyIuZqbiegROOlyx25UZJ7pT6tWQ2IRFnx03pFqk2IGzeUqRfN9b/B
QUoDOYTYYqrfQ1QjimbaWBIThDXZIii8GzB6bJ4wNwR2F/opP415YAxQSkm2iUpj
pS2RNUPKP6KY0vxwfNDxucekUGUoNcH8FJvm07JSS8kkENSq8FKcPLyOzyyYXQZn
r7QO1HLH6NZ1RwrBiFZRQtxLjyvpi8Ryj0lU2/hzv6mUtkDNEEL7E9qiM2QBXUKH
xkSxKo5BfSt7hsYk8jsNTOdteTL/X9JA+xNLDdNfzBWTrR4eL44xdAvtRwWXA6QH
C8bnWhOPi3BEexldRrCD9xGo96dLx5falcMOrs7S+2UtHfCRQ+At2vbP1O980snI
bJO3XbHMoJzHyXQQblRnuYLqoK28xusRTzLUCEI14CM5jrmUoSF+vOdhfehZG5T3
tMhG7uXi7d/64PbLzv41YAPr25mFZa9OzWPvKDUkFq8ln74SA+jKs5iyr5feoWq/
a4C8P8fRoSa7xu3t9TqeR3JalPHkgTQnqZ8us9iMSiAxq+AXTV1gXWeZJDv8RO3v
B54C3s4cPGWuV3QqMOHw5/32atE90PIwQSf9kSB2hIrCKY6IiI59owcTrXWuBE+7
JgqFpoAczW8R4mYs+q9JDnHumgKR9vT4vVmiiNp5ez+kFi11lj0vgyqlnsQ//1DC
fS8caheXkp8HCa+S2crr4GUoxZL9GVKP1TEaJqYW7dHM+le8RVdAzHeefOdgblkp
P5SXy43ddxBBIQjiireHFbvtjuVLYVz7Zr7qy+b8nStK247Kjm+PL7GOje0+0+MC
KUr1QY98eX3xXq4Q6RbX2yr0YBja5IjHQlJ37FF7rdHdZYHN55rjB1vmEmQvPFpq
IMAxSXRNx+3kw5l+wb1yINT8tv9Z6IDqaliXlTjBaZgbYSfhsIG8fW5NhHFRFvta
uqGYCC3uuRViklOwg5iZkULZoVZJdBdWmcfjYaMXwnlVOwhBmZs9Try7IBCAlU9C
tO7XbG9RUNpxSnmZ8M573DEx5aspvs7Vpm2icGFnFydeDMwO6fGEAc2oYems5IZn
Mh6/FEWY7WArStk6A+bdlQOpoKa/Yr/2C9GoI4I6AzdK1GJfajHm9qP5Kt6KlndR
WCAHoA7cDtex7vaTxJgPhuKrBnj+YAcw/7zfN6ihcSas18WPWpXr8OgH0DEI9FR7
jyV+XQVQdq7cvebQOBXn+aPFq/o7aTmM4jVdW4A4Oi9V322I4vWdWKvVWqXwxubQ
xmxM0JeiKif8AjcI3Vb+TdkioZGGVMSijfoddsv1zmGuFAYlvNBptabObybFHWav
VHM5Cg4veXty9UXQkg1574YWNBNgjURAHy+s6R8qNaE+bXvO78Ecp0iBablSNMd6
fpDA+5zoEptbazQ71SO+gE7NTCrsS1+LLQQemMoMOGyjBwbIKCHqLVWZD5By6UlJ
bzW8eyYZH6uoZF2u6t3E3P1ckqWSRlbGlhiPaaUPbKk07hyoFDGFZdWcFTLlVrj6
TrTedTGK35rv1kMMo+LZtHCDCWDwRpn7kKFLAYvpJhuYMWI3M5ugpkvIZ2hr0Zyl
bi+J5ahMQprnjE4Lnh0tyFaCgFmrlqwQFOuBfSfr2+AAq48eChY2gxlBK/erXsCg
8ol1DTjoZUEHxZ9PVhaQlldIB2pP5kOEnbYYM7ORLud8h5KEkVoTTwmH9xR5zxCZ
ictrTA3UOi+XdZi3eUDKP5CffWb+kDbpObYlHy9mUTWOT/qSj4NgBwSfPgeLzGyd
qzUMrSq+mVdeCGsp/Pi4oEJ6hQgokygNBRibhqZM9cBoYwfF2E0gJ/o+bXS5EKPN
kfIp7p9ldS7xhv7hjo64uT/3h5jG6dQZSp43asInjYodptDAToEtiJxbQYauuAHi
Lagiq7JIn4VtZ0nPeLflmWl1BpipgrpuYnEFB/mHwUgVa8C5BUUHE/T/dbpzCQfu
BrA9vGgIpKJaUVdJHCh0DWcR4MPBmtLUoImC3VVP97UJ4nOdihmjhsaY6WtH8G5S
JZWqppdpR25phuMCtlCB3y+NTBhe6d8P9BeipaVH1LOT2nBqsPjE2EM70nGV3eWz
mQVjKvS4Nnh3kyyxVweg1xktSFlT/mXOTXQN/40aDfBO/8Flh65sVaQau4lPxTPF
spI19ZoyD/C4MRTZEOLPRxqeTnwHUCKnN+yOI4ELQRaz7uQJCLGo6Y3azxQ3N7jg
MqVZoYALSkP3Hcf2XxECPGIMpsoh37DGBrqeEsTriTmoEo/pdL/fwngPaVqToUJq
X0U0Tto3rBm4+jxUWUxcUTNLfm1P8XiKtMT9yHFZjspxEYNVOQdyFaslsOhgifSc
iTv7WjqzbNtYAeHi5abaQygdtyKAL60YvDA5cPWF0xrJRETJlSybc4ntYWPzju7I
Wx48oDHlgE6WN8yNgf+TnCFD9Gt1lNmKYgEj2N20NA7yzMpe1GcFBX9on8SxVuQU
4uaKh7NO36T9Sm/j0D44em1ZfeXcQ1hmK4PUW6Ki0es/cG1h/EjOU3X4YttE/WRG
7Jt96rRvUY2f6YmJK3urK3+8+C/mFSN29DOFKrKYEHss4PHDe5EVqC05lBuU0N8f
YupZeKdAY+CnTEG7frb4qptw6hkqSj9QQYIZXS8rsCQ8i9hUmN5IgFTWufkNTefs
wRJpvCxxKFU1lDhuW6jCDAKZQ808Zc2+/+ccsY4Z0+gvYpJZ+BQTLASTyjKkQSNo
TGKfvXF56Xz9momX9SsTsA0WIK8U207DC/5qabhlhY12FqqSuJwapHkGAwnrvea4
/zugOKjRuZgzIR6u+YTludQtpOuH0dwfJR9bdsbq9oMR9I8YKggcKVVCePmdCg0S
J2rNwJWm7KnboAlrKlN16aldYUb1x+sjdncDcfsSK3Ftu+xY2NuWJfUL3EvHzMd3
8JP23SzzDppxkybsTnq0lamWF5153eMy+Zwj6Vv0/H/JlDJIxu9Z4zrDdHrsaY8O
zMLl6BcrTkCYJiiMmU8zfwy5cku07WcpB3+6cXO9JGLjfghwgwzecE2H2by8tOyR
RpBp21qPt4Zt0QevurGW2NiDtHfDqsxYs0qDtMy664Sk/tl6qaS53VqAaqRZChyB
ykfM6KWo5ezQ6pUAwFGdbfwmPBBtiVpDeVGrCXpfyXvRH4FHcjaJKDNTv3FCN+h0
BuJ6qHmBgLtmJ/j5X4xmwZWCdRcTmIZeh9WX48UQMsJmhv9E+3lKk8ej91erwrcF
XXuXoTDRqw03PzzpuyvHD5DuR/WYTAsWERpvgnN9REOqaJhui7jR6gS8RFkYY/D3
mIGFdgbVRvsQEAu24CwauwnScrQ0FOwcXMWvD9ImgkMuhNfXVDwPH7WgdFamQVCY
pobQmM2U6YWraMOYsa62W0eNYOBTP1X2+DOfav4kjOa3ZjJhzDRe6HHviprCpYZO
Ou4+ujvoEVjmdAi/k4djRES5vwKMplV98d2XCh1ginibNPLyzu7f+HGPF6E6EGRW
A0Cl2xuzB1v03i5qNR/c3/7PEa1QwSGKQx+lhPDfYHbkJUnEsxGhnbKpWjaG3dl8
WPi9g1CgUlFQ+bajYFUB7tuAzsWOBm8SLR1BfZpmviZLj0/H2fEZE/2Kj1OY67sE
BCi93gQsLerl56vhCCZBNe43DSAylPE/KvgNK8rkTcGw5AXcrXLTMjGdTD1iU8a9
lYy7fmIYkQUU6FkMAyColjxCjmh9J3dxY3uXJIJgq9Ar1EcajIABwlISMeNTwMh6
fbBlAcC78qQ5GycYaPQDiB2sC7TUdZBag7RefYvmYIZzMn+ygzg2g9IBmjRLcwE1
Iq84XTn6vMhk1Cz5yTmDRSmUPdRQO6WYosv+gG5ot5LYeBY9QYBV93uqYxa/onIQ
6i2Ry+ItVwFq/nhstRejIR2aSERL6CkIK7Ys+sskJStjbpBm1/LRTnQGIgwYoSUD
Ln7UupFxjiqJEUyhRPyvRqzN51DxKCc5ry6KEYwGoHd4kLAgYg15YRmhj9vqSC2W
dkGpA1GqsEEWk+zFqEtthEcMI+GGq9Qx0wX7yDX0GVqpVCGybJlrl2SccNRrM2Sq
iNS7MKZf9+95EFq+Kkw645cIh43XY50aDn6YxgBmZASPk7xKnxhvtifXUlLc4zBP
E0PYeDJzMMy+i/nRbv/J8w4COFCJDr00f5vNTCr7Bjbh7/H2Xf1fUyy1zLQhVEhf
LkXn4EOOtBwUq40EZZyTcBMbo90dXpaTtlYTWjqg3GQcxZpdJd4NElZoLtInIDio
sitJ18ZEqcQrHkmqV8I5DtHYnA9FtvAuhpaSmXwBkGjvc0QxzbMCCi0dOGurHOl0
a+F+4I+sdr/7/2VgwWSHEQvnvT/p/fh4y7eHJWXXmY3/k3neDeAVcL9QApwadKXw
DKTzoXbcOg/dej5DlwZwj907CrHCakpsB1C+yudwW/nrahZNx6eWwTRyoM8UQZpQ
vvBnlh9mRasZCh6Z9woC4mIuv0QDtVTy5u3wxOIbDOc0jSuBc/UQdhYvHQsgWGBS
fr+bOmGDVTOPJy7yVp2RJRrDS8zJDRwtLiAFrYYc5lK4kYTK1XKaOu8ELqvhxikq
quujRWE5dSqrUv8F9xn05Rh+XaJyTK0Q5KcCtvY7UNpS8+levK/fbCA0Iy/41dQ6
wL1+6+Z2mnz/KYX92cmJIy5r64HPEoIoxFmqlVlDiYX2kRLnO8Cv44uFMrOiRDhZ
uQO7oK8GVRRjDNXT49y3u8IxTEbBGjHtJDwXR+x8SUrYPmuQS2SONmHwPhckNbUL
vLsU0Bk7cznHiSHzMX2RghVOajkymtZdya0uCOwRU7Fg/1mtjAblKPZWG91EzO3y
3B/JMJrv3CQoOJLg7H40v8lEIUbaFTmwj/JMVaX4eWTXgZsP9gF77QvsFaj0Mhbu
QTksDb68zhJmyvn65HJzbs3B+aHiwM0bHtrsUTqCSxyUFEv1VVk8fJTPvZOlLB/h
qOS33YnyQoPpXBYTUZ34GyEzXbhQyykuXQEku0kDGqEOSh9fvQQ35+c/45fVj03j
xyk2x1wuMPRXKYrNW3gP5YTDoOHgapaOLxY/SzA9gm6q+PW3i6ewKKR9r3xLt2KR
HHjKozZR3gjD+Xxw/5/262IjMa/uVNXyA6xL8AzIpRKrwgvOfsf7ArmBCm/TxEAT
7dH8HkgBiQI98qMivGxWdQjMTnU1YwPBE/oJxmIJJlNdsBdPO5IXvTNbmxGrEOKx
xcBTfd5kEztjT79olr0rMZECrNSgFsi8I36hNOG6eTuYvvWnfVdkAUl1x1T3aSTA
xMHsGCLIHw1kDjfY9GbV3xSUJZUoZv8XXFz1Sy+U97/m4L7lT5bTUcor0U+aQftB
RbHjucQHtd/F/2FQFJTZufkzK/CqrUgL4EiHbj46X3UhBNMgK8wlRn6S0vB1zMRY
CtKPBYJZxxL8dt26RWexOSHBlgCeLsIZISTXpHeFzU044hUvkrF7UGgIrgwBemf1
gS5wo+i0++VyVEGV/RAq7q0YCZNBGsrirmbzjIbnL9YPgOWBwKvj939SdSNxW5Vt
OvM4O1U+vomcneW3qPPNoY/Ld60WfCEm8JWoxSQ2Aw/rf2g3PGdDwa9hQoAKnTjS
pvCQK6mFAvqnOVkMe1RqSMKi+XljrVnyE6oVgjYwPRSYUdy+mqWNag7UkSMtrj9I
8UEs6scohUotCbQ6jf01KKqpLa2btGn/ydrr9TEM28i4UrM3IMNAVSE9oyk527rq
spgaTedBYqPxEF40CJ1eoLmqCKxCiu2DS26Y1S+CWRdRkxOrzANYSdSkuFqf4btX
397pLk5mxvBJPtU2lHx81vRn7ADGQhsV5O59231EAZpTrr+h9klRVIA2d6eVVdpy
LtDIve2a5PrpMTm2vlKpS2ah5JcKXiIvOGzZJOXDdN/p3sVcXboQdK7fF7TGLI+2
VWhNLbTYXSnK/HSm//4HS/5Go8NcDZziy5yfroQA0R+SCCb8rYZTQWipKWQFSaE4
twMqseDvCr/Gj6/BiXhNhSMolKHsG/fWbuVeBzg72YWI6xWMmKLZlGIFZua/oSZp
83hkDldHiUExXgVFtUhH/YgO3xZ2m+2DKP0LjlZefGmDklIWcgdgVCIUfUAFP5os
PNP8nwegy9XrBkXRVfeKc8lbsja9Bdp8xi3AV2FN24qOEkMqkiAnLSVSc7f0NhSS
s5+VyY/lIaCC7fjBM5QQJpMTH9Vq2V4CpZX4tWwcq/I6vv65SLwzaVXSQK6ExsRY
6UAZc/6pA1r3+bfVhAnozVLEDHaqd3sXslCtH5c142ZwDrC/MPpNk0bccKpEPrky
8zKGySvcBmm3pHtnA96jmPF1grOp4fEB/pwnyEGGYUdbm2e/X1M/CedRwGDpHj1+
qPsQtaJ4ifv4MsYLpFDuXCq0Jtob/FP67OLvbvwwdq8SywSQCO6axFsC1eleJT4N
pPG9Rt1O1uAdB7xkKNJA9XkOi97inrH537qeamdYD+dM5W/40G8QNEPqTD/VEvOK
W8YlV4j6QlZysiH7LWQQhSHMjvYrWULIJRZsThWTrUnoU03er0piWM/L6zdHdvgc
FI/IqPo8BD83POHlilsOkCnYo615hRmTxrv7mGW/50GqDaCVsLNO381uNB4x6Jnq
C9G4a54W/b3QjR18hm24H5Gn2aIpNJ0rBAtHnaB1fmGc6kmTEgSsEWyM6zq7yn/E
2/0MUqdZSIajmt4TAh4GKmPfHsbtuA+yT9+2q82CYAuxd61jW/PJmgLyJI0RVJ/r
ZX4Q3yvbZu9Yu+ZEzNg5T2ZqLfEU7F5vOwB+fy3HrLAOeNjZz3ZWWqwtWwRbqKVr
JkX7tzxliDfJXc3Ov5K8Emkhf0aR1xDySuscS/Wv74wmTrQLCKDd/9TaHIe1tfYo
zBDhFjETav4NOSMphrVw71lxcijXKBMLdewLeoZr/m60ea5b8XfarVeeWi00Dllm
fRacn53961SqcHgMuphKrMwxkVQ/K+ZZS9pqknt6VNQ2zvcUjfBaEdB3ihFNvcom
M+w3U1UbrpA8Vd5YCJOvbyjEYsmrhNAUCPZ5g7pk+ZoD3e8jmip+TMd+CZeyGdJh
0fFrHKbdeiKui2VXPaD8jwXzzoxQogiox1q8AW59cuF22+um4K1bfHNWEBmSbTBV
uBFXDdz6M/0WZkJAGKD5q+esrpvRbSGXz9IReRDqZ2aNSolV3hbUyaSpsuVkc8Cy
Z8lNJ2DyFTe50FWcGfZ/uG+mHsLfwuSeFn1zXoYWNmU4q9NnQ2ms594jiKiIH7qg
10RRpEGYP7K9Yqj020XLfs5rNocfPB0WWlvm9Mz/4NX3VrLn7urGmQUb2GRh8AYj
4u8tffzL5F49yXuUGQG+qfqyLdmlcsVuG6lARtdWUMCYBpu5+aeVAK5hvt/qrd6z
teG6aJ2ym9NF8W+zyQHlwRtLs2RUdQSNEcmSPq454nJpjKw10dYopSxOy786M2De
IRGVthSE2TrgKOZtvOXFBtRt8DA8SwCCKuDPOcN83sd+df7NfmPk3+oM+UnDNONC
OviXTvY4gYhXqCxZ3Wz+uGWi32JOt7q+wLu0f7kT51mmzKcG+4e2gx8T9KqwkrNw
n/RUakQcnyiC2WsV9//mGMrpOLuPj7h9hCrA3dtJqwRkXX3+qBQ3uvsYS1wVvVDw
axtmjVGxxxx9j0HOBQVqaCwIbQHbW7SZc7Y1xcei536RVOPZ9rkJzGzmlFMoBKHA
k5Ei4YaSstp6om1Ni6welw==
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgDmaPortRecordFlattening.vhd
`protect end_protected