`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwrYbPr1+J3Tl50R2qpolXhBnNh1AUhLYXwyc5pdCrzES
ilWgnx0q+L6/4mHHxwJBeKC7bHipIgwvRM8uyhP6akLZCRh13w1NzdEA6y35JsuS
5s+dn+Exm3ORceuqwM1kSjrqBDCIKxGoe7tQ5+nd4swcK3jpaJBeVRtBK7wgRFUM
iC3VChf4sHfl+I29AM2lF60NFW0UTWSEYazTm7uhxIn99t3CpkmhvrcIphnmn011
uMEi/HELJoRM895e8kKUzCSUVmXwYGzYP46yjqgJzU816D0XZHtqk9sfxq5QVJyt
KocXZwq3qH2gAbGIpMFNGAe7mvVnN4o82ceYC+gi7bQUQIzhFQIMYpYuTmmDY2vn
Ya9/omFVy9n+bT8vwG2PPsAo5f/0qPpI5NEON2waP+fkzPI3oKjSJMWco9Af6D/B
UTE/zQ3mTkZxJwNzuxH7hUvPDh//LmKaQ4LKzuIkdOyj3ggqueX5opKk4Fn5tFB/
TN+IbhF8RLro5vcloOtq0wLIyE8Boz+NBhNAe5XlB95SL4OMdQ5FzuQI3upiYJBS
iR1jcAbxXIpc2YdawnSLxPuaXJGzxEWv0q6OH1aDqTyD3+a3Ru27k/PHEJP2v7zO
MGhzLYA2QOpzTK0V1bHI7jiJoVq+4EdPCcxp/M7kFkEEQKUo5uTB76vkbHJE0Uwx
BfkxbRPUCGsdjCgdZg6EJporgo3VG42bVsEAVBDiITELcMjyrO7Sl983oL8ZciQf
OB+ACDM5MktrYv3G7h6V4Ed5jtDvXyi1vWOtRz2mZ0CP5DmhUW0XaxNjh5szSspI
6etXgv8lkztOwddc4RUzt9IpjRw/WCmGQb5ybN76zRnmAuzcwEenWky9M0IK3XMu
yhTwB71t4HkSJUZwcx9fdwOF+HnYQU9ITjLX56XyvTVwS+ihQElAkbjuAYN5i3qr
WipCDFCOD+KDiUUpGNyx23fpgKR5Dg1YYGbvJhUvOnVUFL+MKrVd4jieBQBbrswE
lHYpc6eeOHr7WnpUKtToEA9SXaQG2xnuup3WzuP6ZOULg3NOdzRIMkHomzDxZAve
kylmNklV0ZjdQfwYt06bKxISZ72BLT5s5NlomqK1sJsDgpO+yZYPa8zYtWL0oOff
BQZw+/VuA5BjwAm4qua1vW3YyoTPQ6fRhuyDIHPnZS+18ffc4hyXUU4SHPVNI/6/
ZY5CMu7EuK57cTcNfXsKwIyR3LeuyY535jW4KhmuJ1XRTp9F+tAScLtmUa0tEyP9
4RRa5Y5RVX7wagl5l2G8RVvgmlHGtIlMZufuJowyjrS806/7ao5+GkT+5Hg1zmtH
dED4wMOa7BXOZqdy4Wu7lr58HZyahhxMR/82uUbVlG32ZFpry7pPuGPyvwKB3QDr
4qhxGMrkT1IFM3+3ZAyqBUm2I/YK5eX1Ff4uaOhjDPjlfyKckjkvxSClKfMZoFG1
/4QNiBfnqSp/kKYWvLNdX4E0QOlwgiHOJT81X9RYFfNCb/b/cKhm/Qae0h/Tb4Hg
ZhWVMovCbkM6zoC8J7su7GD7B5G/jTwQbSWRKq+cuLEdkrFBHKeUvDyEMQ+gEnyH
KTZvnfpyYGwqyThpD+Z+5PZR4CFmDObw2AfJWwIiEMYEjKKU+a9nXC/r8wv3RyoC
yBj5yVmN496d4s5NIdovdSkNJKx31spBB+NEPQ86Kg+/pOgdkwBMQg0vPrgzX0Cm
IrPsJi5gLyI+6sh2eX1G3TqaL5po9/vYk1VifP//x7uPFA0xGh/0QR9SqcHfYPwj
YOk0D0D1h3lLaZ038JeXA/27ETYsfpgoxx8IlRlUz2PjKcESHQChBqJ4ilJ4Lrk8
n10CBlwcgQI+fSZkW1+zTq04wziDqesGDjMu7YmRLaBKfuLjg+wyYy/bk72kiD/5
QNxf9vi7edpflPhWRZ57YDUHlzM2qPO9ZVLQDrsYu8jzP7HyiM+J7c3fUoijTfrt
ASgYZ+75TknQksSc4oCNKYmpwIfDNMjj/ZuSjDfAy1zqgFeWUxkrVFPQKkjQXdBs
gsSqT1Nb6Z2/Ys10E05iy/TJ3D4lD2qSKMl54Rlo6mXQbXQq6Ndl9XSaIMq2gKTy
yq6weCBKdLNFKYyQm+ZXW1/zK2wfKJ73ffvnmpkhD40E4Q/8IMUt7VXs0Le3NN9+
T5dRqK6Fv6IrSBsEPvNbxf89RFdxmWQO3Tsnn4jNVMkIy23cEdinkRjz/BGSnVQd
P5UK6r7F5YqB1RBsIMDgrdHD1swQYzeamXwPHV/CoL0DW5pJzUbc6+YiWmm6wpCe
jGT2SwIY+ooueWZQs6aC66LL7Dafr97F/RHd+rsPzWaRHTCojJo6LArvkyQqSu8t
qNDU+8XzbLo2BzYPDdX1VK3jh7ZiUnQdxw3bm1hNI4gOy9CWJmOyQDRw8o767ls2
X/Jezlo36mc9+zvpMtJYBmB6qJ2gCdYM+jPWdVVrBR56HUFxFBM1Uk+XoIqlJZGh
dW2t87zH+Umh4nwKUQTU5FFKPjNNOs/msoFd5g5QRIBBvFEAoJGuH3NU4hi8FoSo
akKXonUvtoNga0qQaWPOncnCBjzai/fvjnzZBWxkRTQsAtuhr3sdV5rLrR2iggPk
kfQz5CttXDm3RxrUX90UzYhUn0ksCOf9U1L0+RB40UcoYFSxCmeQey/ywQ0KZX6Z
o8SWCVqPgRsJfuTuxWYzSFM1KHzk06o4RTw4DyWS+5L4x9a4F2knx07F2UK5dR5Z
wWMqo8J20lL7aZGO27xYbIv70kwHJmOHWwINogk6WRTEipfVclMJ7lKUhUVqdheT
ROspnzjh7zRW6kZaKaTdeod+p+QQslp+WxD2nTNH8AAPo19SwgOLAq1RSkqwqU7a
qaMUT1DfPdQViayM7ieBPOapbMjWwTxke7lBEpI1ro9+Szu+Vqcefu7K19Rd0ak5
imAny457wBKpKBOebvq6Et3VzhKYppOmkhTSO5hJrp+d/XvtsX6mB5WWgpBJ+3Hz
hCRuIKzAPzvyXvdkLpH0j9sI7bNR3KgM9pj5WOewTdgtux9gmDoNyeFAOTpt0XtU
iz4qSdP3QQn1Z7Knz3lxdhYFmaxfjrMKGHEc0T+Hy0Y1uYc2is0d305UCm5Ue1q6
jJA6eOp1arfdp6ZeJFGZlVGqRwGL2f1NsJ1hRE2sNdrz/lLLE1+qdcNN/a4XD/MV
leYi0aPqXVggtTpOIAzWcvTsDjDbsLxe5dmT4d2+GzyAM1iZGJBFFFRx9YtQGIm7
kNR3JytdZMaKt2J3zCdLCty/u4aQaiuyRQvHV3U2YpWn0B1nfakdb2omUJ62QwH0
ER1v9LEsSlxml2WSSjiOF7Gjyhw84a7XWIvagiFWL2Rvc1KuGGsXgyldkzW2R6dm
0sUWsz9DZowIUqjiePUtUUfSSgCA9WbJMNYbymBeIZFWUockWNZ/1vxrVzcn459x
s9ZCKmdX4SF2kMEXi5d1h5Q/ghreUdM9j12uq359EZJyiJXJdG2H3idAENH9gWjX
UqBwhqsQfQW82sUS5II/6lGXoOp3xsMGT4SsYqK9hpyiYwmtaLquSiKMbSiOF5NJ
csGUjHToJaWESODpe0kbw+v22D4RJx9C+iF3rkZLHuvwS9n4JeJeg+77BSFMujB4
7hsFPoE/uf+PI01V6uaRg5VKy+1XobcmVuoemikAcyXS3+yn0tevEzeUhRhtfruB
Yk4GmAVNLx0yx+J/GPsjnvzGP5b7gXd9g8YeJfpp/rd9fsak6pHjmkvSmqenEtx5
ofGpUy9dH25OCQCajLT0fESlH1c+RlnoyYUfKroRdnc/P6XMSq/ZSGgR91GSGaQd
G66Kzl8IzCYxb8FtLJqJ7Px5McNjMFC1XWPoJP3d+mBO7n9tYdcPKBA0pq3rTJWq
hr1DaJqsRs/aHAudj5SmeVpiJaxx98MhpbAQz7f+9Q5pVJb7JKh/5Hfl1xI3C4dT
j5X6Rlp112aVITrGtoZ0wobu0AcrQKZer4Ojytqk08ZEZiNMiYfVnjzRDQLqu8lt
pvS43ZoTytKRNBvLtpLuV+qigtRFM3aRumI7WgZRmjC6Y6f1y8dSbn6ub+Q0UPae
+2x1ZwRi6LwzdPwvHXDGJP81GmKRE9Skq1obRuFSx7iC41XR4iFNfkU/LCDEB7+F
vDhUlNWcpipt7Fxytmf8JhppD6kFswmoIYQWuCKyY5WaX5yr8Q02npKFkNkOQs0j
mye51uQkIYFiVLMYEFtgasGu51w+x4qcdpYHIWZ+Y/afQIs8vaoT47jWrY3+JH+b
2mEUGbwWIeIEzUnQhTNwCmKg+UDkRdm8xGwK6WTeUkXTEXkqNvYchiOfKOrZlCj4
F97HwPA9m+81FsKSWam/mkh59V5vtZBL1axddQ1aZiCAmK9H3wRAd/IhKYlxObHB
Nd70ZXp8i3e51NSRd6REZm3PooPZQR6O9+eXrRsqp0xFpvf4OUXgHmT+cM3Xz0pL
ue5LUtlVc/Mu0HXLh0CvpS4M3TT5I0Qnca2ApfS4DjkGUayRCpP+gVmOZfwkeSpj
NChd3cpAnML7ph5++P4evurMeSZIXMH61xoVDj5/q8Rxda/phgvB/OMF5m/WGz6F
fQjuAAogWhiu+HB/ItBh7/gzXEnh0qDRT/s1vsomRNRVeunbC7bAB1TKALSCx358
21TcqeTjbYaGXvpH03zRtrpWJljzS/0kuBguYu6Aic0Yk4q8nKQRvSy3p5v8Oj+b
sWCOC3POwXf2Hfx4zvoQOLjxdVz2etGA5IRCl44E2NWsgSavGuFPTTgnLqY81PTi
Mybxc8EOSIYugmuuuru7PmOFzHrEd0qlht6mYclO5u7UzBybjdhz3TJnUKAiTRrT
xzzWS/8TnL1/yECkQdoXobj7AvFltY8j9wTd1fTK8JZdTj93YhTW5JqruLQqVk6t
sFD3SXZq8EFVVenrft7rW+6D1yK2HfT1ChvE0nnaCucfc0R6RuLQ/r8+9KgHArB0
UjkxEeOHnxvZtJTuLuNX9sdkssw9OZEWWe875cyUxYoglGRg7Mv5GG+ON0oNtt7i
q9cmX2mb+1TJU/QtUElBmORdvqaxxnuWkO1EimNaBam2d8j/IhCrKfASS4fkt0ku
gF74cO7MOEBb1LDnmnbYMTpwB7W/mLZqRI61856CeEgYiBqxa9a6gaT9Sx/tZ1ng
HUcUb9XKoeHXbehfcGPYg8BfQvbCvg/8KqKxHDrhlVgFEbc7wl85B51MTfahOKIt
dqJo8jpVL3NdBnUp+3W5/JKc+ywd9WIztf/Hs9wX8U+PBsaExSgwTEecJcQGWW18
ULu/ga1WLMuZ2d1DSH/NsZzVKJr+OaWCeG4F6+mK/UqQjBjMjdPo/b95nxUAnsyc
c5H97wHFnnElcTWTGklqQLlbWM9zSZr538dmO7o81DQjIi6paZtssP8BCEhxXUvr
l9KOjq81/Hc4k5mYxP1STVoG3ZVc8s8U7v7NQzfALU5so6BGcQrBzuHLC0s6aZao
KLYFijKYsix9nsKqyldVlqrQkN3w0hz1XZHFShtLHKrM5ukbPIrsluGoqapaDs2j
EFh169LZKepMRWgHhETo870F1bKA/90du9UKPN1Mel2aRMDRTSHk+ntxajwN8r24
auyUK7JinKgl53EDffEm7lT61eITmnlcBSOV8Vn3BY29FqLHG6M/Yislr+Ho/cMh
PCu00xqPW4KDS7eMJyNcx1l5LC1/oymy0Z9wn3ApaCxNe/Qsf78yV/gF2R8T6Bnd
dY3XJ/6+EjFz6POoh4Dk4/QxPYXb7Sss9wTNPBIOkpxPfzx4w1CHLmMcRAqlyXVB
2+yzeCgz/THkgoKS2DmtbKnCAs5SFjncZVXPFUbvFsn0I71AvQRhmIjHyh/ina70
uwyu57bN/uWniEr/6+EyNQAHr0xGT5Ypv+4jD1o5Uhb6jAMC4Z2Yw3Dqw7KLwXJ1
YWmPAE2mDvIaA2t0lp6+cjykKGvTCtPhFvYYdMdBSaEiM57wCRyCo6sYxQeITLuP
2UM7ZcJfIGoJ67sYgB+kLIyZHUpSaCX0JQk8q05JF2rNFsDbgYnXOZR/QAOfsd8Y
qYIuQQ09u1nfQIXq4kOwJUDROTDWMWVHSQGAnjpER+eTQwSxOPoIhkES3AHOA4Lx
KmruMJH0c74XIu3fNZSz0PNRVqaLHGPs1nAcAfbAEdf+77CAOjAygrYDGm3dChC7
sXU294ywNhtAztglMOL2ltgTiFGcOHl3RkP/QFglR7cchj03IWI7PT+fD/GTvsQI
TekyDv7qSsHjTQTFITMzqgmSFBsS1iVmEBeQ/sUCSlp61MM+NWD1j3wxL0/dZXro
Zv+UjDnGh1Lawg/CgFD6DSg4KWT4zDEFJHDw6Wc8rwyas1qa39nlzIuY3SQQVIpJ
kgQpIwnGOizB2HkTKxikDYNJUk11Y+g8dgGrT+jSxTO7SGgbWl8yj1mhts9r2Ypa
5sJ9TUZgA4JmMQcpfjVTi/EGiyG0cyDU1IRih6yT0SpY8zMOKbiBnGUz8ExQvw+M
0PwAm1hHRPOPh5Ho0OP0n/RXFcGNkEvCpwrb+YDFqKgKUuaQ9Dork0scDbZG66fm
avgH+ZnuvwWruoS4y0WDZXF6cVA+iNrhPNcTrxkGr9TSaLLxnJv/PCeDf9sMjk6P
nMoYVgb6LGAk/aznpDmZBh7b6Eq4H7Y8aVg5fI2Ed2xYeyCT/m8XWvH1PwKJoPV7
LrJ8J3Tnjco/w1eSXc3X3sLd8/mYnNAr/dPZdrJujtVJ5bvAv5twX6Z8QjziPdb7
qbBnb0uiC8EBqOa4ZXkGA4N3CrIdubdJOSBQJnBCzE3gw7pyYnh5wADGLa8PRIaY
wXxWckRXeb0eJeUT0XDtEvvNR1oL4dHnD1oRzsvtyweokqlOngdVWK2i5+4gAldI
htpSywbGGNiDA9FPihjC6rUIWW4iCqqsOUzWXqEYwdeNwMcQaNnMQAq2L+wi5Qyq
EU10KFLR9LMZo14LYq6lXEf0/qW0yjMg1m8RSqdPSiyHch+BY35E88TFBAXN+1aC
L6ZBYj71l+YgKbQB3wGID8O76m5LC57yBniW2NMvqy6pTOLW9rCpxcMatbclsjl8
md224elCrKldbFEfKtGpuZ2g2ZhbOp2h9qsRV9lA92483I1XvhZ3hs10D/LxVIMA
ABKtvmKYp9RrKdZQgFtd+2NWsZSd4rZN43lqRhRAXPJ7FLQglypHS+cQ5BuQXp2+
rpY8lfrxWDYPe2/IojbzJBLwdAgc3aUlzFvU61WND4KPuwkab6gSczcsvOtmNi2H
pkCSH0KuuvW4PhgrWvE7GUHHm3FjjFUpDbEefi53MqWVkuJed+UxoyPxUEpxDhus
QC6u+hrz/+ZOXe3nT1YtTcJzQ02fxDs9TCMTQZDlnguTV+azMvTQdMfKfQYSu7SE
l34ohrAfSJWmHFYCWpI0MLE6TwXSAAmp3MF6DEEEhKsLQFu/1hLG/BGQXangNr/V
CJTW5txJJHmf0HDZTkXFkf1bWu6Zvr+0lfV/HzxT6wCB+00Lpv83rhLAu5BVAE1j
sVJWlA8NWUI9dXz6DPZIA62EKYh1CgD0rOvayPz15mQK294Yhb4nVL82SkrzF3zg
X99vgclRHchIgxtWm6QRc0rRre4MD1Hlip3GxxLmCFyg6HXWIPXrcbwXJDqKVTsZ
mqv9yZsl98wF/Ris8GCcwgcqpZUszVuTc0WmxyBkwNEaxmfpq7Gn293iqVzmWJTl
1Hh5U4byMRc3/YrmIDLM995RRJx0RJShxs25oTvEgYE3PNXM2ra9P9tHWu8c0VFq
QUvLzmUIHrMpAJGzPMiJaL429EfMiRakGFnSXFFOgZvPPrWUWAc/8W4avdiAmpE4
sLpT/0Cjmx8irjXQrbystqPs1WTtToohJUNhW0CtLWoYfpHS5tQIJM2d74/VU67D
HKtrR0Ztr+uokhSvcR4li0MNcvhyglcu1Tv8MY7FyNK7nbAZZZJ+/puBb7h7evzd
OToXdDVuoVgY8ZogCRg9z6GeNbhiy0CpD78l5tpbffFmJYVjxFp+d3blyOfxwnBn
DSSx326KoUwg4FOUYtaePnTQKJjo50XN51qZNvSskVRxO6gAx/MlVvrSwdAjAiiZ
GHLujqus4mXfoqPlxvMIOWJUCZY/dRrwt1/0C9b4imKSYZbQJSFXmM/T2p1tmAnO
7USN9bM/Nb7mYlqpG6wH/OmBlqclu7/ETQkrNYsw9XNaYWzVv6mH/LlB8Ve9TKIl
IhzQ/NuC4gKIAzsi+E/CfK5lqZn3o5uHuZOGr2ch1j2h91WKoZ8oht0ukanwmqyu
/XhQqxV7pOHWcypqScVPuA90V+EqKwQctqCs/qXKvaT9YWhcgw11H7dHVeVn4W8T
SR5OgBlwbyEAjxYcrHX8be7VunkeqRu6zmthm/xEa1KPvCsKMdHFirSoLM/xAG5M
EJ7RaKdqfG2lggv0Uo4QA511ek+Qxvxn6Zof5I/UniHlTanGmUuPgYNZyN9kwKZs
5Feflh7Z6v2QUAZ15Q8YNocyGYeGv9itVnJ2mqzOaGSXhInSHtBLFZ4GisEwNoYH
hCD6r0oL2y7dN7fKl8t8Hx9uSCGrxN0HMtbDT2qnBjBVTvAcXBgATLxE0QTN5rPJ
AKXE6/22K74boWOyRGFpCfqo45pF+ViM3Rjda84zVUqCtf0x5J5c/dohEA8pkQhU
0CWrWooUyW+nxpPhvuGGGcAk7CkNgUIMeqUGiEOiPQ8KM05vFvZv2EXDQi09MJDG
+5h0CS/+nl2WJJ5X2r6qYUBgMDUNDnht+Y1lTObWw5uTt61+j1ykY77Fx0vtmOe4
dNVTnEOa8gUsJ32JpuK9HOsSQcX5+x4ZS/sVZiiDeoElkr8LkkE0x1xI28mbWWwU
3HoSxP+48HE1P3ebkNYli4bqBCi7WZ6rTLniEYq/4KYutrQNAyzQMpjuckCqNfbC
jBEavegpqumZECJv9MRhX/MfG1HgUC/jcjUmDe+dyltMGFNygoUe6M48wAUy7m6g
l0wx5Y6jHPmZ5v+CB0fPJvP1/jK9Uw25rSAJnzvpaoZhnk11nLjnwC/gdK50T02A
M5inlAcwYdRZrgPvY2vacp7jfqyUZgJKTXzWXWYXdFBVFf7bcR20FBj9p0cRhFTK
C5JFXvFG03AA1rC12rpaeW8ZyI762dX5K1Uz+cA7YEdvJ/erbJ5EPvY/Nsv+P+RT
9oGwqd/oh18fH9YCjDioICLElG1xZxwP21/vl58ItAqSCJG+0vWxy7x1RHrjcp5j
EHgV8be3L1txyyPkg8RmGBMdFXOFWqhf/IPshkDq5EZtynkzKowV75yhYVRV5jmr
UrI2uEMxCI4+IX3EtSAgx3WB7sfp4+VUgIJxB08a668nIHi8VA4iAb5sHsUgL9Iu
xMcxx/zN548oYRGm9kCfP7Y9Zi+8RuQhqScHOun+OVKgnr0LUGDXVNYLY0TOXPU6
N35EmSST1qFW2hS9txkIKtpon3qsdnNdfSwFj9HZLrwQm7erVaGBGGUHToUvJPDj
NQ2EblB4SKzXo9X7lwzHGwTMt/CGDJypf3Rq8p3PEVIVVB9rW+Q8c42XQfWapmSg
XxkWjRkeGdizYNsePzbNHCeNdwwck6TvbjHZ2JQ6PkrrVQxVlYR/yprUhyGff2aL
66jJ21aDeWlWKVIWe+T9lChPFzYis1Y7CjOBkY9y25wHXKpYf4VkGBQ4iQp05aVg
hca5kmbNGcF4oX/rIkn7c5EVDKgf9O2HRR4km5TzaTCmbnHzzBC5drBVm6t8bmgO
yLKvfPEW+YS5KSutd2ydSPdZ71OzLfeZQvXdzstlDzJczdVDVqJx1dZyPpFFvxEd
8bE7Bk0U25xmDfzhsEyi4D6FWHTiiK4zcrebXfMTlVwcRD1J451MAwpNqTXSsjmk
F/6fIoNi9cBgYLvhjpUJHKSUp9HlJrYUQiyNthBGnh8gUTZyCGr6ljzMNhwfFWxa
Jj1VhBG4VUxw/0ECaiEbRUgzWWrMLTlJawfp0zeKv+xrahW7e8EmoF3QStbLBgWJ
d+P6+gcwxwl4fpSVIzb2M8lnUnMCv9T9lNZjj9EhOckBYGiS3L8hhWzFxse6Whkq
92lu3bKMQcG6X4YksSUCfAWlQRs+n22PUxezUXQXH/pUEF16QMZcXfWTIuRIzwW8
8RspzE59x6o7wg7mAw5RUj2eA3bgyG6QCKMn1MAv0uegM4vWO1ZjsZMFE5ZB5yb/
AqRp0kQYcVVww+q+FzTwMMspnhAon01Wb13wayTNBeTNArA/jQERcEtCCp1UXPvx
X9p52SVDRRSMz6Or7oLEQvCnmVc2xXXxd5KyjRebmPvVPG0icU0Av+LX4yD/6l6z
tWUBa10v0dqOicbMJU/oXaWN4QvWZQJSKnFX0e7RzBHLK1tZWEEZ4VdUZoXAizmn
H4lkPOfy1ExOSzLM4i6qkf52/IX924KvzeCw0BQr0qQcRV/BFoXPGS7zC57ATns6
/uZA6AZX0gzp230q2r85x+BvOpQjnqpesIiUTUfAlXvd4TjqRgQEGx+MBKgH8ITK
75B0hxzfvtYbGvCrzKWktrOnNbMkHjoGouaMSe/1yXNcntsI2Mkr5PLTNTLMiBIy
AwosKhMLAM3B7xgPxuPGKqoFDcZfeF5drnfk2BJueaqiCAb2/rSr598+0CQyQGJx
OugewD5d0eQ1r39nTVoGyDZtLYKQ4kVBCPyP3T7Ic7IOStERCEmXcqpBvQ46N2Lo
mIMSemmKBMpjBb2zVCeUNFCiyuoSSDT37bkPNhdrkdNkuVmRIhwAS99yUIv9bfVU
enKXmHt806jw1mfpLBlODrZZixcrWHfaap70zXepcA+15G51T0aaJzdmUJ3bcnfX
ApSl4w+lOeAz9Iy9iw4zeOJ+8OrvLRSLM2hvwYknPhCgKD3UQyTEAWCSBlK+uXdD
zv7k8WbuapL3ScAfoxCYcwaYqG3Y0jvhqXEhIQ7Xz/ipV5zJUHJaI3h+oZ24SDzY
9pUjCeTwds7J/BXoEfYCDZam3fGUI/6k+yIAZxLp20JoQW2lpb6wTSLGMf1w3+FH
6zJ6MePcab/nS6UL/C4f2khEVOBQosL32OSrGYjcSLGyuPjQO2SeSDpUluzQCI2+
LjVUWw6ZgCDBeMhzzk76UCVXk6gNT7Zj2C0TbHrH77FXYZUHwInaKE66Lcft/MgI
OiPq9fzORGfz39Zi2zecmV7/cPj48EnkIwlZg4d13p6JjhsdbgbBSa69drtKjYA+
4eONAYN07hopItb9hFlGh5fuHon60GQme39CV1yWnegR+yxn+KJJkTwysiG2aMgP
Mqg89tuPBIhbaEKrFy1B0JUPmf2Kl3Z4Lfu/bJ9qcqwSSSRTW88gTG00Yt7sFeO3
iQ6tvyuGWF7Ps2tdEn8Bhp4UiXJClW1bb39oZljiGJf2FbseIkxghkr/m0v0kkXt
kkt5WRpS3UeEPoV+R105PhBccL2OMU6Lyv4gA3S5bRJN65DEIV/OKERLGVW12nAI
vSTjhXiv+dcIZSimEOmPdazyO/p65ocoj14hg/XnIe9Zair0E3Rp6pQbDMx8WryM
LPh//yWRBJ4efthW0ItYegQTg7AEq9hYL+JgIF+jUJEAG2/VSeqbT0XaX7bUZTd5
tl7gDDggbwFhTuzAtImXeAJ+a+ENP1+6QtRapkHujLY++nItE8286Kppc7tfrhuP
fmNmcqviPFTRqFfainA+Rv9GV4vYU89nzB4XnlZvDlFXiFxY0LC4Tw+HJzS2aJud
j2BF7Yc7Uwlj4YkPDjeVahCW3EVp1Zyv94xx5El9CDFhGXMiYjaO7iyLvDEwXbl3
FyEfi1+lZ8nxD/6y1UnhHyNxYV4xPjpMljAMEN+vZYEuLq5j+s8eYOy92IvjQ7Jg
9oUDidJJ5hLJCYFp1rmsuJiI98ppqMZsgdFlsYAaU4scsfrLowB5r2t0a0ZfYYUL
G79ziCSHta+LrL95NLyoWKv87PtqJN6rL+U1p34cDcyI0gM8JtM6btQjPECgaqmV
idlyHV9OsuUO1bmxh1MkZ18jRjFiTY/AMhXerRawdBQyS/+oM7CxMB1oID8dv0gY
VALXcmoYp01tkSbVi4V8ZepG/Svq6ud0xfF1HDNXRKFhOydJKHjgoSkj3jMMfCyv
g2ZOkB8lO5W3pFJwz5gkn6AgFalipCaCuW1sSIhioaiTfhjIfo/WV55/xsmtNVT9
FqZmx9HAqbAqO1WeebgN/6C4WS0b9O2SWkXVjZO9vJD8qhfnD6CxyjuztSWP5bt4
vpxj3OwgqcHmudiZLOhme5RvAh9nIftWKd0zoiqZhtQA4bQUa6Q6Js1LoTYUtZQP
SBTu7uWGUhjzeBTNpUT/CBA2cD0nd+KSMqtd7H81J5JQp3a85B5jn69IkKvB0f9B
rf9q+tceU+EVvvChQhYtKrfZge61nQ5nLcva2pUONgpvbTAR1gXw0Qhf/Eda9yjL
TS7ClSLmvOStwfGUz4vhIi7MYJmtUc8zaubRmOb2+6x53d/oMJo1YYLVvZ66sFDM
87rgQB44Hpl/lmU3baYSid0L6xkMbraiTGbsGzZdlE8H1hpHQuDLvJ4fQV0OiZn/
06LYJ1O9g/ue2LXDNMN4F54NAiMryB8TvSxR5vfyy7n/9UMrBSnYARwwTV1FJtFs
JgYMGOKb5wWEyz/tTJGll3PnhjfkKPeeZwIaeug3dVGiefRD+xs9CZcdKcYeMeY3
ok0N1jvgfdFLVLBtl6itEGMT+t6AdfCfUG8swXsuhJCjMGALjyna+BaN4VnPNjOX
/qF6TFhc+uXYI0CX2mmrsBXjYvuWD7uqaPzHdO3SUo23npJMRMgULsV+fuYbsMzs
I2O47w20lYsx82xsW5UzcEUcLqKuC1hYbP4UeNQ87K7Rb2lrIofYj2SXMyLDYc2u
REZ+URu6PRkc35Zxfmup554At7Wt3dmA3FeP/cq4T/7HOO4iW1FA/KwNgO7gYlc0
TVFOQDH6Yz4brDq7bW3E3KV5JTvcdxNPJYxcKbsj/KFNRBN3GAvgj22IbFBvZOkv
STeFrgMEr/IdOnK9GR2Zj/Dwxx56+1jpZg6QXDbQd8bKHuioDPW9nQLaxhP5szu+
sTI5oNakt6ogyP9w7IPTLN1b+IuhyF5w3Rg/6ggatAloU1qId+wUIZlrd/9BJlhg
paYogFGYAZbdlAIzF26g1zDpVF4vsjBvHt/tFe355Bf7Gudz2P+z9bzTiWu3bdVA
1AGHX8coTfQkQ9auUW9g8F7RSf2Qt+0Lyf+D8VhqtSCQneRNlLemEyH3jUPslz+A
CDVUUVBi+D2cMBHyrQu9EShaY1sjPBffN5gdgG+QulGSMujJImZYhGvEDwMTgDiM
SEayFqeGiq1QyLkyAD6oOOMQi7uw5Y2eHcX1OS2imGc2r1ItFXkStmWEzZn8NEeZ
CdxLWCpgxzCpCfJclUW+6rGMWL24zBsv4/dPWCA9ynP9dlRflrZ+IktaBh93+N/V
nRyG2ylKK9UXkg1W/norQTeXVxKFmzkvEGzlpYprAcjmGtJKplXw7QSuaXHPWBz8
q9z+eisTfz4T1DglKdt0YSyT0o3Lrw+ZkRSSeiEehoHk6SqG7dTTxXrBt0StcuLz
s2Gq96IQIDfEJNE4vqowtEZ2Y2icP0xpKTbahQkoyYVtOWSgEd8M19EMYn1oVwHp
q/ywsDmqug/hfYulHl5iiKsyyomAMYqLGLKJRjcZwqEbmOIpcizN6r6fm00UwzAQ
G7gJs8GCgeG7L4fiwMUe3txLHShEXaH15sKnDkQDtAXgmZ6zEvP6bUK6AsyyD+Y6
y3+YLdyfE2rP32zrAO1PuwLfZfR4rRGrFzsxwXjIAemlpkmoSKsl2+Xi1+raENd1
JsRErKGuqL8qaWB59liPGO7HNOrvgN1LCWJQKUSuhOHwzHKu2zQF8m2euuyaKk59
VDWaKJXHL7Nxz9cJDdgJCBuQJ4SnqCjTMZbyeiBr95G61w8heSV91lrON0ccpvlI
JtVW/GGEqFxaagoTxPHRdTACS/qzRt1emeE1Oi0LeEDGV9QhN4lcui/wqF7AB6GV
M0L2H1hTH7+yFBuvroXOcJwRWzfrWKX5jkHMSlN4sJYzbPMCPbxEX8ah27ZOEzSk
sTR5mpxjlONJ99C7W248eDxWeiSJF5ZEIRi/44fX2HVtqo3VtOV/1n9sZkMfh9VR
cgWfcsON/ig7IK7i9Fz9OOatKBXBUQbYhTfClnleK0A+3wYU/LDmtauvv2irj7/5
arrcID36HU4bj4EBIQ9Q/FUjJbkoZtOX/91BHfAMwdIBxicdyYCbvrvkrYCQFFEP
cor4ByJwgR7WQpx8IlGFLJAN1opAoO+c+vNvJNZ1FZq2aTbrrnLd2SlLe91CubGG
/RSZhPtwINcZeWLWd+FSPHCcGYjQE4z5pI4Y+fu1sCbNcIGVJmmqRJOCoyE7xn4H
rRlnm8OerMpldkc63MQ8adgU1vxqOD+x8R8s80hafOmKuaRY5Nsql+vx0utlrti+
rJApF9+zrDIH4Qy0861wIYwtySk0bSpWcgMCwjYhaoxkeJWEFMr7hIQLKzqjDD1t
IXj0ZpGz+OXITMvFcZreH/pVTmrM3462oP7bkR6PfosdfbaQE6WpHVQBAlbsJXZK
6oEE43IR9S8MjEf+Mof9vtXXIT8FnHUYn2rB6UQV65EB3zeNJsc2dh7pm5KuIvFN
6KmFMHnXTJOoTayQh6o5zGoNtWxX3BN+zHfPIAKW603b/KO+zGkZHH3rPxtMUoj1
Qm/NaNcR0p5oVu/w8MyCgj1UR4h5otfiD13AAjsJREqS4NJ8/63Rk9+gUZnobXQo
xdWKWUU722krOBgclzHug53MylEw5Vso8VyizeFPtaqueGCzxr1CHaQ4KMib/ljq
pRPP8WVLrWvGDQeEWjBrPWneQQ4Oubqs5gCJX4rGERrYxJu9O5y1clQ61lrCCAHT
KUF2g8hvrWVlb9TvWQVBEh4a8THZPy3WFSx+bhgrqxyFgJVDlXTUPoJiHn0szQ7r
YWJKh1JD7BB4CiViS8+rqA4BEz8OWEzy9o5V6Hgrl2yjr58g9EmLdZvsSUdkvoSo
pmpCg667CkV/l757zSfCKvvmuCVMgwDJsecd3F6oCcwFm65f1He3lCAQqOyadP81
5Mti+kOF+8iaBeymPmCydLYmh8lRm7daI7JIZeWog8TBNBiPwM/AgnOkALPzBkUp
4gkYpl2KnJT9v4VR/1uwuP+6yNH9vAHB0kFuyV8oWQP0VPLZYIphqAYW7iEDiFo8
zf/SDZxP1JTxP/+FRt5awJmamdkEOBWKIgxTxcUgTE1B0AQD0GDi4o350e60sXkH
5xjeM6l1BecdKdtKsWcUWg/TGYPenuIYpBRTcJnfQjdF7jkg1W0aaU2C6iJLIexS
hNPhG3drhhw45xOnZtnYGKBZKRBhJe2bCVz7R8gVOuST0OQodZrLxDd3M+Fxnd9C
d5K6+2bjnSYhctKwDR4tlAMlvNUPFoE4K2ZGPX7dLZCpI9ljkxHBLiFmu/FYW8cK
pfOySk30z9S5mzkLOXHRROgTv4GjNBcnwJh8yrpReC5q4Vv674aIy4Wf8NW+93HV
I27t7ZTyl3l7bJyme//CQFJTYVhz9REV9rrJggO+/xVUJReHQs0RYL+cRQcVJ5Y4
qpGSGQ/rr9Gs5Txlos8ipdIqC6Pyn28LxhyMm/FUMwG8nkogzifJZNmG4R1XDo6Q
vaLYL29pYq4A88+0FFI5Mripiyy2KhuWUlbbvulzQ5GMEfk/fjeFIF3pCTTfBdZn
57Uuf4zpqHV63R7Gv9FiV+UIQM8zwsNwjRiOdjBrHOgonVsL5WUaRFic3AdPaRIy
xc8sB/kD6Rd3CjF+dORGcMp1wzAD5xfuxfBMhV1B3Quhmon3U0OO+y6SYnRsho1i
pPVVTcs1x1aNgT7zFIR1cfIs2yIQEyjBWRRmJY6mpWFXWPdTCEKfPmkhjTa1vm9k
DaEl1VrVXcFRvp8+JL/2VEl6WtCFCzPq502Mz+w17BJc+VBfJKmkwMRJ+pgM4C2g
zPLIn8Kn6agY3Ek5tnYWIw==
`protect end_protected