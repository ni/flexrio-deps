`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1872 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/aWAU50mVQMRYzJ8ifGqH3qUjzMlXtPPhHWFffjQ3qjY
nAuxFgoyMpN5LeEL71WmwZd+xW4yAK36siNt/jGGEWJN4NFqshxCiUKj5UTyvWRD
tN9G4fXpc7jHp0pFYIp+K74QIpTrAHpwlFXLnKZ6Kd+AVayN4dezPzyz75PsBjiz
kZFpPx5ZGxdqr6nodKZbUGybphZydDHDTWmJChU9c8eQgTmNBpODoo7NhvFcmeQL
F+pieVh76mAks2SfyVgyBbzniQ317ZBQ5Lnce4ewzXklih2S62XQmx0TEsn88ai5
JfKUjDYys4EI0IymQp5J/WAvthyhu3hcQNCJjCFbby6OKzOXDoaSoRPGRL161htv
8BoYe6tkYtfETAFDYYGh7u0AaIgaF7VuSboHXHa4XksiWg4RndXoGP+RQLHR78iT
DbBeolorZYl5Fc/2CPSYmbeIxh1/k40Al5nwsMw6zF+T16sPNciGBU1YRr10sRon
AdI2gVY25pa92RdQ/Hfs94xzlNcWrk2pSzx+WfjYFJK1H3sVPX9iy9w8phiRfxq0
IFg3K5hM8N6r3zi2uTtHhhs5IupnkzK/Guzd8R/SYJ/yTHDZgIPuMamfDTmd8QqF
L9rai65NtcKNmONuc1mmGpbkVsyek8gpoM8otQqefYrFeBwrKS7+gGqF4qcbSWcB
2jv70gMDlbT2ay0efll6RU5rUvSMgxKLa1ifYXAiLatfKtfK35ECGqPeR5JrBmvB
iXpltm4hFJmHfQhu9/KzWN2BhSXch+ddFf+Q/Hc6unjeh0l8DYARQIzxTMp+t5kK
+R0USbYUkpYuSuRIm7iWJwLnjmWUZ2bF+9sjqgLj9JdV+5w6fccEeksrZbuiOW8Q
zvL44SEZAR6vpBsqyfqkqCBkdzvn2WVE7cliBiexc+MjeVRzHEVezdBBoxE3iadQ
hCnZ4IdOJWXBz27/NebxRgSHSxT3kAJlTA5+GUox4Tf/EwNHbK5CCxEjePLytQPB
FdbHFZqRLmkterw9i2d9gzvVrU/yHLhgdYI0zm4F+B/Hv+KH0vTVnF2QqFwpDlvj
3GUTlCZ9kFSN+Y4VyFT2opqOr6M7IbQRhe1NEUS0XID29rCiw6dQeHYzHKcl7O2m
jzWNs1enXT9m/ikW4kcteldb/BQqyr54vcJ/wTefl/Hap6jKSSWyMrgezq4bHhfO
gBB4A5iJYfrI2acAFmR+aKDtAwp9brNgjop0MT2OnqUw9QnXqdh/ICeYNQ0c6Sbn
t3tOzRyypJXHAJCpMq5qYXcmZz2ZVhyEHyQOMDjpcM3m79fC47xvJg0YOz2oCYRq
jsuxGsoKa4Z/QeBa+TL+5Zqx5mCKS0i50/a3Nl0YjQyWjyZUisnyAbEP7O5VQR6e
nQYz+4dr4uI2jAJTYngam7cLe4r++iYCLOZD0l1Gbq9FJFeH4cHnxoal5VlwTdLv
ZVzPkHMudaJiccs2wkZA6Vjy0OW1GJoGhnSgo7wOTThzh3G/VbKhJMbvJrm/YEEh
HU5sL7YtabB+Pmo1TLchCPqKpuVIG+oVAjiPm5lu9vl5U+1SBXgWx4jy3HwJjZCf
nAWZWXi6umT9O335jsh+Qt1+IEGtfVrL7NxtQynh3Fj0iXcX7IeZe83XFTFb1uRe
znzxhI9QxXgyYOlqg59PJYlPA8Bmu5zDHDUMzJMS5MOAzqOLfkh6pyJznZgFAKRi
IaCy+zdGCxT+zy6BfoI6wrmXNxbvCcmHxPvFdu0nzjHRj8QIALFU5vKdOJ8xtYpP
+Qvv9WhqHpFQgYlPu2YPCAGhCI+sbS/+aOjIpk9S6HGvZ2QfT3bGuRXZPA1ixmvP
73UnzrGPM01jJ6l4h7ovIiNNuH8XChz+X99EYjHtAfP3v51+R40V94lToJvEppM6
UF5GItJBXBQrhPqvPdB1pmf4psV/255MnZ1ggGIhVW3290Se3AlQwfXQaqTXoY0Z
2eWP3dNV2MSmOFDVAMOeXoetfOWP1edm5iU7XL2Md+VmKTqbBXKSSnrbw+qyLQ5Q
3tJRXLvDLsWoXvbEDMjcELZq0Yhf24qMqvQaSDbcFfv82Ijuv58tiJuoO93BVK5S
vqOymSKFBH2GMH0qBik/kI7cvpVjn6lSyNkvlID5bS6/amtzvJn1nTYK9gxrDDup
t70WRWEmeHwGR8dHG77PrJPSJw3syAlYKpjnAOp96wnyXAj21yi77IYOrr2H064f
r1KoVvEAgAH9t7Mr9NH1Pwssm00/brtKBnGgTsuNba+1MB6fGM8zSe/eynTWciSo
5SNZQ5tGPFzYtlanpwTmmuvfZvMvc4dk5hS4JrVJoPRD7RbZw31r0x6qWQQGsAEQ
`protect end_protected