`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
VSXhFIuaIjCHh4QnXeHfrLb1srkhQA6YCB5viS0hqHJHzUk0ASGDHri8iTRi7PSx
9dMGtPshH94tfgg7GPbpuawQujzUqM8TjAf/1tjxhpd/cr+4Sp8UXY15g3hTBYgm
fGXnYvyZAaQyOWJKkWH0mbN49R9OPZPSVHqnJsvzv/ggw9/pTa8osuqPIgkzPr0W
1kQHruocfsx+/HM7oNz1Bbqh7ZpW60rwV/Fl3T8ci9PD3ChfuNGozstNs2nX21wK
PASR6t35SjBMJf1zeE5hHQMuknbma3J02K/nV5Cta2VaYELe5eyNpq1Rl444dcs0
Kp1RLW+JuJFlObPepOt6yrwln3Q1JjAji4SxkFeO95DbyzjRdZWIiKOgTE0ZaOS6
UnoJulSgIS1dvE9AkQB9u5RMaoWgBROIz65ipBH6tnM5wVGEX4XEpRjg2a1toF/5
FkhzqwLO7a+DxNjPVj0Uko6uS/2UUmldA58miSDfBLVEQ3LiukKB4ZWKiSYW3iCt
boNhKxck8di+lrslK85mAa5ZWH7Ktutm93D9VJWDhhDZnZMOMP18k89u9jXmEjcX
LLc31wtKIRYwdwwy0QgN7HJfJz4D0+WyQtYeuETo3kKfshzdY0aHUE9MRwTO7rjv
w9xZJm1/a3+nwSm6mL5bbFnnFBz59j2nE3YqAnBmJqRMuwi84bTr9qtUcbiJ1HrA
YxdYxWC11fktstvDdyp0FY467onnqXGNkkivlxHJeXlIY6Nf74wHtAPaUEkksHtx
ymVVdGXBFITw4+t8TRCHHL3GoMY/seDDJ5J3+hDcxalt8pv2a4RqdSRwbimVVXlX
8sMxGyNwFsoS3oid+UouTrNfOdvXKyyA0QMMPys7boYo1DiKz2D1q9KO25WBDDZn
8nYSb3L1KYPCsPGqFX4WYHfw4v1Ulx7aPCbPqhqQ0NS0/Zsr0Vr3pawjfRpG1suh
dphY9BgSdukTsF6Ot3/EhYudEU6ApBOsema4kBu1fBTENiFkUFx/Zb1Zvh9dOPpo
S6etypbslUvQIVdHZWDsOD9coqHd7OBBqepqdwOhy4pYE4f53AJ22BeEeGIzOq60
HIKbHje5ketjBMASe8yayjVBneyV5F7F8M4txvalDQfnyBOqm2wx+giO4rzsPztN
rzJIKmsCDKmbWkDXBZ3xvO356lFqiC9ldBxzJxZcvfhcb+TShrwRqp/oFiFd/oPr
vzEy3kqfGB8R3g7bo/1M0WOBDwChPy9CRqr1+ushPZPN/XS7SwNCYB0V6P4wg+hQ
zI6tv88ht1tvmxWcLdgejkcTHLLoYdluKv6FZFINMahmnvkscSOL6qdKiz80lbSw
5qO3o8r1ChBTOi/VrUmm0If6xC99F0OSvCpfrk7n3YnlFmO0bUWbebXWmHcenbeV
WofJqF1k633xYhfQE/RZLop/51ENtA4hQ4hdBDwf0/D3boRRMwLtERPv2FPIxxZT
rUIwQ/fqWzqtNpb/AIZ+Cf/dXn4qx+AHDu38ahmDY81873RGzcg1ofxh4yueSZ86
M6Mnpfe1xUafjVyNnW4S9Prh7Ge2F3d9g0nIb0b5YVI80Y1rxi9V7GToi/dG2wrj
iMQtRzrpcxwFVKrbtpMFQ0uDdrCFX2CcZ8stCKC4zA/xEUmeueWg6SWGZEi53pU0
kOXGPm1xkQJSO5cIAwWU46JSpSLmx6qc1MA77wW3W81V7ShAYVwnDPtjS6XX01Hd
CKCtmRTFunRI7tCvlvxwurqt2thB84b3/aAwIJr1eLFbwRK8YuZQbBe3g5AMs5Ul
mW5kPm0AqZ+fyR/0KiXHGorFOZ7YcFBsnLqzMi/J3fbBVdjpfob8WDFYRar/NZw0
EfIOgMBkKq6B75x0vssHGA7Lgqsdzd18Oem8p5htsDLqV47LOJcR3lvtlX42K7cP
Y8mkOaK6MGcJNnWclWixYCU7zhqM2M49fgHFdmCK4tyiaywqGQGvWU7vrw4yHsL3
X4pFOZ8Qxu6z61DP3Fj9NaU7keoQwkoL/DFxKqPJyQCVE1pYTSNFpRzRbjVKNQy9
NhMQJIxPgHEM5L9O0oeMVXFD4RukHLXsbeyj6ZLcZea8JmdZQ8QJxDtCDs4cNFax
jcZh9qvEWBGpUrqs83zULv6TUkM95uyqMZAq+N+a4cA2M9XQbfuVvQvQFt8sDTyW
roM/HJtWIv6PicAJMSQTlgkZfnoSJ7iPeiij9g5sCZMBznq467XXMostzeOz+rfg
CDObtj/EoDnx0Kozsy92F2sHPS4W8Hwjj2UJvh0W2+TEVCZCyNf5n0uKTCPcBayd
64p3hftVrOgd6jN1pEGMbDBetXfY4oHxIDSecL1H8abEs6KyYqMtK2crWq8nAlZN
CgnPtCIOxbNrR2PuMYWNFfjLTqg+8VgppPoezTnKqa0a33kwTO+V2SclL3nbaiZD
Hy/VtP7U0O8wVHz9O/vEG5TDXfkp9wDsAeEdmpB6+ZnyjdpVKt5J4/R2KWqz0nWJ
msMJ5aaYwiXDFOGJlQe3id55EzLOA9AWavECI++RCTUBrWRqI1tXDqn580YZEP1h
WZEonfIjcFEXn5XeU9IeoP4gYLeIzEW6zOSQ+wWjKHtDIIPDrzdH+x0aV2NrUFmR
iW0wpFngm1TSlYJYXvvNp43YH3Q3C6ct/kewxDKkcts=
`protect end_protected