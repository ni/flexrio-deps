`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
cXWo8LLcsQOjItIP6iyF0Gsc8hp1T4cunLRdRXz2u2A+RoKzG43RyUFA265u24Rf
E3nP+PDWaA6jjtNnEdoVaG0d9zbZdPekKAWXOQZxrj2Nh4/Er8cRU4WpSGKAMUzb
Tgh457HmYasjHF/AtyWzuODwYBnngUR26SanLVnp7wMaDaD32pnll2F6CHafLW10
Xn1RWhgMwM8eS/AaicGWYBA9iWEnodU8USzg9IzFEAinV3ULC+W3Cy2EcMtGqbDQ
Z3H+P8yAkPhI/gH5ad0dRmpSVdFLU6vT1WyxTCZKkZNUm4OAZ/nHM02eIpbA3LP4
xbjM1s7HdC/DfR3++hY1OQembbBoL3vu3oACyodg8w9GI+8/oeOOXE0aZRTvGMDu
JgL/e1E9jvTi1s7ef2a/g3t/7kciGce6zThtf2+xorUUPLuX4e7dX2bMGgXUzjuU
dgeNJllRZObjs7b/SDALJGqc9cLOGM1xylTNq+RC5ZEfkLQ+v9nQ5yiJyboLyQcs
OK0Y/vqqkrtcB8qdv4IRqyn61WIql+NkVjluK52YUNm1oIo7JSN8BSV8xzlk17Ty
rgzTWjkvzjYMxk4f/G/mfq1SZMK5NUeD/d8gkaJU1xgwl5AeIKu0yHj88glA5EwI
HntGQbKny+V8Cdp+ZVrWrUUlR2WuZNe+zV8XB2EPa234UWNacf6+js2usV9GeOWK
A+1E6dtdlB75WWcd5srhO7mJCiHgKLEjPaD2N2yt9ZnPCOMsDugER4OrpD2Uw3dk
gbdUw2qaiS2iZQMpjfiB7PLq7Hj1vq10dSRJL5+6WfpMNeyXoATEaMV/3FWu/a4S
7vJKfpqRAEcCfzHfraaBEsMPzIEzX346deRf3Pro/F12E55VA+kZHXrEiuy0kGjr
YQO4tSNtPQJn81wEN07R8rgQ3aWmh9YevwDFM4bZI1/SVWdS5yYacksCfwn/dI8i
fa/doLynmvrrO+kscERWi6jjw1vahSgn7cbEhKASV1AW41jyKPE57E/tTphJnnCc
f2B9mzLT5l9m1e+4g9GlQPd8yoeAv2kOa8j/qZC0nbRkvIIwKsfYsiDZUavvyHkY
7AX1NaipUbFnDxkH6otEy6lOgyDhoWH+daZsCgfOQzZtkiQb6aH6ry6PX1oBs3hu
bLUBdMt1dC4suBN+vRji7B4GbWGjFw0kZHOe+vFNm1x+zOugXnS+LL01UW5p1RXf
YNeA1SsGUXhL9WjcZWtpBX45MicWBsIu0D1TzIvDpcYQ8Atk/hqetoED7t/yghwM
imoJbB+9XfhcnYeXH8iGZXuH/yiZajzijdNh+oLvuVM57WNPBOrPZbncluoYVEmz
3vJBedOnwoj2uP2rY/ZO+O17tCkCNtyQk8Y1D7DP6swK0trwy4OGG0qrpfPbspPg
nzxynYXzR2Yj0BglZ2FEbvC857D8hofi4bk6EA8FLB0spuGT/NCCMfyYv6y72II3
0ckMSbyV5fPW9NpLd1XHMtDI0zyOibDm78qfJe+9IjtaiV3+re+ppFXTGwrfdmty
sqjkV8dPqAkuTUw1nIiGVvJVQExoTyTn4BNSMhUOs30nf1ULVQXM2tsryaGrdmWA
Ul691rHFbuk5PGa+sbDEEeuJUIebDvrrv/nEILfMXZZ7OLHIbcrZRrSwKSWzELoz
eQWk7xJ07iyFjIrAsN7Bgww37qkxodzaMzek/7euZV7NUT98UlqvpShk7wOO4Dok
0VJBKR5LEx7yluewWcRc6TxXthOBkicVNgHVST1WEfPzaZpc53CKU+TPJFrB5Ghs
bYc3mNLL7YMmTCmNfhn3RCOaQS6xB7lL52VCnX2e6j9Ka+shGMisySsD5ySADyp1
tb6SUdKdvcMJSSj8sZwninUCgG7vg5HkUvQTnmxjHnY0ihS0A/dVo0vr96f7aF7f
+BDUX2693vIYylVlMrPAR5R5P9aVAa5D8IuuwMZolu80G789zgLN2tgbq0FpEgIC
oQI6QpDpLOglqPdSn3SXa0P5StKQBsk0iuUBJ81QS55WdErZDa9DgEfnRP8AfJ5Y
GUjRl4EErQDDZF0SbsUisobbjY6nnTH3QeGjx2QEnYKKA5tlHWQ9MSTmcyn7YK9U
nC/yYG5nmTEWHQ8iL5DK3rywQWYluctNT3+0wNpZDSTGCcnY71hW8qbPyRrvs/RB
s67GyaZ7XImCsE2YsDoi6NVSOnZ/AIB/FOIWyq4+YNFaEHEL6VQ29hGpRThhKi/o
nRR0QIwNfud7+NOhmUhNspnn5R8w+9pq/L+8AmnHo00edkieew4m54C+oNVR94Tb
VBulSuQTvwxMmd2bzGMpefUxZUWs4KRzcOQoTgfutCT5X/1bYW5AI9Z6+nFAz0yA
cHEwX7O2ZaesMVuIvI/IIGnprVMO0/5w725CfrUpfK5VVr+1mGJkIfVKi/tuvKlD
0kJf6Yv7JVPfG8OvOrkwHzVjanTylVRQ/DW/iIKhcfPw+Gt46xrf9CKgbuWVDJ/8
Elbv3i1eS52S4DGG3424B03Gfsv/eAPf1rfAZy14lQmJdQO2iiB4xGdQVYyWXILt
bgndlXedRWFIYfDhdnrMGpJNwHSx8MgeNFiUoJqGM2i2p4Heen3x7aH9T0gT+AKg
x9OQRlUoEK3wxrL2PY4Fs9k54EX5V9C14YsXU1/inB2L0nIVE7fNkWxqpKWsxDG+
Gs4S9yHFPY6vSNEL85X8grqGX6Lqp+6gBjuJDLC48n69MuOWuD80wtzMNaBSM8cq
dyIEdHumTTiiiTB2/g1uCaqS/yrrW+SCA6J7lXYTeBOhajadUBxoLQPHu3z4lgpJ
/HCjDFGelZ9RhjDRn6xNZnLRIjnbadrfWltVl5fkm6eTTshNK3LjOUjSTL1aNVur
GigyYcRaOYxiLSBzZtNZ2e6AM3+7BoLDHZfyacART5/WY4HVypHC811HL87m8C3X
bl+ZEXP7WwmqZjaD2scbr3jq1wX2h8Dt2XfUNc/etyDZLhNHKXR0p5ldnsrhBZk/
AZ2Qaa6ha33qXuluF4MXfKWHJofbNC2QqSpl5tCxMzrMEA1z7CjwvnKC5X0jkVNZ
S9i6UDhRAmi1xzQeKzCY63xZsfmW19Ba6qF/3nrm6h3YxkGwYVpkfJ3ohi+KMW/T
MRxGCyZ/toTeteTZZAH1ogzwEhlwZgkVwEET8OjERYCj5gztXyqpVEnkcUDSXmch
vNjCovh0pCfkPD5vbRBZ5mC/wJXvJh9ILY4goQzS/6ixiPbpLMmPN44ZNdrjwxLB
KIkAKl0x5SXajmke68D01XliKRGhFygypzfpUkkgJmGr8aAq0HGl5LRHbbUyH5gi
FjujphJNduXFj9VvyuvT2oGHR2ZqEsEeJwUXPhoRjPjDL+W3DB2rP4OMMxHfQd87
EcyeGBvW0+XaltmkxHGQaKEGuev65U0sHCwgGFy3h4Ob2PHEUKpqOX1xkWOlMJy2
vIqWXVC9wBefSnqbHAUMDql49LIHaeKjdw33ashlm+7vhn+pErZ6Kn4IfiRZTX5f
i2ei/ZFuOnxNFJZ+Y0Hv6VUeHjUhYnd3RgAduhOtDw2D//5q5Eej0hX8VVClckfS
ULzhXoq1zd7zJsr3/NFd4Whoud9hvGoTJNv001Cs+rA7dmckJbRZNwjXaLubZzQS
2Rm/WfK1i58Xc59fKNxpQhzpypUHAQ4vDobI+NoUA2QlSQkwEqbzxoHFcdWzTc8G
JJ/3s+8ADNrxrG6oVc1MNPtRfPuRYPIHvNX4UyZao0wK0pozXPTknBPsurzn/MHX
TMKgIBIvdamH56qr6ingKO2ZBmW66aSdCgbUCLg0TWKKgZXGfYaDK2J23X40C1SC
3+hHv/FzQ0KjHLJgrp6obtJEzyKhBv0bKKEq5HkHeGdlseB4NsGdLsOtoSslF5aA
7NT5Lv7Bk674BH8OsohwA2uwUWpAr/BjzZwpRVy/M+KW6LwrzyNxmU80OrlfOA4M
LkZoGOoSiPIbsoaX3dttfmAeqOTcL0qBHiZMNo8IhLJJJCJ79jGxx/0QQrBxCMep
tqklVRVxguVEjjsnZcLukYmEnbcFk1ml0TWgfJUk2+At7TubdhWPzt4l7SK/f1Bf
Dj1duKKQZ+DtfHQG33BIYvFXpycWEcGaOyux9e3UG2wObeLePc7Vs6yw6d49odUN
pHN0PRKbWY2NFepzHoFy6b28GgWT9341eHAyFbaaplhoiYvs5LH9c96HBbKbER7Y
7JxQj/AxGXyytS6WuBvXSOVgAxwBKOIGlYM+lC1bsIDRl3DxfOMdSLnDkH5ytvY4
fVDltbJGTN5s5hV5j5Q8lP0ixqEz34kPDTTdhSijd0Gw0Jw8f4JLT9KAF8NFugdT
diztaY/0pc92ib89gRyCUJn8OUl4yUyPGKN8U3e+1fWJ8W+4ZTgy7gxmLqWQdMxZ
NmsuCoiDTqrTPrBCaIks+aEfu+h35x8cD8bEO0ehXW3/HQBVenGsFqEvjiHkk/g3
ZcZAYqPQjIAw15AcoZ2YQXHmG38e/wwwn0LfVkRMup27DDMvhiZdlszmsJAkM7NZ
g29HDs6+TXUYKpNZEA/dM1Src5GwD0ge/Wa4LrUibwQusDX7viom7+Dnrtv7Z83Z
s7KzzKtSrxL4T415VQvUxnE3cOgRpJDx0cBMOh/fClhAErVv15tagCwk4U9CW9u4
1PAmInlTrdA1A/k4AOHz0VtGHtvognSnFRNm65O+wgLusoWU8sUQ2H9FDgA4xnsl
Vc8nOGdPOa7vKpKl424ivfzgHRs+F4BRGlWM78Sb62QPFp7cwpW75rZUwuCc5jAp
2fWY5+v6FLyTqwqOShYivBmj8fTWnS1y/ax5bMLc57U2n02S5JBCvgxb26s4KQgG
zEOsvK3dTnJb9LBIu4OKqFvUyPuSoXmidv+XPb/fdPO0sf2lk05OijdBpa7zlkcA
c+PxDNSY2yyRGQ81QuXCzV8z2HKcgnn+dDrcqy9WAVq/edantyZZAUMQaHgRdRfM
7NfS2mw89LfDopJDSjSFEh5u2y6qZo+DodxFfAoS0BnSJd8mz/nvcSDUlhq9/2S+
nOrKLVotvei3BceEZy4iNl8iWDCcGFqQ+i3qEpzuant5ZGng1APFE3kT0mugniYl
k/B9NqEo22qc3oOsjHzi+tU7tPXovlDUQRJI/cz9xi9cjRpbYQ4Rw9H2VmnNRS/Z
r45nWMGd5p19EFIaccYjMdPf2JXAGV6q7UtGerwF45I/TeNsPuooa1JSYFBeJLE7
WBR/U6JcMkqXTr5WQZaYvoqkl9oI70unqfn5fe5N5Qq0Esm5HCj+GJEBK16LSmkO
5YJ4GEfEoox9sWy23Gnq5y0ag4Flvr/rYaHcpFcPvpFtbQBrxqtz0HdAgWD9ms1s
PRGv3k6zw0yjglGIPF/+XiB/vZZ4rE9YY7pkR8VvQzcHV5jEJI1GdLhRR1UCHTUF
LesSn7hjMiJ+hszWdajPEF/0V9ndY1I5fIqD8CjhAIz3U3NPMV5dst/Qlvfaj4bD
1UOPdpi+7XsllQSDRWVM+z2rZcMkyQYCmlHhGw69O39Bz+PKyWawVlub3rjTGw0q
0KHG86zIdfJKI1jkabyk8PQqGBwJ3YRRCWpG0O+qQRNIy6GV5Sojl5bM45+tiYEQ
o4uHwV/+RAEVLJxonjeLrNLcuv0c92ZJas0ghq3H+EIXnIBSIZBr2Z3hBZb37jZY
MsPh/fSg2z/8YGZuwjYFE0qS6J7G47IKPGr6+xlBEZtjypM/kJWOu37ZsZq1mYLK
EC4XOguO+50YvbOeeKzqyX0eaxFqApzsxs2c72viHbEX44czv/3BZTdqwcrhbwBf
jTu4VaNl5k2Oge0EWq+3luNqJFWPFhNnLJ3ixZk5A0y5WjWd+BxbbZaja1OljI0M
KfFLHxiLshUAcZgk2g34w81fC7MM1+5pIpPDY8KNoJAHYZFPZaVfGEXrZNu68UhG
hYNZrScF7AVKEParMS2JQsnQABiD3a+VsG55n78/xzgjJam7Bg9KMCKu/2U6ckmD
hfIQ++sXTqWUGZV5/BBB7glaWTpdCmuIyjCIbW9u1uYCfxNz8n2PSsBHYwMc5TQ6
+fsHR8daJSirO2ZB6qB2GODZro3CAWDbozCtd04bdyZmP/jdEkYrYNhkoWZzt9Kc
kg7BzgTvGH3XHAW9G7glE7m3+H6tpTtByprxSCOZJcjZiTsK9GSkmHvFdPEq1N5d
4HpjRm8ZOwf0Ms4+SooHpdHTAPfh3IWSGfljFhtV+UlM5hcQJ+4gTMXLEp3Sn9W+
604znvms+fAUrd8WMlRp5+ZiDeNPlWrQPSUX1Om0ewr6k3DGz0t9V0hsiQZgj4Mx
+HeA/zut0FDP4z3EmNEVup4iFlbk6O8bIZEF2azb0FsZKQDQeJexzJsV2B3YqhLK
L92sEi988hXldsuSmNyr/69RMnEPU4En7oaZY2H4Cjc/jAJ6hubqX9/WZ+kb1duD
/Jp7EE5JP6+8c0kTTiCLe7jrEpjdF3o12BddWLzfcTb224MAEEE9OLsD5St14QUh
5R2dIeReJeZ4sRyfyKjFkZXB3ZU5AKtDOCYYrxGrwLvRRb3FYhSIwnPDxQtgbsrz
x/22uzuRMc7RRm1/qDdwIBOnnAm/SngSeS5A3TZqfz6O3LyNXtpyW9pKnp08RPlV
g9TTYDu/jXwhNiMaZc4/5MBjNDeF7c+C7TOzAje85h5FXNNR6hnyIoeNF3C/v2dZ
SeRELR9+RIGI5LRjKr3kq5EJ+++7T9EWyjovy/8Ig5uJn1kDlWf01BsRcz60HjdY
9yvSUGx7p5+z0jRKo2rUU5s4wf7YM2mu7HQ/bjO87ubsE4Do6/mIxUYvb5EgpQwj
q6gC2V6O3o4dtbYbgrxmW01ZbjGDTaava7gm0bX+ic479jdzUIAJvZN0FjRWe6RS
LkJG5dblB4oSQTu5OLflzgZ5Ic0g6v6/cp+haGO7KkNL1TZHGNOxwWvZXRfkMyhX
o6+D6+cPUrtguaxQITi+kBCg7cmdmGhLKmS+9ZYMy462X480UM7Hz3bsZd8ED0tz
9QdnzJEv7vmWClj4/4C6yxQcXRlrXZR8dg46dx/K3tKxuRV2ZTDjuUUE2PokeFpK
KDORdMMRecatfOTLM5isAvBLl3j2u8Ls1fLrOggB6np+0ckxtzPDcCXsLTljm0R6
DtwLEXEqGZJIJifZ2uNEBN6iGJUbZuVZAIdcwNzR/uPEW46RqOqIhrBtoaVry5Ju
aad64wmGb8b8XnU7Ormm+GRpqDiBb+vPQa+rTw2rI34FC/3NqJ3p0t7VBxATQUFB
v5MIcW3SkUfNb4igtnqZ19ReYWzZ4XS9501X4weCYngFCnqda0jHfXloplaGKxzr
lSzVNUQUALttbeuyVlQ7xU+a9HMuzs1aNqmWNJjsbfdVLlb2BPNY19LPbBiJJ9Ny
XSZdD+FRgaGqci45dRbWHDlglvLAvQcoqD72iAFSO1HZxeeub3S3WbIAEtNy57ja
k3OE4QyIO5pSPkh9I0tKqFWHcNtDvx2A3qWu4qzNwRg5dInyffk9oJfH39di//Kn
C7biK5YsbPtz+O3MwfFseVTGV7hgrc/WVQjhOGfvRu6Pq7lCd+Pe+BO6J08aoUzd
2IkJyWcx5qvYiR/ijA8k+nnqtomvVCvxT4dabUdCqpIEC6whAH3+sJ0TLTyXSPw6
ko3meyYXdIMaU+lT+0Keaim27hp63RcBqxxFMwwmJegPUM//YQ5um/7WibtFmnrC
TljgFfIlz/QlYS+9I4+ZaV09fsVlBguqgrE0HB7eQlKFm2scneQyTSVHts2aUnsF
yW9otCfak0xd+8gVt4oWrfSQDXrVZ4BZdNc2fmdDVa8drKkxscyMRga15IstWdpg
sPS+W2Uc6r7hIC0sTRDd2LDppKN0/HvDHzryU1TDR98gO1DbX/C3rEIMjtykvLDi
Q2fja8zkNDMvhhaJzGrUW34qDKrlpow8lHBw8X6p/LUYMlbVwT1TrmPwgTnvTSYu
dgK8U3sKBWqT6AwC/kX6tYUIaXbWbHdGRdHlKeXSbGOm1HO6JCQHIueI0YO15ZwT
j2qrvDeVNr/G6y7WboAhaZlwl4fWFeDXbwOM4ijQhumTzgReuu6pD3SgO/7kfTK1
XDlXc2MzOyU70kDu559UH4tKp9Y5gUGoqhrbvgNfWPLjt0xCViRLv8VSXIbvEef0
9HS3xLKvcKuqZxka9PnKkepsmUwZ1RDiSi0cCqhgoz1Dk8vVbd2tZaCSwnHdDo3B
VbdkL1DyaULPCLyREyienjjDAhgO0LIJIb0ysfaziDkbT0IhrklvpjusegHhsq6P
xiChgmQYXYLmzFY9YPR6pVR4toHarX2Pb3/FCySZYnYnmsLI5ft1k7wpvDlEuCcI
XyQQYL4xC7GecCjjnnT/QlwtAQtV7c+IbmSe8x0Z4+V0zjbdkrS58vBKYQVdH+hR
HBOo842gZ4zyx4bW9SaQLBy3IX324qtGeq8CfUFHXHpYKx71qy1ZyTA9wZFF1J/w
EeVtrUmqmc9Vnlp5b6xgVESJMI8lwYOiiynMJDtnEJAofVArJ5bP6k2wLOvMsM+M
bRGxw1frRzFKTsINokxFG7XYWPRVA2KPRqir/OLHYkplz0OnmsVfZQDndLTNNWK7
nK9imk1o1M9B8dZSMwrq/PRGrwsFHgxfAuqU9RPpc4axTumZgiLBe9ZJ183F2kSp
HHD9yZhNy8VkdHsCGj9/jYv2lImQaGiouFMvKgVyZdblvDjfEwDs0qvcCPJHS7T4
K0zj6gSIyXeNkzhNZ8v4Yv/E/8o96dRP+Zi1c4FShm1ejssqIV3aMseiRgEkrEdJ
ynEShGuafb81VJ3h11g8TqneUvOASt7wsftkiEY+dYZuOI08v5CA6q+rRYXp46zQ
qkxz2MZvlCZVMQ613VujwN4zeWi8BEEHsdbtQ9PNJegYcqj/fbRCWr71d21nPLi0
/91zxjeke4+KQqhfj5fe+cWSAwmG4QG8xHZe53dXaYentlTGKo6Oxnbs0Rt6/6JJ
ii/M8Qy6nPN7UbHNNSNPop6GjG3YjIhuqr1Q+k6gb4KYfwMCXWLffiElnWgPH4db
3ki+SkjiUMLiLROkp1mFL42R/zcQNvSOT/7Ze+qxEleGkUr529SN//9MbNxqxmm9
1hp5/FVcx6LRaESs3JpfpRFjyw6T0ZhJI3a7uMdsQCMHZmQMfW+lJ44UVx6UGWgh
yPmDJ5WgeLAiC0AsU4icdhpn1Hj1Lm/W3s4WtOR5FVY/XX+TEBpoh81wnNdUAaqu
LFzO9o9XE3Q3IvMcvLWbqvpmIxOYsJFjTJrFvRK/ja7qMck+AVTVwZ7hgSrJOOoI
CN/lQguTGs/QVz/PAsaCwvbaJYRzoVKbw9LDJsLWr3Mk2lprK23xiYuYa6zIbtuJ
zM0HSEDbkl2KYI5eCNbeuws1cvptRWvQLRKnGfuGV4kH1pzfKPMwR37te2feUmeT
c2g1FhxvJ+oFK0rS2TR0oyDP9bXS2TuDDpGoz6LJ+afbTTJsE5sSqjmXfbaWdv7b
Tn86aGUxpTmzpf3NIGE4ZiP433WJ3/aBZjiyKj/nHSzIGcJxMO3cloO8/1E6W+Ef
VKf+xqNxiRCsZ4thAkm++1NY4rFk4IWhYuO2uFe8hW5Oq4pZyGRM9gbTV1+cdywr
YIEc7UG9042GtTJoOvjM5ue+7UdyLp8hCNWTUKyvm67doJu+setqEWlFN0FEn1dO
sAbHGAMOKJN8mjXE5pK7Y1YakbvnIIDO5zdx/YIvOhII4YB96dYOgZFmNJtI4+Mg
q5B8mCSFWz3mzCkMiV16Uq/9zUZkHErbgX1fG4uV/yKA80jlklO00yfx2nTeDUC2
Fm2StzGvPP+QdD42cMybFKVDL8FAOaAuKQjiXWUJ7hR8tecp7algdb83hbFcCmIm
PxFZZX63a5S9MlSGQ6uXDllqZTxTHeQ/XuMqGMgK5y44pUrhdNGOLBVTph58jEi5
j9g43Ad8yg5gimu+rvibhQ6IAH39v/0XqTpn6NBY9DWpbuWBa1J0f9YeT5YWdpX/
xY2Q6+fdrJ2cfil1deP2WRX/1oIzdV4ar4PQFXrH08U5v2l7n7InrxpPr+gyoohF
OQdR9som/QVhQF0b2WTtpOPTF87e6GtbY7de1A/X03Y0cuADn8PacAPqzERJ4gSD
LEQ+D0Oqhjj8zWe8PMTR+IlAxVHRqaRbx0W6tQco0SjzJaE3kEmg+sFInpvFm0IH
iLiA2nSxC5iZTdRO4xQt0ayEZSOS0M4Zz0Tn7Ec9ZixQGn11Y6V2ooiJKOnY8sji
4wYiLGcQ9GJrSlw/gmFM5cO0RB/1yOqgvwG4qoIcxyiWstI7wk77zfaYcylniXt+
NQTCcuTSDCIizF4BHiWcl0LNVUFLpv2kap57lWEKNjwuV6Xlm4scWWiug3oI3EtJ
Qt6aoVBBV1WnjbXRtaKOlk+H98TuEMQ0P+Qd9PJK1z3GNx/RIEELC95dM4KGx9uH
k+SvBPMJUe6xf+G6bQav3CX1ZGgZxdeHbHAYn7tBgFGX007KrpGAWKVP+3hPDq87
b2oy31F9O3/xE/Bz1O4KhZsJ+p6gZTx4tIfmOO92TiHOvKaRarJsfmO3UfytLmEY
CckKg1PX8+L6z1uz/RUpjNfW+AsGcxiv+gUvY/CWnXJlCAhrIj9S+9WEEC+HCwVX
xcloWr+dvQfn6qFM+CcsPEhw4S19IiNeY+Q5tVgBtYMgBsdhF3Izkpfm1ODtdh5j
qF1XamkEU7imfzHuhAsZLl+bxRow2FT5K7EeHrOj0vDaeBQDB+KFXSLB25ffzbAk
sCALA6xpvd2E+kt9kK/8QCLmwm9VLHjonKqOuAlJvaRI4rBFFkRDCiFAlBlYpF8R
i96nv3ZWfqUdHmtZ89WZ2A5s/b/sy7JX5rbUX4IQvB+bh968X4HAGEBI8wOb2/Gb
DbThrQ1UdWx5D1xH/DJVGCFpfzMK/x9sCniM3ozd8vnaNw9vOu53Qi3YUHytZbzq
h4tfNlnP4UwDM+F1qrq68lnvMj/9rfMWnpty+Qce08YETbmdefnkC0VXtlRq3T7Q
MEj8GY8Jm/8YwozUVg5Xif///5KlnDvPsikT2E9ftWPV5iQUH9lbh5MhIix1+vn8
8ocMFl6c4nz//JouRPFPOsqLi9bXr2LJec1uj6G8ZGFuBNHQ7EmcF3lPvbyYWerE
NnPJr9SI8C403MCdIcBwddy4W7myfDWf0lR64ERPz4MkYmv5l7CIjS8Fapuk9Bmm
isHzZL9JCpiUNara+0LWZ9/aef1RRFUACcCyOMoWeD5MPYsRGfliUT0bIJVHc7XA
rHVI48KI5F+f5PbUNGzD4y+R7DSFLva/sK/VHK6ViijLy4AsiLWfiYfO7SZZo+H0
flsoTCQGpbWMyl9h7QsZRHPnOTjGjBOmZmpHcvCq2KG67+CM81P7LNZQ/CBLv0b9
i6+IW5e2NyKcRjq3Rr3TiCd3Kv4U+Yj4r1x1SGz05zGedA2M6bWaGekNncIBSvWD
7EP8PaCRApWnULNbegWXplfcNPQMFOL9BK2Hij4oZ5s+IIep2iTlAfxkjmEIHeSN
Fey8exs/C6V3djFvWrK/Pf3Jxk01O78QCzOxpH97pV+vZB2uDBh6nrL+4VJy6E5+
bw7v3KlQJeoVK0pd437vaBeUjRwVKXiyIDmFeYNSN7allGFykk6rTPGCGnKULgug
ARS4Erz/yzDDtkIrbNoPJ65LFznF+/hfmcwmabNY3DryWt/fapprzmaoHXYFxL68
Y5kTKRWV4v9fJp7mZtxH4L4XYVMgN6fBVPnjUxd+py3GntrcG++wP49p3V9UbAqS
3UfRDqgprnu51+yrmeErEU2MTc9+4TRtBHRwcQZHu/1iD1MeJgy9zQ9jbS56oWun
uQHvQuoraiMUnW9vKYHUts0JDeEHqmwUH9+dFytf4/jmLabJTSMUjaqjRS7rEGx3
v1SAlb1F1YLMjKn/oSAEitytTiaAzEFxd6UoUL1P88BQjHdoUD6hpR91mUpObuJy
h4UIYTGT1hgwgQMuLvXSxJQygGKjy0GvIs3b+FpPVBxnek6Xej8SDDf3vyDNeria
S3CtK0MK90CZuoTPtSwbwYKWkq8ltCd8yMRS8h4+r+eCAXPeowzWj5HvGeicWCVH
4dOWTbHTEsUTXzqwjgJUPtzaJPpu8m6bqV0vn9kZa1ONdGXuYevPamoYWjsWY+rH
N1F4AcAi0nI2WpdSHXDhyR/c0vcY42vm5u591UUMTxKVyNo2B1auw9U3bkfBb6MC
aSeDEmqEIy05zTuFGD+WPzFTmTKnHYnArd442xnKEqWKFNvTNXVAVFfRhqqYSPyT
rmi2ktKh+fpoT4d1XDAGl7T+TfoGrNFUHuxa3/ZEVfSGabXPZK0ylIWsAhj6Ookz
L1uqI8Mf1lYwul+wP3zw3NShanDYC0zo/AWSorDdaZWV72Rgu3VdatmA/WhV0rcI
ezJVip/gXhN2eFvTvXsx7OyVqx6Fd6vjZ2WK9UpWKrF/sR+XTm7/vd+90ys5zXgy
ht9NlBQ5X0UOqJEKjWwwXqHkgh3W1MvQzX6FdSbkcWAH2qlRzZmmVoJWZvfb+Zgh
AD6aKh1oRoig7I8L8tiFKKO47QL2RKAF80/Ao/6AH2EMCfWjKrrjyaaAzIpaaPEN
1gat6HHgS+kgG1Q6j6l4HD1ad/ksGTHkVaeOhSBgfFW/0w6fCc8dOHIlJWayD1X5
WrgAZqsbgXMT+eyP3YYqKvN5KL8njuAUH35+JMeLbVTYH4lfylS5G5pvge5R87hg
FG2ZneTNcUMw80hjtBZ7BjUZxyUVzLVmRbMSYSHGUIVmddwHxNrN3ZszLXWrQT7I
UHXDDVYdJ6UMyp0CPSkscp4/zl4Em9BQZHlltCd7zUAftyiudbSBbCHh3N2cj1AV
BZhGpLJKmo9p03cOCf3a9OEEoMLwAvbB0egmVyNQLMHuh8kg/qbLfPXp2CukQ+G3
L+nEjMpbm5qpSSLszDBEyWA5TH++sXTpC2ALsKOWQ+IrhcDnFCqz4QYH2EB2cKEV
E8RR64U8lHvTmnvtvWGKQkO4m9c15SKCO/Mp47DUgyXCP/nQ3iXgU7/TCq8Dw7Cr
z4fsGNwzqh3bwaA22PeUS1/gKwir18a4y471Noo/V8GvXMvI/Vk9BgO4t80pRjWP
af+nzrZr2lURIUdhncrDgZoCMvWj9DDfiJCme+jcczS6k4oxjbHRirjLik3Ad7e0
2AbQIiDU/hGL6sXaRelEoPd0XDqJrun9vF+LVb+uyr6XtuTzrZkXo+ca+tsyxEnt
EBdAjcOQq00M1QMcZZZ2IO3i2TE28pdopVNIwBtSOyPybQWHtjDwfqO9102zk0Zy
ztiWWzdzs8uJOcEE6cgblI2TG99OdG3i+F3k9xugLVBpcewihWIZk3jcRTyptc7K
iyYf+SDleRHpVoSOwP9gZJNZK+epfz/BPcNUe67c2VzjvTs44KpTUmb7NhlyzP2c
z9ZYN0bLpjMVFlO2xgAInF5T7EMFZEuGkDlVBXYlkApD0ETaPxP0F6RsumFRI+Sb
BsI1Wn2HMvGaFceHBf67f5h2MGjE+Z9Ia6MhSDLTQO5F3OjCFDXxKki+u6Lnj3Gn
UcKyRNPkXtP/r+QP/LRO9LerwDVVTnA/lN95mluVGnZDahQGguUj/d/gRUreRqu5
mCr0GaeXZJb7JHt3W2UxBUSeFct+Nx+I5WCkWyOts62V/Ai0jWNHLKRX5VmNUz5J
HDCKpn1eztpQqqKyvFUgj1QpVD6fkHZ1z0y1sPK7wKa6jOsruShQzEjiIZ/xm+De
Btlyf2Yy4Huab6Ltlax3xqWBvncUMoRYE1Kg8PlBfbwQkimbJpsezXhAU9n3G8kf
5nyaVEn/PtJe5RhzBy4yR8XOpgqSDONR85tk5ZlZXO75+2IWAyzYMvLnU4bgBqPG
DArMZgZ/5ggs7fRNbXQ7Px6eTHKErroDvoLNqa+Qm1ona9Ki7IRUfwSy92O9lJxJ
B3bL6Rx0X40lpBQpouIVR/PeM+U3cD+cTjehfNiPHVGN0rHTcFPf2pG/JyRvt/qH
cxgp25txhux9Gmqg0/1xvTRWoU8r3Rl5M6JXyqtbZ54NTou42BAs1db6fvf86OFI
Aje/4gDR5gk14k9w3fgzn6KuWAX7XILtUnLE5VN8zSOpw7H6F/j9YdB6eHJJ8wOl
eLOSuD6TiKul84f4+gTEw6xL0SQW17MdfsvJy6ENNrs6igBglTgaHRVLzSWyO4Pj
/LGqpGcNVGHm89K2Gp+EUoU7lsA3aA3JYN5XaSa5tHzQlIebQxKhHuGEFiZ+gqe+
qH5io2jKZK9B04dJT8pSGH2H3QNlYoUdCir7T0R3w6qtIrNTWvPgIBPeEfKQQTX9
5NZ/6PuWrgwDOwk58UNovTpo8WYz9vIz8Cs+KX+qXrDx0ZhxezOXotga6LIj8tpL
ZC2gR3jAa5WYqO2f62Yt0OBQzI9OnGraHVoTWxiyxKhcs9vRqYtSlfCfVxoiaC6s
nc5aanAtsU/i5t4Iv7jLIugtBXmIPFn1o4tGO1wRLuZahqs0iFJoW4iOcZYq6GCZ
bHpuI/TQsjUcLt+8436YET/+X2nrWdz2OHF8236lCB4JvrR4gX4nAOSiwE/8cXtZ
J5g3fLGDeyNRAO4yfuy4N4HkSGFPYAY1K0PGoa7FV8aFIdHEMmB+Ya6ISHkyYNpH
KVnxj0CU1rt6BFRDmVN5sWCPbWt/fy8h91J/DSqog6h6iKCwtX7NtFlphivP0zx2
EQPcgikNET4KlKl/h+zWZaTi987JOYEq62vI11mVz1FjQQGm2tnIA3Ps/6fcv7vm
fyLef0vtlT8iR6VFSXBguZynek6Utgj7o5wmbirniV3ucJ/y0DUIuMKQYsAfLWPF
KavPbbwdPYIuYUAyd8GPdGN+6VQWR4wG2NkiMDrGLDrgCRA1N7cctOi4Z6Yck2YZ
wGEIrB9U+7iNBzDjI+pVVOR95LI6EftwJxVIcnbNH3aH9VWp0jj5i8UNB0gRfuL0
tUs3qRJDCne9shE+qnR8Zd1nOiLd/VkP81RMOoWXanLn6hRWk1noSeNhKmxlzjgs
aQOxRec7A8Zsjlf8mmN316pcHvjFXXZ6V7bs1aRQdS3/JpkAJIvHVMEYufqt9PCW
CuZUBDso8l4JlscZKWSddvo4+vqu2J18Ys4RNoh7O8CmGjxH9vpDR2F+9qlg3gxu
LYgRaI4hmRTWUFKeE7hQAVxuaul/jYuOEJjpE9uEAD3znNiYv4ovBQhN1zXX8OtK
pszZ8smX2NaX2QNcIDdCrUWCcI4eVo5z+zB/r14wH9VJysOcUwFoE9EDI/zSW46B
hutBLQo3/qccxHenQZlf6XYRn/4t0LX0mtJkP5qaRN+Z628AkWhxKS8Gq4xn4/T9
U6BA0PIrSahXkgLdmoURUu6sciMvFQl8o/ZDV/QRCbtNjpa6oDx3IfusPCW+Ogsw
PTVGctq0vDQiIDeBJLgmq5QloNGDW1Epb4AdAEWhJEWBRWBQn5nf9u9Lkqm6WPXz
X87aRrwdubnFpaVvg39NCaPChCxlfHD+v66q987xZWTgN50NZhDLL462qUOn9MFy
0QPnwLKs6rWV42boJrUTtD9hOW3qHphhCPwjwfA8b9O885zN1/WHIm+eLH/0Xaaj
/o+QgWUz4JIW4BAjuF7L8aWnZ1knJ9Jiqe9tHgcmvK7bg/T9l/1GWBZVk5Eektls
JDvZYOMzmelyqlYzseT4Pk+LEvVQn8hkIX9UOQAYlb6sw99f9BE+jc0g1ewcv+3k
Q5UPrAlfu5Vx+NOArkr2sDXniQNGZMofkuPHMWAs6NyHZO4qF79n3/nffc3k9V8Q
gk/p0sluxW14nUv1OiPuxj+XJXIHTFuu/FWrXRZLTJBjMAJWn0DtKuXulLa601kI
c2fA0fUXNRlYVyAjSRYJ3sr11HNtOkfAEc3ADhvImMDeMCTL5NYSDiSzzC7QPKDt
L4xZtrlcXpXAosugo4h1rgPyzr3bfmbpzVcJwQxfZEurRC5/AtHRj5mgCr2Yx4wm
1pCaq0qKCsixLFWM5DoQi5d9wNEgttvLTfc8szC9qUpe7hsbMeKDDB4VtaI/Gu2d
tsA4ujJX2WFc6DTOfyuboNfvqD/sRxWxA+FS1y/s28DV2YWGEKYBi1vFch3EcBkZ
SybAKgEX4wiF6cxvXWhw7oqtS6uTqG7waJ09d+I2tqxWjaXZ21h6sB0yDuDQYwOj
GbHbkuk7hb0AW0vlYMPmSFMMvT3SVIoLjrRFHNGpAwS4HtO/AHrYxs65IdGh611Q
IT9JXHzrQsjpLbziZPJVBPqmp85BqgFp5OvBpp59GQHrFhABYsOq0YnOtFjf7NnV
yQk/Y95Awic1PwC81ll7InYEO9MEvSv6K3Pd43Ws0nbQWcdIV9Swy2+ry3suI5cE
skzNWCVAthaK3WIXeK6a65m1e0+95auAHgq6zfmILMSdHq3Z3tbZsc4QQviMcrtR
P90Y2Y1u6cz4ipswEhlFGd2KUb/QtUh4LMOztF9AgnCyMwwGl0eRhhphQ9akVPVH
jT0HRfR3M6xSTfqs1gcsepKK+g6a5kfx4+qQO5UQpmNKIUI8EzFIzkFiNaDvFXXR
8Bp4vtlfzra1dRt9iP2Qvg6zsEArptg/SayAeXmidFpnflQO2ww/nXze6WzZSg/E
XcIiK74ZRzpHmtPiR13LSdcN4zAcFRp/8P5tSrNC879cDJFno/qh0svp0O2uQYwR
eVVkCDQzvU9AYLwVgp9DBNC/lg/2Yzga5Mf8POeEgOoeQjF86sqtOzaWlXnVTJJH
ouHRm3p0feHPu11ho0t7P3jltwqi2VeOBYSR6NbaJJtlfySi1JZH1CX9IJlzUeWJ
Pg6S58o8EsRyDpGbCZvNSzvf0Ew/hAHgb77SAOqUwrMYNILwfPa9l4vWi3jOyEp6
DNQaaO0C9TPbOVjAbFU710Dh5BOwxg3yHX7/peZnPF9JzPVW9kB8+1WudDXZ/72Y
foAAwOGWaXQyYb5V1wU+HNSxSMlw3+YfGoMAttO6agKBdlDoV9cQUKoq4ld0HbIW
/Y6OI4IUhAdGw2uNmxIOxS2EtMKvNP6WM5c23HHOf6TqZ7JC6PaqbJvu8oyWybki
p+HmeNES1sqoc27p2kiATlZ3+gHKKiuFe9Q0y67i7nnL79oO+wUsjb9wB7KWV2HF
w4vdumTmbVShiu6Bk7ZYQswgbpG/CVzemPkTXWBRYpq7GTuzivQGnqRH1gGZJEYM
mNyvchh63avqQV3tZ7XtRayO3/sLHGem7UB0o2ndtNC4tSDTkk4XPZHoQQ3EH11n
PB+2txsxpv3TCkkEDgbax21g6zfl35fa3EeIl0kWMQb4LRi2q9Swz/QzUhL/O1en
x+qovFvJf+LgyFJWjqaxAcAt7iKhnYgiml9YMJbLZolsY9CQdwG61GHdNH4KaK3/
QnKXiciA/vn1XeGKcypz8suNKL7S26fZonxDeXXeyGuLyv9v+EEXINYmJi52C/CA
xeIRRpCFtfOP8gEgreTM+JkYJA4V9w37FalVdT7xANh0xz7pkZKTHjWlDfwfCORm
vIUYZCmtprKXc/dGZ2laHkD3tZfZntmhAVwPUSLVzUk3vnHtaB7xD8XIL8akkE+E
Gw4D2+F8Q3Gz7MemzEuhjud+R4Iy034u/T2fwfFKHjwVcZV9nwIPq1u615xkg49Z
HoVsq3oBrhPgyaqotYScaK/Fu2LluF74SxqN489uj3gvnDi8NiKdThys7an+7Sj7
xIYBubBQZoy0qPcOXg0ybvApbhi4xE2qrhIXKe2HA/1j7vahgxx/AJ5cy1lFfnfw
afsLGj1kAq1mND2i/4qwGl445nSnKRNAKMNGEyK4hVSSACaHIqYazOgBH0f9/bG+
Z+4UG5lz3rG63aDIn9B3s0ZLRCNMatMAf9LqJiVoMUF/L2Z/ojB6UYayBIac9zPc
lWpTdfpu8PZVeIKy2zAuFPsA74XdhKbCRU7ddqrmSb5YRiiwmtu4DXWCzjL9/RGR
iVGv/7OnoobmIuum4XMDiQujulQOwbf2jC1sYQCSWJ1zTzCfOIDCPlmSD4wI27mR
RQPnVFk4bRoSi02tqD5JCW+JuF0Z12jGGFgvVSbDGdYK2Wh4YBMoZpKYv6DfuaSv
c9oFLh7VQHtfPiySSaZ9tpOO6+1vRWJ/jobMr5yYI3tVL9AdHpHvx6FCd7RHEqOw
bQYBJ80JCt+cJjPjHRQal4Gi3Ib3RDkvkJ/k7Utt9elu4t0YYkB70OZf5LH5KIjg
wEnEfHM9N+cDTci4hEBEcyBrykcevdOtlNxepzoo8eaR3gPYACLHjNbiNTNyT7cB
kLohAZZ5QjvNDVQg9jhogRDvnabhDS3autf/H6m+jNyeCIqwjf5VxUpyAgX97RUV
41SAVQuAjebtAYOw4S4nDMWUzFvOZ54vsSNhxbC4RARn2H0DADnkd7jjsZGS4iYm
U2ehvfOE4OMkNxhqVWWhj31zV4ePTPXA4Y1ggFizisvCkdRDeJtm4+fgo6DFjmNZ
9FmBqZcRTlNramy+Jkf+E2a/wBkhEoeJMuQaGHpuW296VlxTXPANqtOpgxQaKJ0u
0hLbAAG/GFsmGFlcx994IjlSOEJvCGblmyC4eagDZ0XVbgFlhTSaWhCNU5L5uW8Q
9kLCjNcayNgsUZ4CF6QtJkZpXYQC1Nsy0/8E7AJ03M8yuy+4gy1WROZQIsiw1+65
Q2fF6RrTyUL4pADct9QIz9ne/4MEwUeB0HMZH0gKXt74dd+nDjzpa7kZ8FqCuaOQ
6FjKc+6lP8anwueoQgmnvNI+k3QmD+oT95pDzgvi/DTN6+vD2HSKFwcLZEDWTeJq
xOIjzUFtCx4IDvAGR6gFDiRaZYHSSBAGe0tJ/+EfqOxAOaDJu4OSX+vvZU7D371v
ZBifqVU1MSxv5FpHgcRZYvqEpQdduxKOAti0xADgCMySzr4zUEywPNWRMsLkOI0T
gTNtTv2Xn8NHTAZqxptnhrP7gtTIdXmwF1Ner6GwhJxT4uUW1+a/ifuHqLE/fpYf
4nWR2e7103H0TF2Dq7P+McurjXZwQ5YmrUKdTZAec8vXTcLPzDpVxHTzlk+7LAFx
mBihh4wCp2QVE4thlkOv2rgoOjwPOzZJsznaLwl61VrTTy1LsyB0cVJPnfoEZ4Bj
7rntacOVtBSyKHNNttK9X4ItK9gpwoL2L3kTkhhJbDM3lsX2iD0IH2TxmYUvgjQ/
aCf2grn5cD9FsapggoV4gt5GcjvDunGiKTK3I6ZL6ui1sPWuU0N9kiJV1xkv/cIe
df4nVGUXb1wYUSk37dRtW9HG+Oel5lHsGlmrq+oznLX5WDsRH0CDrQP8gBtvgzke
llhfsGDIWOcc37nvj5xxPG+zK/zfckhXwk53E6tFmfoX5X2wYpSI+zzSNAHqns7O
1WpxGtYLfrhd1zE1bd2NtkC1OiRVMUN48bayAZHFIiWBxu+3M7PBeQwh48KSgHX4
5V9QDSSdrssSH7VVv+vJxYHgFwXXArIC/b565lh/jQ+Q4FZm2SJCMl8sQ5wgfSzc
vdRFcy4z5PkupfveS/ljj++egh1DxsAA7r7Ob7IJFJuabX1DdZEzgCcWzCL2RXgv
XnHSTeuXFSfqYK4iR+lv09KMYKJ/iZU3Ol37z/nTdodS9qmdZNUlsCDJGNG5H8ZI
XMU11F2Z3GHAyXQzGAiQ4Fqh20y6Yws8eWXmtUsFuuY4U90XfZ9SpQjFxb/jU76i
MXGrWMUbkC7GgpnbBPGnZUy2M0MN5RmZkFH+QoW1FbJ4OmAAaKP2ZkgphqzLJd1A
wkXVOwLZDy9uph6eMX19aX6sRehVkKuRmZ2SiBUDk0EMpqCjqjtOwjl+4YcVYmum
qsLopW+YgGqozv97YfmviQgROnGbgEaKRztUwNFZC0e2LJw2TPjA2D0FWKf/zDZe
SRL1cA3C2shCanYat4xtR59hdtn3dWIeybXPVKSY8E5yDEp1uQbo47raTafui9Mg
WJWew8WXhvMeIzYnOxSWp847PV26jTI7L7VipNpn0lGS341r+6RhicDEubtnluxt
MGu+MwrUEH9WuH/ShKAuEYuk9JWCn3e8l1X4SUzJINI10tIoTyU2VokhWoisivsu
4UppSKpTArEFaOsueZUTzMJrogj9cZ7yyfW75bYw4DH0/ShwVM7orXYWKNrIHKjf
tVny05RVrebyDIWYDfeY18GnA7PRp8tUwoIr/t4uGtpH2T8dC/6nNQxSBpwwLC7d
14q6cqgygcdFbHzKv36PhhzsdY8A43fpbYDrjLamYKn3Gcwjm6tnGn8efxA1xoYj
MOqlc3Wg3liebvyYPZa0uINaOqCLQKK3dd1yV0+nhxh4EvkOz+qQRrmlmzEk/bRD
znn3vfKLPIts5Ty4xuvBjHhRAwKI+mCYRFFiJ/k9DhgptObUAknOlUYvnSkJQFqz
wUtUM4TgWtAU0d/9hR9eGzM1ONSGvaIzmxoNNg83z+EoJFr5F1M508hiEkVT4b59
r8drotkuoUZqvk7/wlN4B32ccENdjzbwFKwaufiOQw4Xe7p24di9JlrUz3oeZ9DE
2yTfahCFMSrse/17Rb4CsEy4APncipwYTGW5ezykp1ZeowadYuCIsWHjwThp8VrF
8r2eRVpF/QHCw50WVsB74i675LZm/CNHuklZ4oGhfIMk4JRLVmZpUqiscCuBpyAW
3LLHzErKAOt+KmlnWQYEXd09bMQs8++/hua+Go8VGMZYncpeE+sTf0C4OegtZMiO
I9F6Uy+4OUtd5Z0XmFAmRPfP2QhE4i0w7chJjN93+ssnOG7pXW8XJYOJjrO9IuMP
ydCfGmLR2FECg9D+ihPOyGu7oxN0eYbptfpPaCto2XVaXteLDn0oNm3mLztdzBdy
EHJGxflCVDpdyZZsO111/Wai+tono8JqYIOACkVAccP/C0nRYusL1SyeI9vJvzQq
JSYo1BLlOmjSzRtcdngDMRUn/7iqx3t42xKcqGSa55YgohD19xSBcj0OxaTQuL2I
RXnc4wyWqZAd1eVk8fja0/wab9uenHitZ19Cr8pqts1zVjtcTKnKMHT+d5rtN6QV
59XbMYuD4E5RbLkRVXaPJz/9tCdPhzI7wmCgjJWphzMJGV8PWw74wsbZ21Kjogx8
4seek4Frjobi4hPnB2t/3g3qyvQSmfLLstwOhc/7LI/s1AkRslQXmbMv9evXaw3V
Zl9zfgkLsBXpSE58vjbtB2S2tRpEPzBWiv/qX3yu9xFHhLh92IL0LN5G886EeA1h
ykDcxVd7F6I6Fi2oAqlII0+NH97gyEwQ28aIO4pvKS03sgL95f8AKaHOZ+Wp8g9i
qNxI85doJ6N867ReZ7bJWu4gIIMaHtM39P6mT7ZMY4yU04sV6Zqglp6cVcPcZvPZ
qAMMvWZvldrTuP8ttIAxTavlSS4hzTpaCcg6FXH003gGddOiADfYjcs4ZhvmCTt3
pcu9FIL6bPnRpAiv26r31LPJ7tazSJVFpd9NeKEQTwE2zVSHF0u6d+fbSN64AvIv
09rcgIFBi25h9NT1aIrgtx6qQFwWex4LrA/Tuzib/ax2JM4/HLqhNvGqUB/V3JaX
YJPZleHmX59tWtCxqhFU9X0sMwo5MeRnCwkCWHLTP6/cR0HXIkUUzIySgWg3GpnR
qvZY6v0Yy5OlOKKHfsePPC7pvcPzyE9+WNxqe4fh4Qr3uKYCmxNXJsRHI0+agMDC
Y59AazxyAstyAIREJ78l77lf6VF/cRado50wFMW7+2Dmi3ZTMvMKf25OBXVhNktb
rXZYVjAsKq838RW7LzAraFSwTZayvSN62fJzjvMUNvjshl1s0uNxRT4KOd7QOs/a
8wA63jM+OS5ME01Y/5USlidNBQB3NH3iAkkmQoejEleoctifMP6EEVyjl8Cv2xvc
mwM6VVNHTQ8vveq/DWUHfuoAOX3m6FMPzmugV3fG6P+3uZV9mj0pb4+fBUu8A96Z
Dz+ZCGACrxC/LzJ5j4P0keF29cRSlB5ngE7agMsK8oHlBcSsFkas91iXAxIh43sH
w9JrnNWPpYG9ky4f13HtOuuJZXIB+D8/8yvsJHoUDrUZWFJFPnkX1uOWAEaWLg19
b0pLj5mAXjQgDnI0NQrJz1KSIdmpWUmOzOYmyj8K4GFQPkiZoclfhSKXu+sbvmfj
K1ENlSoAAATL/0h+nrHrJfcuwk9OI+Iri0Lm5MzmbVQOR7HWbMxiGg2awNFLgpXK
8uXbOFp3D8DnDuxbsEVpRWHISMqNlb+AqU/9ltR4hkEuX05sNUA84Qy1OF5Cpj6J
3a5psT7FCePaoW4X/t9urcdItW4I5kHpv8f8++jMImhD+NA6Qbi9Hl15b9iEgtss
eZPaIpQu8cnh+COL/mXnIbta+/zrjhclMFhn4p2FyXzjeM2oi+9YrJ4QyMYrhiIM
8e+IudZKi6xMuCxdgitRxzQuBSgE5p+m7Gk9JHGVhePX8rXzqtj1/yqf7PBudXCC
/hLW7YEJ9NHDf8fnpe/NPCMS3231P4DUpwBKs8PPlVHSQKjAgfj+QMrRcFdVUq/N
h5JO56roKprkCoWsLRTx2NFjma5AZlpucjobRA5wR1IfGzGFtUM+y1A4KoDF99pN
gWu+dcZqDkGrGQA/B9vxOGeILCOp4yYp04fkg6z5eaX7gAmcp0lKOBFy6M6pe1nX
IbgqtpD7i07Rq1pM+GJXYDj9nJC3PZt+qmnTlL/1Zy3NgjdASP2KjmAouHW1Z6vL
3JzyUx3I569qKeKuYTF36r/Kuh7ymk4dfbLJ1UU9+Jjq6HOHmDGK1LRIoWrUr2vz
zWrkjn7VSrog/tEy9ErPkXL5joSCiRpRNBGzYBvxEjEP57oiTS43Js/jX2kqBFgy
10nrKx0JCb+qPnIPU0yjrOng/XlL05OGIdwt8K6G400jEN0NZfsMKTbO08UBcUm/
OGwzqH16HbWUaSpxKhWGMQXw9nzAuwpxjlj+C81UtLGIB2SIpeZyIuaW2P7SG4qM
I1+3RF6FfMdUvTw030xipwf70oTTR0CDID8U+VePlxD5cgj1G4gEhO91fSyYLMO+
0ofBvdCNx74pqZY3vpQSreny2UqG+9v2Ft72Jwq7DN2lJMpYsm+roIRS/3gHizP+
JXdl5RSdIveaL56P/DPlEGXwxwWe2goxrqV5NVI0/rJWjlWkgscaxvWlQz9BJXl6
No8IWtLAzJumHbXxQ2WJC91pAVpaODYbN5lZioaMS+ll6y9BMgR+g/A+wZQLZf4X
PlfJhFvu4Mh2c73z2ZZJTnEmIQ+3gaak2MB0AZz/dbgdTtsGEWnfnsz5M63rM2do
kCeacvkbKvthaRzDCwbOi/t0k4DLuWJkG2FzpKMzw2B4ZoDTNM/XsnknB24g12N6
nHxpxPsUQXUHf5GNoKfArWttaCg6XMNpRpVTb6mi09sVK7D58fQo9QBpqMu8zWRn
pZhj6CIp3tUKptL59WFT3zFDB7Jn7l/y1U96hUOwcnOWAqQsmYZ1lJQeqfNAOwrN
atKF1cJXDSoaEqwZ/DByqOkyvosEs4L0vnHYDx57Pe7nL5BDgTlepusn/WoE/S6M
QQfCUKGohBa7RFkCmReQ0eEB6QeoHAzJ91fqOhfmKzJwg4My5OT2tFbBf9b3Uw4Q
blMX9QjrrhzzCP0JdKFclsF6P0u+P6DPNedPMuR9vPHSw0OlxZjIzU9q1T9N6zoa
Qrjt349/nUNlflPHqLeDJLOoSVUEW2VCliCYP/gh4oY/1GWj8ZxU+vcfuOVUCYZM
xdU1OOivE/UqBmAh7Qcom1DMq2RlK+IJzk7xcZXh4T9kJd2twglxXFDqaIAjW07I
W6SapqfcnEb1JPQjdO8bIKRVORz13hZJ6pCuGz91gGWsdSrGdiRvwX2Uhr3y7qLQ
/QnZmoSP0ADQ/BrS7JPzpPWz8/++V/xJc9SrFwVKku8j0ZjB+qv59fZLxdwtqAeE
aLyDQ87O/GANrWNQcr/WIDqAep3k3AsbIJWe35yhYyvh7dZTSzwVis8u2MZ0X8rB
4rLfWSbo8pl74i7jv6S9G6qjD7s4O5eUE49n+3y6BNSRQBZBiz5wM/LXCu2y/4bU
fB7dTdrMRUEeMDgEEReuxpJISOddtu5Ps7VU39UDLTbiO+Bor0IbGZ9W5WutvdX4
hD1EA6KlMSYo+asiuU/HW5PEObxgOEctu0RQZVZ1TJw3iDhBtfiPY9MS4xuBhSHN
jGk3+Q4G1j+nxWAgD05nOMxd81dU/KhXBoRR00w542lW/6BpBxz8aig602oSBQ15
iHKqJViRwsjxOk/4dxcP64YEjy9BH6vt3ZVKifpLwaqLEDLaSgDJBrUvC6qB0ZuU
oYaGr/12MfcFcQDE/WQeCwj6/bfDoUp3ZH/eBvhFWSyDYWoKoCc51wR8/A9Wobm3
IKkKyCdmdgsieJaBkzvhNXvk5qZH+5oGLP+kOhp6N0mFLyJ6NlHsgfj+N5CqAdid
r3vuSR0RupxQMoBxxqgHANb+4IpOJaWIyC/SOSAbshFCg6jdP4iloszlX6VcBPvz
QdV9OW/jKot4xqKyF2Djdudkb4fooZDjA7KTxI3qHhp9z2RxX736FIH64YmP6nSN
C3XU9h6zt3d58HKjj1UaZhGHrk4SnYUCvfgg485pKoPIuw7HAa3KTnGRvh/D3NRx
dM/FED4/i02oELOQPLbSEu4wNy6vHoSq/R96vFd2iTiMvUaD2kX9GQYJ0IalMWKe
PBuCIrmd0YTX0rGjEXS4mfG0xGPM22HHLvzxShJUQn7wpvrwl4uAWfksbHJ2tg7H
dnN1qy3X6c6E697jZrZ2otZPAv4eABbk6ixMz6pkzNdzxzMQXI+04uVCTnAdaAet
S8IatXTOOFr4pGfy715JA++Ots5WRcbjsE9Cf8oJa7ISWV4U1BiJIYouaURqN16k
sWCNQBmEVNtrrtwrnyplS2nN+RohuHIq8anp9DDNT8BbCrNGzK0dpFkzujdwI/0y
NBl/mR6KWs8R/+BL2CAjY9MOMguMPOCohojvbNMS+21oLX0cSYhhM77bNjO0ZzTF
0szYSsSRAP6GeZffLffgm259z8aKCngKCaF7S1NOdaRXq2zwwhFhyPBqn4cCQ69l
XxjaOocRlqNx2GazpzArXnv5eYzCIXnNubkk+hO6t8XdXsv2qiws0IdzizbrsUuf
Pp6oAKmJRqvt12MulNWyQseFLuYO7tLfYBLZIlbLh/NzX1GYPAP4eh/pn6Qjdb86
HPOfPQW66AglKOhepqIGsnGUI60ChtdvEKj622qix10pJEM3uhhMhaD0pzZ7oBe5
nN/v15pmnlIoW9N7IjDVdfgzrW6Js5KVReoUU3mXZmNnzKvaptILc4rTaiIlAsel
7Ne+xIDRl47sgcfjSQYpn/nE3S5mFKkrnKuIpTXVdDhQJtphJ+gOCZv4cgbmDAK+
TPhI/m5kZlX1BE5RcZySSGO0KrWu9aSyJKpDo7xdJUhCdCSoeUJnIASdo81uZRQJ
a6cfKZrc5jpSwX8OcTXb4bwIWelegGoJeS1x5ZY8DnblL5M3Csr0HMMASNJZtHh2
XY3nSxNijcOCSLj8fgbbyIUXgVKZ2oI+16Dx6oUZoewd7aLySiMu8+k+inmcGYlt
1Ok9JrCuH3IgESK3kBO5UfRuUevouPK0YhvF2VMlDCN+Pn84vfYdWipxsR6qiHC6
b8dF9HOfjBhvSdN6xoRyYVpEzm40DhFTzAf8PdfoI2vkk5S3bhYAiDgH3kUAg0A6
8Kaa4RhfSsdxFHV+6Qp/X4RNFHXih7QITOLEcqnkUK7KNK4qllZBgXpx0TI2TTGx
8G3Z7GuGp65qVXkUgggx3T7zPkWE1mffpJj6SB++FHgK+SHESSq0UjowiWyAFmPV
/8lygqJXcvS5Yq6rGO91r2LK00wIQWCdGk2Ec1J7+NhxJMijDIhtU1agbOdi9N6W
rdUtqB56X5RDrByzRarC0wq72T7qbttjAVHMM2i1qf2QW1uUo7uAkvKAKhdqhKRW
eABhwp5zExpo40q36PCEbBImgr7Ot0DRZcyV9jcBwgCifgimHprOlXAsdIhFT/67
kb9Nd0ojiX2zkeAgh+XhIaLd5cqIE5RhQR5AzzekOzjwPx4abb+ouR2wGS0ze2F5
gUviiBsyNhCJzknTVvY88aCflR0d0oI1SAoj28tI7uig7OiONvpjaZpNUiXYeXVA
j6CFf5NxNoHtH8Bbp0BV4a0kFv/kDeyJoiWDu/nzVwSqQscAjqOxgxtak8lFtvnr
QjKr3QaLWbBK+iY1TlYsd3VakGGojiZJwbGRDITFUNxVhkUfujcz6cazBmMzcjmF
cFcfo+pXftVQSkKG3qU+K0RRL+n1RCUCcZJLeTgkVtMP89xSx6x3RFy+0U4Odoqj
0mW+NZV1hV4ob63AE0roHwo7J0y64XHGV9ssKINhywOwBHbV2xp3vD9eckEwc+rl
EFWm2Hx2xrCj4vNA7E8sGPO9u/9znnt2ip+EZfBCAFDuDAE5O8uhIq3JpzPTv0lD
Ucico5Co3LOJWyel4p+/QcTb5GMinOIFZi/SKsXUBkDlx7hk2jSjexCZ+8CboCdX
WkSieih0FD3jP1aAWTdDyh/iTl+AHs5xJliAhbJJQn5IgHUdae9Q5WKB/p/HG2Fk
sC1dn+fOWQs2UyP+oa/NSFWhwCo3c6b1zF902T0BBsOTSuUfNxq6Eyr87xNt3+JY
9zSqBVTi+KHTGBCFOXjd+Tif6rRzmTeTzn2JC0++WhE+DDUi9TOpbQgF4+buBZ6Y
wQxoSVPPCQ9H5lm26pd/L08bsnInDUZrjEClVGX7s1oYryooQ0MNgY8No/y/ImO7
s/q+s3WP56JOVAloA5EuVWD4Z9SilCeRNnvTDgwjhOeQQHpPdzeXlNc8UgaBOBOv
k8/oMqSN0Rtrb47tdhxDQk+G9xGx3tPfs1iRObMUNGSxJ2Dc+YqXztfT1vRmSDzd
mjJEEKKqUzEM9KhbfqGVEh3/Il5WVEGc9b6O4Fjmay0SigHzqZEAPDHm/QP1WOWG
hOcihXl0PbviJvnF7drLj0Rm+BhzSqYqzKPzvDwfR3xYOh5DJqhqiYc1gKHbyNrY
Ea+eJ6ZqBugig2bz89OtI18NBFSNEXA/9VBklNhSbpqRS4uYnlTR0kEgHEtuSCjW
3enSJ6+/pm5JAprg8dUgB32Viz6nvMCDuc8BRV4X05t1sUzY3fWqeoXE1jUEU7HG
6/ey+uUO9YvFS09faLNaY/r/wFI817A5aVakYREczBqKyvzP00QL0aYybDQ4weTy
/we9PcdMzC9zApq5KBq49EQhdIDRpMIFnZnS8ALSbBLp0dM0S6/RsULQYJdZg8wU
GvQjeLcvWQsIgAaYys63MoLq8npXwNm9n5Av3sFQF/3M3kI5wlV96jpOvj9ZsZ1K
ZeHCTxiPpmM7OJReUqjaRqvGMcEhfRlZe/UH6DK2S8JvFzXBEVb87uycSs18bq1F
M7gjbJOlf1fUGGTJvYmrGHuJVSK8PY0OxyjhXfFZ/5gbiBmI1zYKOZoCZ4d10LJa
z7KJ7nh1viojl1ZUGy4HWegRMljkgsT07J6ix26fzKwN5cLI6x/guk5z/UzEyEmU
e5tR7hMWH3LYGI08Ck8/K0vPL9T9ZYkHGUdrCyU2zNTS6E+qiaPDgqrdVxePhVTc
iC5XdTPKK4/cjd8dubpbXOEH8qYNu4z1XRCkvLvLQDYgaqUAMAwqgP78hcctwn9t
8b5S8ymhNzgz3wMBJwDcZfnWTP/8I2wfHwMlT5X0aMw+K6Fdu5oPdG9dqcxwul2w
1HSTHpuQyw3P0qy5hgDg4MS9LnTzs+W8FxfzesubXsS7bfkHrc3GOyjIcCfXsmXz
++AoZmEkcdLoIVLTO6doVsIDVa6/o/on1MzL/P1HxWY6fVxclifGUWVf2HLm4woy
H1+R1sa0VLNMq2pa4RzIFShTNLyMR5B2kPZwFPhb7eZ3FKLz0zp2/eNYR4FNsIWq
lqEP4mz6QHUVoe97XjKsEnISu8Nwsbnz+U4FilL0AJIc/CP8OI1zhWdFD2934mZd
Hj3V0460hAioB2Ue8JzqWawCIVt+VedwuWnOWOZz41hUXVH6B0RxHFC2I47iuoRW
ndQNFD9UOd+O79Iqo3Zu52vjC87DmeD/A7b6HlVKHTlSL5vEAgE1rmptp2IzSkqX
+PXK3FLh9MVgpDPXhswEUytdgyCLb06Y64go5eGpUB6aQVD5V6wqyj2ubd6TiB/5
Htvhe4KsjAgqKS7yQ59krfy9IjMFb/0HzBk7ISHQeSTQtpC9BH3zKBY8aLZxOp1y
ShCF+NwSsvzwgAFvk2AC3cduKs7+hSgRtPEnbZC4XIQmM0zdMCW81OXszR/NEmQK
OxfW+TS6xG/SORWrwPc/yDfbvNTb6x2GS2g+LYtKrrNPQew+4Tb3ShciiBByNdcr
513cy+ALNIkpT7cwOHRUjn/q4xuyJEPFRKP9aa0Dg6yAAhNnKDrMcn96UHmx5+/C
kgLbcCncrZkXYWafjzsmg42EuvdfcVjhKuK31sk1u/32iDhTtXJ62pM0wEj+4pCz
OqgKZnYimN2Bt3XLRvxCSNTI4buDCx3n9gMvV4PyUorANwfDNf4AS+As3PzxU2wa
i1VroHQ+bF0wQfaC0NYD1Ikuo8spTNaKx5zWqldtPxrH6U31vk0Ce1hjGSaD5g4w
GwFsmcrWoEfpyuM18I1D6jmuUKZrzPAFYqt2w4JzWUWJ3+eubuxPQC3Qp4yjPAPp
5m3bTYBttz9xM0ezTRx9BeisBFFiMq6sK9TzmdFzMeXPQyGjx8NcgVnE8uwz4YZE
LMYQsdZOQUMuD2DVDP0pps6Wk1PAZmYTYJ9hx0KbfzvOVWTxqvKaXHSjX36uRu9r
O43ELrIy03hb6MFjxPabNo323MMRY70By3bofRYtMAF4TL8pW58cKtRytbvt3Xni
/upqCoyujdH11Nt0RCE88EtDR3l4no3htv8UChsXUnhnv86nCKswmsrwYS6udeYi
Repww+G/QYVCk6JDsT+FmobDYyS4198/JpKYxVS/h8hNXPGIDIGfghV5Vqnarbdo
vUFQIa9R80XZt2nyUhGvlf6+Gjd+Mc8EIhL/YZlh9EI4z1pqw9CfDh1bwJTzzJrE
DIzAM3cKCmGTGxqolAahx1o6+rvZB9CQLOf5IsSvFJd5atAVYQBplf1cCDbZ7Jd4
9Epkvn1pbcAjQSulgUJZwkoUrE+TO6uQWPFgXP/Gdm7ydXro1IJpfv1ymN3T/WrJ
DBzaIcn8IulsIZ9CdtbmcQV+ulqLVWKbdE5GvADpZYX3GoRIOC7dELvkUB5+Hkci
RTPTbPNZ2W/+bVvbCcfTs5pRexLnw6BEvU1AkySuvmZb+LEe9QkghlE1oKrHjFrZ
x3MkqbH5/zadUVKUJIwCxHZ8V6JPtWzLeGV8YesYyIKiuxAFaV8uVIR5zOCbflqj
CJFXImeCWs/8i6vrhT5TQZ6fh1iXlOHbw7p7xckjxB8KEDLcNTnkPfhRIMCZB/0r
Z5P+ZcMJNyyFK+04OxQK6xF94ZPDngbmf1UgOLCyhUthGcartBXwQCsE1yUHKme2
1u+2NtHokUspnscC5WBo1gIUfoqoFG2+liPuHEP/ReE7TqOLvAh5GupvgIxL6Axz
hPyIIWTjoPmwzNSUBbmsgZOtBqsbpy9ZoCyMpSsaobZLBbeD8eGrPr5oEH5aglyW
pvZ8SlXJOo4u64leS3BGfd1fJh55FnobxWrtPDPK968IBhGuhBRCe/ZGFFq87Wto
vj6AMt1FCkxtwT9mehnJDqWxnAQRUsQjhpDgC8+isNG1PHzqyO0X5DozOc8JozmJ
xg0kd5UWuyy5kxFxfJBukXTc0n8sGjq/voOzAsSkYo4H+jTMqaSMu+ygiecf3aKI
nwUXfHOlVyxmnU4e2md259V1p039q2JWX3o5kIQ4QRdgeBM9P/UrfXZ66B9GsKML
h2j8LZk9SJA0lr4n5wEFRyTiT+swqKebVbx+wCF5iq9qiptQkx6JFe2tKJtcCEV6
tCf9XD9EhZYFPu/OnnTrH+J9ZLP1WzVvSo0r0dFrhEWV/fu5Z+nAIIF1CvXi6o87
X/KYPRWmbeYeNZWc0fdnkiPTEu05XU8KlmyusZAs1t5DUoJQn791e8++nDDe0Psm
5DfIpNyhj/EUQJqdjRwN013SFJg4khnISKyqCYpEb9IsfaSJq3vM9d8eeEUfDYwE
AQSJFrQKmimQpGeIp1CySruPt+0ZPOsNaAS3bEL4k6d7YhYw0qOCkbeEu9OSpyPn
EIQWm2B3riFhxXUpTlI/WB1JHDIjvpNFV2NdTyIxGfwBpy8CPPmqk5bOhplzLReM
DQzx5Owd3KyAT99Xlw1xiYjDv5qvZHMNLXPwO3BsyB5+hicP3CQrQwtRRBQa/rJd
8rshxsWFimseqTLkDkzFN7mLJFm5ac0GvfdIyB16uQbmzf6g4LWO+TCQ5it11glA
0nV98zoelNdjMyhRPpoyk6krEz4m5Y+EGBqjx+kth4ZwByoyz3MiU/9OcUSW+8ta
OwQ4p2lX4AviFkhweaPU2b1dGx3b2B31q8CB5Ce76hUVxaQGUWflvg4qU4DlKPdL
hgth+Iz8zQp1y4DOMnaenI+KjJK0aTXsMvx/yxhAtupUcQcYAPRmjkpQOzYp34Or
ocujsDubxMPGdLRwUG7jM7oaJ6ufKGLBfelDQRXw3KymTTKVIRZNluM0K13y7k+3
nfQiyaJWbBbWa4ciJeInlAOCpHJ7E8XZdfkiH+6iE3h30kXfdn50UwMWTJDPy5SB
S1+QsLwrqdTdNmicP5kXfuTA6/4tuutB0ixIDCSMA1/RBASMGcQvhy67xne+NXla
9tLEku4Ik+yOUxSKZ0bqq8RQ2zDxEclSGsFA3PkmOQB+fclqDgABB3MKYTdP3MOp
ay8QuRZTeVXx1r0SUBowhbnTeVX0mb58mHdkhov7ShF7Byan1cfLgCvR8n5JLOBb
snuUY/mwPDOXRz3uvmHS5pQcHM+u9Ebh4tCfV8EPiIKHtJG77SNPNUXreKHw0l8/
emHkMlAEIirjIaTFgfZgwXVA9YXpnwB5QFBLMhl4bko4j1XmH2dwOT2AVDR6HXzw
OeKLtk5bEeE5YDMy7uFd9gWVeasIhHbqP+VkgjW4fpqMyYg98y6+ar1pwe92Mrgz
RcHdpeQC2d1PBO/ZEae51TI4ZrdNkIlNR6Zt1oajSO7jpCqgyIHPxUHKvVj9Qi+F
6WTy7oOBmYqz8JQRyBhrjLjBWWdOOkGQUhaP3Q/z9GWhqsZZps2PWWI7PFvISLKY
xAMjYEoAl28IwTfKy1UcZe+O4CYz6uo3jWiavgX9WS8bl7oUZb+7xcOjSqA1Zuc0
CY/i/KcPYJl+6dgoB0cFvVQYH332oMGrkO76L3T780TOShuBlKYBm33xJfApE4Zd
Abwn6wF0hd49dq2Q+X/k90b8fYZpHn+La3t0BlXOdvl1uD1Yh9LMxy/O6l/uwJe/
dcwvOgiWaIrAxkHu51euGbtQZo7xB3j+TzpGcBMCt8sUmpOerldVCpzsFsET7uJw
kUUzXN/QOVgndyRq2K2Y7SiR6Wu/hKY7gJTHrP+WFtWkBpFipTC9QkzBROJpxp/2
XapgYErvVSo7ZZBUq67W88Ok/bV/L8feDYlxEPQplgKdfitYN8vIyDzaWkNqHjhK
FDA2mqLPzBCuFyQ8bKnxVE28TjRjpEMji94iBZPaDXGdQsbmfmA+9uNFgoei3UtH
n9lC+qJJFEn/C3mYfvEYgXpikHO5d4BrPhCVPQL05MMq8mYk6926BUdE/TAoET4u
iCF5+18zxiqb+N7LaCJAH6Ag2o6iopqadsG7k/sc3lZCRMEUYuQPTD2028v7Osjq
F72SsnPR4G6MTc3ZMALI3koE8ajBhzqpQhN3KFHMSHcPbThZ9D/miPDeOsT2taz6
A99H5hRKXKRTVhyujKtGX0Mr/Vhne0zgozIdyRlRE8dyMx3iYq1YLpMkzwLbgBaH
JfeIBUb25HAo+QVchXshtV6QMJfA0aFnbn/O9bGPNj9BQPR1lMd6kMnihktvVRuO
KN+nOtzIPkl7t03UPVq71BR5T/Ow+QqwArInH3DynDDDVNo3Ep6dIexhJTlu00So
hlfKnAnZZhhP3rHTy5HfzjxO+L/YPP9N8a6FGlgRJV9oNVYaTlzX8DtRPA1Et8YJ
9frOQNlBCzqp5oUXhNwfpVirspQrSCSlNRnmcxog9HpAM0+gStwQY5vsPI2lQPjA
VZnfAQdoBjf8biOSpUzzkbHXV8UucPIfs9KQZQl6wfgXflwW/edEF91YSCmVdvWu
daBB/bF5+FmdoSUlRnujBrRTNvdkJUyVQZhb7uWh0djR8RiUWDWWA8UFTQE8u5Mo
LUMAGKfhSY+q9r7Ohaiy2/b3af+esJKwD7g0TKHOHuDWFVOFduVXkXgknRNMpCnj
8/wn/eLTfNA0H2U/p7etWAdDLk9mCCUCTK0YmhrxxuF2K8cldm9l7O5TqV/hGAS9
cL3+gMddBzCnOIIZIcAlKLAx+pek3MTu8hf6Jw8ittICvn1QegES/G/merQCI9sV
ATLIU9l7X2x37PuCHKpzRPXRTotcmAWFc5g96tglwo3txVxh+9UdwWWcoWI9tZer
09rGa6vpAVVa0bGC9WzNqmiQKNHlnwqrl1McMiCHDEO4YOD3Mm8KC8Di6QSG+x+A
NARfnQCi/nJM71cuenwLiljq3fMx3mLQWud+D4+0DPBCuHCoaBUiFr6KR0XGjVzJ
IUD5cohhgdhOKmblpoqbzTYyWA53Wix3tk4hm36wbg0wEidVo7d8q6maAa2nHru7
rBfMirWEfdDa4To2DV8HzoEwqG0er1BaThr6rOBtIx52KpA9zXBHw+eCjMXZTuOj
Rt9PO1PupKoTGsQJkPd5fFgLoJWID2/ZCTIdy5NaGu+clysHz4FSZOeVTmA/Ckb9
sejUTozA8v0mrR4Kup/4Luy8try43O+iejV3n2tjCXv960pf+G4SMiQuiigVcWMI
CiU8Hd4ok1efI/xE0culnrtGYPUVPjx5urbHndpZhpD1ix0f+CDu9+muUfCvRjzI
sQ67yCYqOn42HDYYjLLXsvSU3oZ5Ts6YV5Cyx6t71k1f3BxukZZ8+JfvXzUKWczV
V6TRTnEyq7F7xcffpsVP7kSz8F2eYSTz0xk1h1y6G+g6pm5WT+VGNVriRAc4eD2N
h6+KnpnyzRVfrySTv5I4OAup6nkUfkc1cBzd41MXbrkqZVPHo6UUp8AHV/QL/2Bc
a0RDEqasdO+95bwd9zPETawvWKHPx2z+i821jUPGSPJeI3diOzWJ3ezsvEpFoUBi
nY0C3KmaLEMOWEW7ejcos21a+gEslhyUPbqWhzTDe4WrK9v02lRcz1T76u8dDPIq
WJCY+KR6s4KxXJunRVXIoWRwIkWG7M1K0TIUI/i/VKP+//Spx6N68QPCy/ucJEM0
BGMwyIQHTZGCNPzt920g3rp3H86zw4qMxAP5AAljHKtD2M8M213U8/nc8gr4AIsS
2+xqoBO04mktD/slhe2kH0wgf+CUZzMHvr9gWVDrVCoVjFAV0picwDen2LHSeZeZ
lrGnUhtRM7WwH0jwv9/L1zPgxVaN6AdaJBlpA3LOkROumRvc3roWtdVcfE+Xze40
u2JDyJO9bDyaJcmdiqAgGHX35fIwExb7vpJvcbsySXifT7X4d9y5HwSFj/lH1pTd
xy4oIQ7CeWcUgxxcivDUj5OI0BxwDHAt6NVYvSTbb9F+gDKvXoLTkmRXHzo2YpGh
tKjjxfqfM9WjhRDawiQYQH9qKd8WLcEOOIWH3Os2ZC+TSh9HXWkaW9YpFPoFTesU
48B+tTIyv3XAUGUSu7/yHd+o/tcwza2XgUN7huZlGpcywNICLJ4Q5LzPL/bE34JI
Y+beD8hmmQDu/q+YmLI88yA5HwxNGL0Hitcvsr2vnRVcx0UogAoTNqFG3lacVLVB
3UVrTrE7ClxVQJ63ILnD3bYoSxDcs3WrsIdPfv7utu7xcVgRPCbgp+6NmXEk49mV
o4qd41+zpUaizFeCh1wJVEoTCBmep21iH/rM5weWAy02lLrpdPnPAuaJky+vIXTj
dBUgkyY9K+VIPaySrS+y7b7jZnzOlk1WH4iV6t5B0fXc3kotTRjYUGaOSJrbbaJp
4YTMMDSbRx+caa9hUTklRvXkmkkPLdX8dvV6P77xFYc2sPad2QMLLfl3MxCJXyKQ
8Y4HKxQ+skyjn/wUqHZVt3K61NPBwcPsc6KI6H5K6z8QV65nuXHVOnZN6r1m1kpL
MUGrkmprdI5BH0VesGYHN/vgvd8YjkwyXXsFE6Zqap8M963UdPf8QAMCotBiTnSS
2MNji6Lk9pBJ4dPlrsaIpfoRndZqZHc994VgXGSnJXR+GqU5n2oRPK+Zclttpn+b
Ldp0ujX6A6qt9HhTPpVNoARY536uZVc4ZF0kZuvBlzIsGYxgzqqgQIBUSAquAZEh
zqbd8Eyc7jKbGLo4QREeqrntbi3tVnAMBz019K2ntXNzhjw+jLtJtQgGdSrXY4sK
IvdkloUAJjxakewSEqjYyVvn4MciQiYpzlFlJtOU8b5fGKkZZnwAZ5HMJVMSa9oZ
NgYr0U5wDecfcrdRUdrpW1r7neUv7OPbQ2/ev2ZfC2p3z+r9CPieCxqPtjBkf7kG
hpo7Kw/oMA6pMp3wEds/bNzSL3oBks984nyht33YtGUF5ufZDRhCe+aE8/QdhAG2
uAr4CFYdUvIP0WhUD0/h2iLPV7x0aLcVduKB/pTEzazLVbsgQN1byYeYt8jfdOVI
o4fxEQ0IU6RneZpxgHLE71psxqJb9MS4t4D5YFEeQ6tq6miG63ftKlUyjnJF3L+i
8NPw/i9suJY0Z4CQKdUddB9xBMKY3xlHHWW54VqrO0CfmfB8jS/A3jC1NwiN27T8
LNylNakaHXjBzxZ6iKXOkltpNNZhz7HG/CXxWFcjlAmCeL6aKUHmjpC9kuEtI0H2
lRRK1w9zWRApXKNJKLY4g8rOREmzJ5Qv+WJVl8Iq2kLby0L+qFzc7ilF9jMVloXp
mHl2JimciBdBZ4WmIsR3h3ejMJ4eUTjAHNcxbOHW/BmTkuHqsbN3Mitft4iE6Prb
mCGKlXJzT4Tc8m8iJLL3nBdevi/8sIEm8Iy3NJgK9K/Ux9RBt6DZ/sDvv9dbNfay
cAyerRvas9iHJOhgtgcCtOv8tCM2ayoNBz+/Jx20gBvi53CKDoIO09NnEeOIaK2P
l6gGKmvLVFiDAWZFCfiqeJq9go/9qpoSTCPZK8+T8qTw0OXMMzjgL33MVZsYDAZP
5JiZGiyTelOAkwOg6WaAFsm/kNxP4FAq3Ts2eKcXcXDn9GNOSTqXGygjOdkyVds9
niFCozUH9mNb9CRVeMApoSUt1DUN4mUjHJcAae6EkQh+VU3kuAWZbIqjEpmjyikP
xtVLaiup0MrPHXQW0VuTaHCb56OwZ5scSrBz0izarNNdRST5hYxLB1IoWhzhAKMv
njHGRcxn6hJMIqERx3giFhkG6HdlEf7SyQEnfod1YWVQNqtwzt/G9i/MiainD6VO
5M2CVxNHxI4PFjmlbEzq0a2m0upNVkaWzDe+nxTNCGcu6EDDQUHF/nV6Xmi5APz4
3p45t99xVyBKgVtCBy8zuRL6BEfwnb+hh1T5O/IVAs6DeU99xFjw770qioLaJfGa
FifSQuDedVID4hnI5qL2CskPIpMjhQ2loNy74ICTzR+ktJDQhkrGTjmZUenBHlj0
NetEj+7DNcq2+lCw75LCCv7Oud8gScLqAG9tLZgfP2YjUnx0GJzP7pa5TFAroy9b
lJ5OVnCw682C91M+U4rWXVX31Vp8Pj7vaOHiJ0hBh6l/U17SPLh/yrEotHjw5x2H
LRqBooR7UTRKwvrtCv5xD4wu2zJhSVHPUmzl5L9dVKfxbmaTMVHpqlhmdmKiTgKz
mvWc7DhHeo3V437fGMFle5UVhkXGpHZ9Z9tSuT3FMp6rx+Wa8QHT83hkl4iJbtCm
E52mZ/Vs9QyE8ynqdhypU0GhGABXbFiumayuDSt5730r3Z6n6aHEqhhoucOPzVMR
OT2xaIAD/RPRPliwafU5pqI9CV5DirlmGCr3CV0lEQqM1de2c7SY99TNmm7xXUI2
dMtEThhCrcjoLQpyYrkiIsJb5KDhQjZp+Y9IWFz6HMosyY20ZSEXxPBCadb+pFmC
KFNZLfeiI2Y5MMHu2fcDi+MYf6IvkLIMq7rGa9hSRcOozBOy9c8e4GuXBL4adBlm
ia6lb/wW37x8eFJxkdaNkHWPdftnxB5K7OCIiBWQkrL7Dx4wLrm2Kf1VEoYXG3f+
i8ZBolM0RhzuWbYeRNnqiTHv1A0mXjz6pnppeANWKfhk87Vod5KgCIXXS4aQWSW+
Is/lonXkuLChgeyLWO0vnf/sRWr5ua/fqz+XE4+aWf2kQUM23U002CfsmBE3FVzx
+LmSgjoGYg2bmixsGl2ar9XR9VShRLL1XDgPiK0/XeKHTlFLjR+ONMMpqXrtOI9d
WeJ6Rb8BA5Ze9FLzKnn7MszG5fqA1CR7mpFG9XGVtph8KW8Uhvw7SgPtx7dcNWzx
oVZ30KHnAbdNMPDJSlE7vsJYyEqrPIjxSXqRdDAyg52l+WGRCXOMXwOlKMq3kckm
4t/hsxcGvxYW1AuL9Yhp8uyK76/6+hua7WlDuMUB5BaJZpS8vJRZcREkUYUtMzhB
W9kEKmhAuaMbwdSb76BcMoU4vq7KihJTxr0iAw6Rk96eeOF8JIRKunZEWfJwoRhY
d/JWoURQc52dky0EOvNwJ8h6tU1TFb+PDv8BH/IXLI8bfc4mtObvsr6DlVJrRr6o
FcKBeQPaRaBbqz3W2EtImJHxA7uFeK6OJjKFnmzK/pFCsJvv0VyKZJplYPULljca
HVh03un+SwvU5yfd94/IxdxFu2fww77dxbT7o0DwBob4dU7cRdpvzRPgLgay3pbI
Ljj7FjEm4JEytd9IbKh9ghz0FQxWJWE2bKIXOuRrsyuCMkVod39X6e43RdA8ksZ8
a2EeXwnV20+u+QY/nuV5MJjlpt0llz9+cQafGaz/sg1pJgppzT5yEKP0mZ4G+xn1
ovX9uAEkJ0wE+A+GIHSjOKGnd47uqzLZSMZbTOc+VXuD2ri00rusZHCbCFU+2s6Y
NNV/c92bKYrYFDmd9V2urC9LMy/HJ4aQxwRQrIAtl+396V9u0HDLuJVE6XJo8gRJ
D9fhB0MTkUq3PJ7w6qIvFxHhOxCuRpI5hH40hczb6gLU7G/1bJB2yVdpbmt+0GgZ
O5UN48GDH/U6/4y5BCtryc0quOOmpU3yH3yQS9bAa9EUO3qB1EZpbpyuER43giz8
QWhMofM1VP5N5Q6UBS2QJ6lDn2OfcpjLcHRn+lYMD7VC9fP6LF90sXIU2Lk8TVx9
QrA6rpf9zjSVg85pgqbKS4eiVYdAnMAwj2dvjmvXLUF1RE1/Ml51ENAXXn/prFFy
WoavmzkgLWql9mchLktZlLtUtHcYXKqlMzQ8S653rgrULaezhgvvq8LA14lPlZ7/
5Fsf23modZ99ztgOcoNh7PNW5PYZWq0mn/3TtqQWc46hpxw5DEmORcKuSujDV0Ix
TS6dQiLiBFpr+O4QN9jOh5ltAnvaoaEz7NOY+AB6W6EznqQrJruSiLKylPAQAPTY
3fW6Ylybuwj0R94eG872yH6DQ2JZEs+IbSxKlngIk/y3kIPTU0bG3g2EfnvXtgCN
EMp+s+a7EhtuONUTvF/qnobr1GbjG5dAM+BALqga8fdIVdKJ7Ph/UAyg0g0QIGoC
Xhcspo4inSei+iNWDM2BW4+w63qXggAq0av2R/jo/2dUBR8ipK3hN8Xm5FZ/Bm4w
ABIlVtbY7uEFIQA+c75PAA/6ooOPVRvHKWEFPk81LQPsQcgeSqDdrnDq9w7oVAIf
FNdlMIMeguU4CcmHfxLbmzivDEntiuVblO8gRXVldlxsMylTCoDmtdLT1fKT52F+
3RsHX39X0YfZuhjfYUyuS1aoKYGWgSWY6G4CvLBWBj5J3v9i7DEKJdyvLHts0oUh
wwvCdb+IYvqCyotNC9Umpy/awkVmWAwcWnYGRUb15Uo1o7S4wLly6ErujTfKqNl9
xhLJYibGhuGhFCcs8hk+r8wbXI8NlwTuAi4WwdAKifZykg96snO4E0JK+KjigBXq
rFjwT5gD3D9TefC4L7LF3aOQ2P1B0oevH/iG4ji/mQskMk94+iPblIBJrNdu3gZn
hlYLhSthj4yWhpKzMlGMdni5wK+ft0PUXypzKwfVHZzNqdwzgYpJXLN2nUuyjg+1
xoKwWszfS+DCdDG0RzoDbVpU4wXn3HFOe8mDvDICMXQT6KGMEd213XBe5yeKZAoB
BD4UYE3+Btd9Au7eYaRqd4sysleME+iOig8wjPFHeWwxvH7SrVbc21b69G1Z/UaE
1wkcEkFflE8tsFCgMgr80dwRBPBWvYZNc6r/6wLOpvVNyZtS+qJdSpo8QWcuJmGN
Sid3CATgXMZRnMAFDhZ1m47+GIIhKkmgIy7VFxNvjXfH/mxju3HmnGEstJtCQ6+q
/s3fFqMTQ173rpzkL0XHnBKthQH7P3nuDorzxy/ujBhbrrgnwxAhI5O7kbgc3tkm
njwhbGLwtrmFwJgJxM9qNwLJ8wsgGrLD1OTu0S+78DZv9n9wKwhWzHd0bMKcE2SF
VMGizSP5lhkvDnv1a+Re6xPTbtkgfn2UNNXgfMF6KaV9wx5/7w7/SygwXvr5g3ez
a+xhZODgLBkjf5l/EuFohr7dId72banhe/cdE+bb+vEbATRreCCz84Cf5URHTaay
5wgsoM3o1U2ZZnyIJi0i4OaQfKTHUlrxrC/A/c5buuHGBC17UiXDUnNsJEoXpAw3
lGPHifi+O4ewU0Y+g4ut3zRaV+tNL7ry8HU9ntiv4ExBL34FAVepMcvp+VaUTrF/
7WnxLlpo9UNuiw40tg5PYcGxhPBBnxIq2Lrm7csZ/HB5JyNm7gQx/s58Cs2tDjy3
g0ys9hmhALtlYQd3zuuwbBI3rdXpYxduvAcEifxpKfDwqWW2MFn2SV5VCqhZzwfH
+QaqyPqv/tEVqWPeF2Nhbq4uvka1Dagv507nnHo2ioG0QV9OUqdotlhyYxBIZjP3
OAzMqzfovy2vKfeWjUwHzr6rBtpeNwSJGsf2FXAAi4zwvbqbrzpHoFir7eNMaO9O
Rpb6q0tPkGZs+etMQNV0crGF4kRh0Qe/D70Wpf1bWW5MEFfManazJLfp+c70jSaQ
QTxMDQCvfplPopymNdtVFuJdjIYleJJlWncL0GbysFSJohXuVlnd4OdCtLoH5Hsv
4a/IQJrhgvMBW4ef1C8I/uu9Eg9G0DOhFgy5FSEGeOMbJTK7azm/f2FKu/uFx6/E
9dH2uWxC+NIHQj5BLsiENcmPbPxHIfYSn+hCXWr3GgZ9GWxN5niZ9huoPtgIVeb5
IKNKbJ+wNh/5hdFd/P5nevZByauwXx6uw/ctKCYRPYHG9pr2chaK8Ql37OwBPX8y
BuCHQHIHKXbSL9waaBL2CE7+cLyFE4JlwygsoaGplvkSL1FdF9bTa9WVLP6mgmDL
+ZJ4HzrSxiOawHcbA2yPVxuFGonhT8ctjgGfm9KicuyE9GOurG62DgRQPoPlt6yz
97er5+LmH+a9KBxdK0EgnVbb2uxx7603r4kDjBK/2OeuU2HJcGGAzqM9ZSzBGO0w
fMQyY7aYakOVqUhJ9FvhhVO8L95QocGi5fhPZsU46PDiMY/tu+CVoE6ILDf4jOJW
7Xncv2Qdeb65K6dBxdj+QUYsFMqcfI4ondxIsu84hdDwdCmueqH06ybSlgmWrDou
Hh2qcWGx5ka1UCcisckT6VRvszJHWEZIP3PEihinvyz53GLlpGmMsM94S53BGwaE
3tkuQuDfd9GQ2nUDJZKQRcwK8yb1hvulGqWfMskiUVTNztIsH8z1brXlZ7gwWW+V
+XuFy7xUp69JzY5gCeMgtXPswCU7apPAUQbb46FjlJIoCBGEq++LSTBngcfwevJq
XQKtSPrulfPtOVckbQ8TfPE7z+vrDEZ4nX+qFOrbdij7askw8deJe/xr1rS15bko
mBjMWTJurQklXaGMRdwm5pGLM9T6ko/z9Fp5X9qSlE3duVCKzsqJ2wBUtbWNerhu
Kv3hidcXN9Pww2nsdSrOxYpNkJHx3SpIX/m3ak3YQPEGv4ymTXnPWlvY8eQVXqW5
LRz4oYaOpkqBk60MF1+pWukNLQaFINfYTw/pcArQCSfjzQSk02LKfWGNuLbChvqh
Uf9GwKQySA4bIgAbwa6UwC2N9e7xFyXI0yIlXJGRshtO3nidTm7FHaJDdlRrGJZ9
M01cE0fljFcQaCtrlcFva7P3RAThh7h8SW2Cc9I8j7ROhk/lzWxMal/f84erpRy1
HH1dmF2pwMQLyLWMZvR7tw38KZA84LApbROtY9b2Ok/W+hV68zvkIOtnLYQrBej6
O5hXsByUiiw7hxdqKLaKEHJDxg3uoJlEd3utUxVkjBTeYYjSniPCqeMhq1YXufcB
Igk+jKC4RH9GSadVe2gwB+KOwijN/1y6kgFIqakaRLxAihvYfDfsx41dArhrhne4
99hrM7U0u072D8sBLMaCDC/aWiMHQR++4K8tgeSc0lJFTCAUpli565Qj7uXVLSQk
AdDQtQ9UGoMBrIosjuUa8/8D1+lxX1ktD/eTEEZ1mS8YbjcPOF1QklfSBcHuW3Gp
HMsB1eW29W9Pw4TQuzc9jbXF3MtZTdvmee+psxIM0ZfgNv7inl9b6nPKu24qZhE2
uGKm1t9i2A6mhL0U3FiByNa9UZVvoubY2cZdf5AE1gIqCKH3hhUWJfiFZO0pYEh8
zW4F+LgmyxeTsjP4xeTiSpr79ju9evsKAtEwrcx0ISaArS4KNIstaVCp/DCtStlV
+RxzY1xNCvT4KmAy78a8iD+ofHcFX20ffEr6oI1xcWabkflDbz67XmNXK/UTiKD2
+OhRMxrVZARJoiZsUlvGDCrAVKYuhkgSpI5zrj2wfHUTeaZ5NWCbVs5GdNy+/OGn
MXiScefJnYC4WhTO2diZnX3sZk1x3CH+goPA4MDyU8UtkI5Pnp+x35GrrMr4xf0i
Tb325k1UI5Il0+8dNitEQQjtTF6NhTV33bX+bMjD9V1vtQRQFkgicaLxrZW13hcc
UdwgOyEf/BZPzvEjwCoI04i452sycEJ3MEv2bJaFp3msFrAxOqar0q6Zaa0oUVzt
1CzxYaDtzprBkrDlYBc2o6UNeCuKxpjWDbIF3bxBalfHthqaKqDjMlCiD/bfyQbi
AnPkxgRzLwssHJTy/Z3eB1f1wsWF4wTDAd2kyD6DdHR7qbgVuU0mDxmjcPCy8+aK
8HNfpnY4RZus4uyG4w8vpf6nrcWR/vAh7Iwb9h8K/pCFYtS08YQxv6YZIa6NOeDg
I5xnzncEDA0Vibrtbct1PPLRfYIvLhaN9SZ35FIr0OseAORqW8nDmGEuR3jUMvSO
BGzl9MhIpaKuzXquTtld7/cAX3x8ikUaYqwxxRfMybmWivc/bfMjdzOdsNA/1MTn
9UyUBAVxeElK8pVeM3OxKuiL9ENrKuXGUFJFNBdrP3vR7adQUc9uXAGipzMd/t2u
7JFdzCF6sxB1h29+MrjIf+/pSXWYiPch2dm9F6UAKLA8O2cDd+KYuZpDdlwdZvbJ
U5EsxQg5wHAaZ/kVVxAhcmaKBtQctC+rG8RoI6hviV9zXlkaWBnS7F/UtZrtki3j
l+BlouA90C3CSvBd170leAHa2XAGe+BxMQxxKzo+1etfES14sU5cgodUXhTBgXR/
7AqeF4GAR6DIU6cxpYHmBy4mHZtMhV+Iuw5qQc3dt5r9ynnJQAlL6ATucovHNIIy
paMidKMD02H32HwO/qCyjtVjCDoW6HTNUrHdNZRZMl/6FGXzgeI7K94DqWrN3e0M
I8Xsy366rfcStkOSyOePK8MomshrKKOijb7qC+e9F/sX00f7Djz5ZkalcAzfrkg2
j43eg3KFPJMAAo91zTxlibdJQq6XEZpCUCOJtGiib52Jfp8W5IZiyG7+tVYLSQ3/
ARyUQA0Zr3u/70NSX+qb6aW1x8SH1Jwcb0pzmbT1vNAsngskmulIhY2FPhXCbptM
oi/RZ0QQzr5xLZc271GcaPIzLmCJ9KGjL9KkstTQrLHoup/0yosfII7l8jt1esit
npBfGBHnA15TBpVUpdl932SrlYu73r0FMPfGt/cr+lRLhRxYuYrcfkST1s/PWQsz
U4u4WCqazjq9VO0k0wLy11TN8Z7TKEUh+5sOwnkiPTxzvVRRmGDzKWc9mLOrgOig
2g3H2vY1keN77mnlrdjBKV2TWr4f0waxhykt8RYZzl5P/mFOeyVGSBoP3B/3mZ8h
3fn4gQvozRnLnpHQ39Fmuu9Xn3Mku6hisyIh3IIOb1e3YdxyZxF0Qd09Jf9jeFdG
Fesdi/zGVWKlWpjBY2t3cEie93vRXDXouoKm4fzbcKqAR/dAyaPVAEDHOZ6N/65k
2PZnT2+WODXPO0NE0nx/6J95VPwvvAU2CkRGysfRt0bLozAowZYGLMWUTpifTyQr
KC0cIta7nVlOBdBfHTIuJ20UDtDWgfzsOoeLsy+kpzbo75msWYhbwB+4PUof0ATN
dRNVs8UEc3ZqTEzFLe6MqORbduesJWBJ9zct3JuIp5P75MsWmzz07hkwc4AcbxFi
TKFrsa0pEJX6B92A/3wfvh3MI/U6DSHzgsuC2KD905/wIn6+4Jl40rsz5BtiAw40
yUoa84Y/vhX5uJeqmezCVr6fQ3O/5ajUQRq0Q7h+Y4gp6pamFcf0Bvx2pJpaAkTa
htfftzCs0HLezKLsa/O3jTC5ZbjVRh5pDKK+UKmtGqQL/0EmKdLVv5XAGrzZlIqL
fxg//rU3IcN0eFt8CE1zVdz8BAyxaBtx9XpHRsjQGY9rGM6w2fUeFpSAF0sb6+dM
+rDhU988wZ3U0KxPha+XOQhxo1qra3ZiIXEgqp4V7VkMRm+ykkFHtBCNsvK4twX2
5SUDAcuRrdrtbafzdjmpV4JmRQDfezb7TSzEcTMw28cF1O8/RWpC0spZ3cBjm8tD
gQY7eX2e0UQ3PnJT3X0efPdm1xfcC9l4OKn3Mk2WtXGtBwaT87j5cQeLF4F2y0c7
j4j2aI3dcfUq2CM4HjgIdC9M9gqW5/+1Xjsp5A5yHNCGjHmrMEM2F7Qn/1dGWc+N
74khrOIrNFJENOd6pwHDlUmKeUS6wA4XM9I4Qjamfy2W/34hYsqdj49fv99MV0aq
q9YL2Qyx7cdwakzGF1nsydz/kKj8we0iF0TPVgspE/uqAkzhT2PqCSnPtIiPOJKR
aXj/5eKZQ0vDFc/JGeYz2MtTFy/pmxDaN7OOEycxguVO3ml9+ClpOmqakYyv1X/v
pWTbosO+QvJ70kKX3E8aVihVwnN8vhkHjerYeByvu7fDwpwp6iTvRcDD1aOduMvL
M0kCBQIF5xh+r/BxDRj4+ZYUDPnqa5Gdbbf5Wd6OcbmFYYRFzFbz9ZtjQ+VB7Ace
uPuNs6gY+yaqHsRv4qbngMcjko/L+SIS1nt+9HM1yxpETS9YFPsZvsj87/7rqq5h
VyZwX78KmNHu+kcHVuPhYT6qcBiQLrPXkyv83d5h37QxvHd8Qe7yxnak+0P4cxFd
h5VlaOyWWJC92puvOY/kyvmzrMCyWl+l8aoPWjsK1fL227/eqKxPsTALcvvI0qdL
VKfDRXmSl4vvejdQ8OemVHCbnq05pp86NJv0Bu/EWi5QRnmWWqWYRTPGIWGGDeLY
7DrRDt7CuH1/4UMRqSfHr6TnGFdXXDIuoDkZU87UKeHgfGm1kJaLyefrHcQou8wz
JXnhTrLZHE2iQtgSIwd6Al7OsILp+Q5CpRSWUX9NY9dm18Xbh6u6EHKvJ+Z4ENcs
f+8p6ykv6Mt12XBfGWmSqcGFcLWgehnAFmvpctRNjEHSVywZYgOUiDa+XG4JtV6Q
84JVoCEPH7j1M4dQMsd70oXDchFmXSp78bKAlYfFPi2GeMLUJ+QcL9xSFTJ9WY2O
NPcJgrqluzuAX2BjDyz8E4yHUquCmQdJRn5ed5ehDrjVSzZVOslHqPphe4cToskE
pe69cSQxabcfUMIk61wkgUClC0H9JfhMQIRz2h123jjhPPI8fDC/1Kk4pi6BgUcp
aOJRE2zC7Ac13jA/tN3oWueqz08W+qvvWVX8ldln25INIhgkczGOd+xZAJC5P5R9
anJCbLxGcviu/yENmmQ3O22jEbAPh5/8DZ3GjUPX2pZ2EDNJ6dEsm6+B4Jv1x0yZ
GKg8ABSFWWuGvDgwH/y1uSLqMX5FiFaL5shtosbP9oYwyBWJzXuYtH/gtGIRbWp9
fXl1xjCHD0CDmyFx2bB0eOhcMHZ9/bY5XTzTKnykMUEVIGApxGqhXEb8z232LASJ
d0i65VCA74AwHhJY+VzN0b5itx7stMepgSCSc/8XM3k+o4x9QnquE9OThR49pMHv
JLss+dfIFmlsz1Rm8bF7r3SbQgt2KarGE3CzoTfIO0GGS4PlX/4LcwY9anBG265e
WypPJnd+lUK6fKm375jSf8HbtjW4NIwizoWDUcUy4c5lED1dCmf9WoROuu4lRIQ/
iSj6eAELESBXVuPpQS5CWkFMD9w1dMXiGBB0Yw24Hw4b7w3WQ4n/dROeVn4hcFT1
GdoI/2Lrs0FkoQsSEQ0UWPQwdWxSv/RzqiCYs6b78GWLGFyGfeV3jIop9GVtH8Fe
30AhOILKZvM0glym/9rtZ6C8QdTvmkNn7fTPV8h37qz3u21MjFJHKkHQhf3xOXA+
+Qcc+6O1t7JXoah5+9BqtSZUX9BqD6f/nAGIpsrWa6PXKevR8E6qIjM6pjUlzgIt
/hL5dorsz/XOn71vDDJBUlDYeTMT885XCtBNumXt8ZerjMjp9KOZVyHcO4Dkm5T+
C09BD6swNya9lQY1cF3j+s+lMKX7OajQh56ZWah7C0h6NqvVAo80kDFrzC4JC8lY
dIyWhsQbxLbw8KqMts6croFsOvTPaYTAKXiLNMjzifQIyhnTksLKGt5phm5NYoBd
azAg1uA9/ATn0mgXSBWI8q2HN2Cze3h8x2Cve6xNxF3I+eFiMDTVmjqRI0yX2Io+
rt0ks+Y4Vk92yMPzd6v2RSIfm67Zz1ET6ayp9hAxvtKGRBb5jO7+J8JXBkSp4+MH
GPIflihGlLhmJ/biIH1/oLuawdqhGqE7vt69BQ7OzKktzu8XuagPbFs7C0fBBx9E
LULnzZOK1RACsmtHyge0PHHlUfuJtYxvjR12kgPE8E4N3SYCHsnzdgGAquHjf6bn
Ucl7k1rsuSG5dGlq8B5TbFs41FtnfoXWxpyKKJ6Ngg/FMWp4arZjv+dV8y0WNqz0
o+Cm+bMjs0D8IrSwMyNKhkZCcXsa3Dq4kXrtqK+tzvm3KO01ASvINpo68P6yFcxz
coFt2HKuZbQEHGce8H9FHxs4KpXxMPKWAuQCkZOW3ux3Ls720tcy2nK77Q7azTwN
+ci3LBrgusU/GMdAIN2AsO09zI8QMDV7a+oLtqsJYJai00Pf/W3K4LVCkLMPTfek
Lwa5uelpKuF6CRoPluWieq/YXlHM73zUdQYJYu8HFrLWundwVn3ubr+TsXDHdkbR
hRjxx5/ceFlxFgwrDV51Fu+y1Cu0BGpyT5RkI7EnEtbASESSE9q6CSKcaB8Pj+SB
EnakUAGiBq70HlQH9kEgF2AoZ8QFCQRtqa+v9QvYln0CaAaa2TR3/B/ScaijTjBE
m6T858H6+tnBVpuHJbLPiqymobGLsw+f6M+gUlY1tZZ0867gDFR8ZbgdJ0sCmNOk
2pCnAmvmidkHZLzMDPqVYWwsO5SRss7sBEKMWPVt7EDgb29jPmQ8J/0RThoQPyAG
UgjR1tPaduQIZQMCUMBjwDW2XO92XR9OfG6jJaeFAPHZ2JYxKDTR8cFbwvpM2cDu
xeBQu6Ly7HR1JlF7tItKTmI4IpkRuBohh9IRAsmE3cZHCyMRKzo+qSEwIug0aEcD
mhocIGAy0y5s+hv1j+F6pHYBBLP2rXQJ4ZHh4f1anG7TkDQSkzbKhLmpvd9NRRzt
dcUojekkSesypsZVLaQ8jgGt5OsyOgk6CJ4fgSUVGw23EdLb1cHqEhokm3aXWemw
s6Vrkiuz4HtBTQOSjZsKm2HlqEcFWayk6aXbrxuxFLOdz4xpmfKIiJQmzAU4LRSf
IjbIZuqg2kcVGLJWjQ40SvPa2KjKNwTUi8L7OMU4PZkgv5bHeNrlBZQ6yXuz78Ii
3NlyRzoqNMbGOdNn3ppeTmFevNd9N+znKeabYkA6IG3M44kDmdGAMd/zkXuEllNC
VMCBch1h8JnkkT9jPH02xW/flG3631z6Xt7jl2j5tQPUhItVySqKykR8MNSLUHPa
OBwNptbWEHvLOeYNkAvDxHTH03U04EagiuDXNiuL1nDq5WsYn5WGVQkpHqna4EHK
74Fe8FXyUVIzFHI+FeLgasnqrCVm6Kbpm4Nv3HibvCcwCSKsXfqMzl2j3YMrr1cz
DpJkJVFYpaUEoPEXLWkF4y0msjtAar0TVXXpb23TMegBrNktPFo9GfH934b3oK1J
UjuI3ofjPftvu4cHMoOY9LcXArbZnchjY2NBO07rD+PSwOGMwJHDSDZVHNntgy2/
6HFXNetjSjkOihUU8OpU6rqwKWn2j+elVkJLEvNCj+qRZiDMPh2VpJxXYQKM8SIJ
AhOYK6yTp4m6m8OtBMR5T7w9s3PRzXp4QLwYJR7HvpQv9bbgFAV0kOLa1IOxYyLS
XeWcI/QSvimF5qMB/XG6UKEnIPVZaEkuCARin1M34ZLbzjw4dv1qZ7T0JfKOdi2v
dNIUNrxLGZ+RymQ67cqPWsKHfRRmyN4qClM4WuquC1fpR5OH5uv7KYoLYZbjb9Th
Kg1ENq7X20uEHbHS72PxZJXcTGgWF9T4lsup7mSpRG4UtA9SAC2scBhv8MG5KG5f
oYO5DPPsrcWB0oxQIYTS+RuVAGLb0hWH4eyvXQMksUescFMuo0DLoeHsHiiJp+ee
f8Bl47DQt8eTZlzityLO6QR/MP6hUmn4uzP0ND5pP6hCftYHoJ+UDZTd7i73A7hK
aSFh7qkTT1dFQOWk5s4KwMgUD3kPp5ZrDfOIA7zmtgzokfHCmfAP3thG7ySOefdy
1i9B0ylcpwzExjc3Zp0UabrX/32L6j2LQVrz5Ar/jz4lf+DT8gq85EaKKOF8rHox
VshWDcHKtADHPn/8APsFykKUiB8MiU2aA5oOfaVADYMBH5mnz+/SXxOMZciqjBu+
k8FBAgf1OWNCNtTr/WJPqY/25Y0g5qahayVsm4M013HZUkD+dUyd0mFXZ4dVxDKv
THYzv7eCF39CYW/KEMr2KO/7vhxQMWe/pRDSTMD57976EdJ/6cpicL4N6oDVM+22
tKbp/vGgn7n1jj2dLWsPACv9l2vuthIj65SytrK0WZ9TF6N69gGmzRvldpB0o3q7
hh5T3Eo60JIUFHlVSnOMFhJH5Y+Bn1/oExV5HfgJuXRG1FvQ4OeTPHggoyePuBu8
ySFOiAkubMOhGa5J4pYz4nIvETiMLkcYxqTXD34ueeZqSHOmIS6BYqyeZ5WbFhDG
EAWnFstKBQwa1RoQpxyyvQ24G/AMZcoyg1Bwfkgk1KXXNbaEm5shqWltgVdseE3J
WQA447H7Y9Zsr7tIjoDjeTSyK49yUKW4xLjXFnq7wAb5HBrI/o5g92vyG4TyY0cz
7epmaCfAqkFHGS/X6KRs25Ml2vA7WKQscPF4toH7c6HMJ7sCXm7WWP0QcE/Epp6x
l/LmzH8+3L9FY59nOkQlLoY8StD3Qrba/D5LmFZ62utaIzmks34+l4Ibe+j57K/U
8ZfX54FYePZLUdso6bx2crCd/Y1P1RKdxia9PVpUiagFJtsiGmu6N6Giax412j0V
8+ac0/i2O/hPH64qvyKmWpEflL5h1TDBAjAmmI9AN5wwrfOEamGiV4FjIgCXpibV
oOHj4BQLoz4bEuvpVLAZqH0Iuh65MkSk0loPz36VH2eTA22ChzweURZwJHYj//Lh
w6lwh1aYf2hK8/B1HziKzDud/Mr5zvFYVqMygkhNVqEk7eU6wdF6YcgZZ+uiSzua
5fCAlKQn0Ny9ALVscaoNkJJRd3Ou9Aax62b0MNu01ZaqMOsqVS9JRyzKA0aXCH5y
CRIfjhow6rWHmWr6AFaO8JzrQwnba2op3y2FFCXDx547aY81lMXEoDzXGwjAE49F
TW2dFgOWvQVrK85RSpyUlNVdg0v3c0PiKdEAQ3O31PTaJiOW8IxFXK7S6jqG8m7Z
zlLPNR+ZnrJjlX0XVv13OIYgGsViQSDTSmh/e3uWoappgoMEdQeBRONp3RwETTtJ
q3tz0g73NaAS1mWrNV56gkOEv1QkGIeeDXqHvfmzf01TKJaGcAYlRdt4Z9ukeRBm
qZwmrFCVQqsnaEMklMDCy3EE9ribvtTJilwg+3OZ/tfvX+3LRKkkf7NuJzMrfghW
jSGTUYLxo7IFkOB+0mnO5X5+ygbBu29w2OZocDIN4HmR+2M1aEURni7FgR9MrMVf
QBbLLjqH7TjqZAJeGGCXs+WWAoI7Q88RMD9X2oNVsUYqtdU6ojBpnYu+2CX79ey7
RRdACtn5s+V3581VpJ35gSmDbSpsr4mYg5KCEDe2hGU=
`protect end_protected