`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
Uy4DmKguuKHGYwV9sMd7gnMzpfgQ7qkLgS47cm4aWk5h39OtoYEpx/egHEQGtHUq
kZyGSqogHmXjazMq86VMGlRvkvy+mROn/0yVQ1MkR0i3c2nfArvaX7bcDd8JNC+S
ypcIYVdseslGmPQjel6hM2CQkDyDh5fHmdU26Dpixo/+HaB7qlVIXD0Itdq9x3mm
RVjuwGu942H+kvfd2Bn3aLL08lR75vfz/knEVhfsD5yBC+iS5U1gSJCWtViL+ThG
mHkGt9rsnuvSf+PY8NIWKOqqAMcM27HUA0uwEcBS43kqVFcNCthvWBw3olu1qcO3
RenFjVKMRRxVng7O+6X6nZAgenTNSdUgNmzPdYoHBAGWzAM46Xld4k4sodN+veYI
BHDoABH8bjbW6os1zH5wTCChsuAFI9r5hJgJSFKa0H8MxoMIz1gEoW5x7FQTX8A1
Z9qOIaSEhH1DKNuVFc2AfMJQ4qzeaaNeLIwQR2GtBkteZUPCui9VB7cKN75pYC2i
ViZXFBm0866uYCSY02b0hdvNIg7ak6sPWxBqkO6c+qUT1ZrZMTfvWbPN4hgmxbNi
Fx1Md2yhgJBgO8ZhhbQtOcQl8lbi9MndwkNlouRm263L22YGCzOPLA/iWFh7ElMM
gaQQR35Wgmum9AVL6L/HZpVLV00Xc0syuuxlyV3BDF5wTjtYsZLzFJ8Y1TSYJCCH
ta3aUNttq3bdX0qiS+zGkvJIRwoYV9djr63PrkCul8VKXJGbj9VEG5OfhYiRfm1E
0NnMyphR6O+3FDx6alrt/ld+YJem5WCeycoTey+umJIkS+7YwgZ2UzdfAvuHRVlN
3l2P6724Yc3ATF16nJl7iyzOQtjfwrtRddB3sRRwtjInJprmkqbZDh+PfZtQELlC
PFZLLHXuysPeQ3jchzfx7e716GCr1EVwIkMLYGfgl9o5k9nMLy9wgBcdgYCRrGKa
oactMJwI9tKHSY8gU1jaz51jQnUUI1bFTdeddrZDdmjzKGJ0vWQpZknW5VGSh7eb
j6D2k0hlLDh+QgsFgU4PDxWI8Fb+wPvE5HWAkoHT3cr5H7uc7sqp+PLRsbr645sL
ptgwzCQw+ZZ9Q4wi8+pIpvvZbrSWpBWtMfzFHquNfsuaGPfBkquvgpMTBYzh5oBE
LAHKT9QqgMNoXCIgKfQgBIPI1CEFvlrTVvTHEXZYgJymL+pizEKgkGkO3QXMhiAO
FVB4+uiIPtV28LM71rx9qB1fc0ofIkwPLpIuH+vlDE3Zl6cncAMepbixzw39FWVr
NWZv9YO89f1TC//6su0LQ0oh7De822xbtGvV9BRJ38f/KwJmVN4G5sMWjTNzgsjN
0gHG5PAfQ+2BxO9og+nPwadLSrgUEAAnE6sQaSnINxTZhrhLpHmrRU5yGihix6/0
ph1r4t+vS9pFbV8u2/PlFhYGy2ZwxZHj1Dul5ir7758Mye/TnPSfKrmmWldhPXbR
dj+cudOV0khl9wPy4pjquD+atkqL2UYLIjVmooq+U74e2XQnT+VbgfImqByJ5E1P
FWkqs8JYkpgZgzSdY2hbEc3u1RoEm+b8dSDa1jOb+KXUHVizHB2Ywgt4OGnm/Ftx
bfO9rt5TSZcQeXYySouh1yMOFPz782H5bFJrxOVIVvnDaDYd2CbeNibHTLy0j7in
yFCe3KLCoO3lGgLbV+/MFxCZdVaiB6zBXy70Hay7CUyeFC0DblgMGNdns6zpruQI
CYdJm61KdY/7B/giThu+nSJbrrGwcEW5uO5gkV4WDludMb6NgAsaZQtoOLz/0RMx
oAz56EWuIcDOqyymUPRWKkN9hr3SHKansURViFDYVBj654AumgHmA9Eufvop8zgt
08O/aMZkMM0PndeCcZXhrj+0DDN9elJJKz2GeaU276BxAuOY8XZGAxOogpNr/cVa
kLFLeYAPqedoDwywEjoKHK+oSQ3Bplw+welrn3u8ENTTep8QsViXFECToP69x1bS
WogaCNl1QcT7HNVZ0X1NwDXsyTF9EcaNFIwEe2xvcly8JidekN+ByclpopyGAqcb
2jvA6HyWVDG9ZnQJWvvayAVudZAljchNmNhUHt6xgaFPeDmeVKKztye3pbir8Dz+
UtSffouloBbuq8K39vzAZEv6CMORA7SpYuhGddwPEVvabVJirQwn5o5WfxWT78RY
WuRAHv+4dCrmokFhQSwSAf8mVpTDtqzyIFX0FUT9NU7h4Q24wDfIIk5ARxdm9nj5
D67SFeB+oodaXJebp16+MklQX8hzeiTrcoRcR35UWAgY4iRe4CLz/v4WjlFrh9rl
Nptqto6tzhILikb694eY/mcDB5rehaB8L2vQLNdPBHYFv4fBSCCiylrYM1ON37Z6
aTxAqnvihjwGJ80yHF50WX11ZVCUDWOAXFxlxvB3zagBSjp9sNz+YEHhoGHTtKQV
DLMf5ZF13IOPR2ss+8dS0DbM07SOnk5m6Qv5vIYzAVo0zxZLK8Dws70evmh8t5ol
9KPNuP5OcqJOCjFvpXypDz2LKb/6ZcxUYdchwx/0rD9WiTGfQHEjskaq2DhtlNLS
9iB75TGGk1Tz5Tps5xNhGbct6nE+C0YLTv5lU0R6IuJMLDsxjOE6MO7HveJRyls7
11bzlG1clsg8RJwL25eZvd7LoUzktXJxL3r0nMDoWyNfl7eN3ry9bexJRH0Yj1P8
bJDW59JQ5S7UDXZg27MctHd59D9bLmj+3TJdA6jNetkgDDlGEInnI+dvDieF+hTi
Mpwwi9X2JIWVDFZ9E8NY9spfHuM4p44ELv8EmVqxCbeK9vCc0er/orZTYUdmdCV+
jfUei3KjRgd0xCfBrPG7j5esZy+2ZWOUYJ5fu8aQJkwrjpHsS16gdU1MxTXlOniT
tSomlwo+e4oh7flT/jrQxsQYIN2npHVyKbIp+V2xmaRk9Tpo+1ZCvQHt5wl8/e4g
WVPVTQnOswF7VJJbPqe5A9oRR7eXT1yYg/ab65sa7qk0brKsITv0HuKGLANfxxOZ
+gulnlLBoebFufZDHRvYDOdVSxWiPnrsZWacytArTwgKy0JCy5WPhIUAGSiLQYxu
izr0bg4K+gSalwYMRhuiRyhry/dLgfboWBy2k0GhGtDTeDmRDfYDrPB8SJUWED8V
i4ryxXlcXhTdkDPzUTvOfH9pceROD5EVYLRXYlWng90T9iGXCYMwLTd7DC/jTowA
yJZ/waCX0B6Bue8L8GlZm2dYeDkjssJqrBAslis+3ZWW3XvsTUffmVrwhYsIvoh5
BgoS95S7qBP2a7fEFeUY6L8d4/6xyC1PX+ppDqIbCjAiRfQWBw4Sukw8AI9/HbMH
wl8xU2koDBq5NgOYCIEFIRchZFtehTU89m4X3KY/nMN80ltNCUDuBu/cKnpKCZ+R
upznYAEJePf8kGOnD+eWDOG+5v7X4MKIkQZJ9/hJhJlJtuR8r2kGAY44GtLK6khI
LZ6kA0vXsGMOwPmN15ZIHw3fsBlQQer/ycvr5GY+1ivtFR3A3oh+ZHNYUtLEQiAL
pJxh6gBFRaqz+Q90yb+nubCgm+YUv0BPeDKHP+5QM3aQLAOnYF5FUtMYvsYJ2arZ
xGjaAFR+QMcvXsmuYJ2/XLLDYjV1fkZDL05BoF2taw2YERkxioO9FfzyXjrDW1HY
3r617FrT1wE4FyztnD17NZZ+s+5shTPFbg+X5choit2+PE4cyJCqwjY0sV+MaQQt
UPDUg1qP0i5gEd9NkK64kJfCRuUNrjo+Hn7gN4eZY+k3QN5x1Z5MNsFnYDPOOYk9
IWKcvLUNhlpE/eQS+eKpX9C2+OGxH338WAnQxQENMhTOLeUxvt6LgBFkHzGo5flL
dpZFLk321f7bQvwodfW9GrUqu9J9DCKsYEre8Kan0w0i2EfnRQjI7ugCkt2rroDh
WQ9kACAtbSNn2X7XZhqKqdaQQhCgc29ujUEG8aCMpv5OQB8Gu2di0eI4skFZxxAF
qKGMYUVCWPOZPevjLGF5+4APjuYoHJQ0zmLwk1t+kBKcF+nZb3PVybjtp+3STeBQ
CJlwCGrQSjR1oH/gKUrO5AykhabOEVPpEi0nYNBDcvyaNIlm+KDy3uoa5hzEormP
6FsJeWY3gf0URu/+7l0Nln4/yxZcowTZ3pN4/fWYbrg0eVX4bijVCRPff35YHEo0
KxP2oXKlSF0CtikuAh+gysuhGd8oeT/Xx47GvbXsA6fffyvmMwLqO9Rqrz8ss5Sc
Ybn5slX900EK+iatf5rxL6/2Z2H01EZEUuQ6LCOuUmSPsxphd4g2c/CIFXXOkHiK
MjKU5nu4K5WsBAkLW0fTEE0qyyUg4TsgKHyXAc4NnlfVBXi8E01Rhq7NI4V8lSJk
cIDKqXiLDlpXPP0cv97qOxQ9fLCKLh5TPZJVO38hb+lbETyJxour5ZzP2qkAg2qk
d1Lkjyrf5r4MOkvO5yFzV34SOoH+fDzfy1zOprCMoAQspGDyR596w6kKfncrx2Pn
Vb6Oi4ibbS+VCppcSOEY+AaXXJJczUhs4OTIxo572Nk27qSoE9ic6J8eycGuXaRA
5u0q0tCId7oeo3+J6Aw6GGbSoInkyhxgIrwC2lQAkTu/E+QWQX33pickPaSSP4Sx
N8Fq4LMF8lFsVw/rFvN7vlljr8a65DSIVWtucZSgMajMOphYNSKW9Rkcajc+Mnq/
MyiViV0VrlFnSlKqWKpud3pSdYemCg1a6WHF3+tGN8f8xL18MTdUwaR4nDmRxFq7
SnvErgHC8TH5ARgfFMV7+EdiPaPesRGoLDUGBPeHRjgWJqeVOrWmtDiDvshlHeMD
bKliG49K4vcFF+oeycn9gE8o3016mWsOuuixrRk8ILN6x4K7+sn57hL1RUlDVPjj
eG5C+l9XR5LVlq/q3UnB32maeWQlNRMTu0YVvAm7sW4F1tmi4MI7KQgZ6mPC7Vsn
sDfv9UC/phR7UtSqgjvDZKPBgLPKBv3Sbj2tcCG/LaVtaGNgF6tcjGIGLsynyOBF
C7NuQTIZ9dIUyV6Bf7GGWmfFslP+aDVsgwncIjolLXEGnwSTxU5lqBwdqc7wPRy0
jDJcXTzkU7arZ4zG9SNDKTNCpz6F5F9b5UQ+4qBZ66Bb2sTXjbWISMD9+1NIlcyR
xPDfCgwbTP2z7tdD3pNfDEpNwtoGwNWXoymwQ2lmwI/pacrrwDU7zKeEFHWQ0pKD
9ICVHFdlzmWwWWBlTkEw4Pa8KOfkxWW1tX45WA2ALFBypAQfJBpbIdy/RuFUsqn4
u+1iZFivmd0cWnTXfUrVFPSWiH31KnMo6jOz7KQkvd4YDh2W3lxr/o33bfaadTAx
0p6+fvCWSnWIdIvFV84hjUvzarbJFHEJZdCtjPvT9osZp0JsekTcauN4H0lWSq/s
jfdXi34SqjbhI8nrUUAADfDVcFGIBPsof+x9vw7pDDJN6j5Hbx7CByrJ7XRr8oxl
YzTR0knA6wjh9bkg9orp2kTXvFb3WOEeAQbz2osT/Yu++gYz1q8tjDjJBkxiK7qP
oYUCbQLNzVLm3oyu+MZcMWpwIyoVNF9NIitLo9GBzPoFwstZMU4+ZlGInf6p2K+M
V5jrP1KNOFqeA0D9jWR+H67yuhny56t22FBP1D7T9GTd+xcx1WFEhAaz33F8Gosp
ZNeGXndz46CzIPFa9qss9yhaVX2dPDjZUSMnbjYzafMHt2q+5qDDpdZpfyL+WvMw
OgzqdqTGRJnulzPHTO1nZoxKSqvdTz8+KAT0X1mI2ULJoJdKuQsf/NS8ne1rKadJ
L17wwwsEzox6fRI17qDxsQ0U4/KRgEGVhgC73joYDfs8E1opCt1PMYT/hvozn4OO
0pW0TptTAV8k2opyDFFbCEm1p1Dco98UOt0iLwLv83cloSXO9IeJR1Q9jWicMGjP
pQwHydW34whOg7d8MkulXPiLA++/4gMDweBE4Yf+c/+V8WK2TZpYzwmLcbECiPps
iLKLiS+4c5J5dxKo7Zr5mr+QDEulKOba03g1qJP3XVy0ZjKErI0BVYur2p/hPxu6
ED1UQKOK5YhUJKU1iKzewlpEYNyoMG/O2hR344LcFALVVvs/jQqqpYwF3smq+GT0
Vsd1fdsija3KOBdRSCy8ZyhrPc7YXCPu4lkYRAdlUF3O3PFIGd6M/DDS4EShbxZO
cm24juFoPhGg8ONMNJhFxowe/9RTecmpKMGarzCiTy60Exh6eVJDhB2C/5KLkeOh
12O3LmwWg5nhbuG3y20yu7znEALJzarDJPUOj/tYVX8x+GsHD7arQzdYkJucNXyV
l5xufYyHTVHpBxiU8eAonOAXE1T4H9lBJ1AlG0s5xaWS8470zKlLlS3SDPWdLlCm
7fmvgvPV21Hwzf/tlYWZzXxB3Q42x05ZnzCzdRqxWp+OlsTCHw76l1KIYuXWHskb
JDG4rpT48BctnPy5YSnBxiN0dezBrMbcw835p6o5K2vhW2xVqqNgjn2dnAUND4U+
jzf677RZEsmosFx5lV2qDDvMXWSsfeJG4fvuvdyIXmK9BDn0AhuE3zyeT89ljaCy
8F23aCRRC6BNCIlOUDSQHKSxl9s/QcqLtu6eep9+YWVTaSFh/D8VNR5GFmcbiRm/
szn6qnpvoYu/O4RIAKLPO3yC8bgSt1gCa1Mx4WybJ13n9J3EVCtrspP953HYTUUo
hpU+S3hYBViFChZZIyZMrosrfpwjMGm5vDbfmGX6UFiXiTaDuS+G10JdwRNbRDWN
BuuL01TWcpu0Lc0p8ZuYZiOVe92aa7DJ/TxQ4jULfIYqJ49fOZ2FRS6bP2xLVLLg
JpRs2U3AQRC0xdrn+XGxPoYW52H4RwenQTJzulY8b0+BkeWNmQch99IR7HSCtWo9
6DiR+d/WcZvsfqAnojF6YmfG7/5fOBt1SxR7CIXCQr8sXgKDL6JW1RlJuxki+64I
TGIYNPkMVxkOoUzY1ja+qprKU3KrV6bIL81cJBFILJ4i/BSQIL4sKmHg4+Ybll1c
3Aan3p82Je1mZqZVt6qjYXksrCMk//BiqTJHup29R48myU0nKVU/EU5c0wD74jGM
JzAC3EOaXWSH51tydsQAqsB7l43qX7G0Rjh5Q9equTtLRYYkkavzZ6+8ZmoWorR+
aZOaS2KtcLf/QOZ5dRoAzqDMs0CyTQh2P+PMT816UFDoSn6Binp9W4fSvx51oWvA
vgw0dJ6m0IQzE347klQIpHRjZtSdZIq8zbrS5gj23x+kYOVaOw7S75GMDQxYlXzQ
e8FOuZmxRSHHxtk4eWS+6hsan3J8EduQuH8xdWMl8MpZAKVWnvVLBSG4/076eQec
WToZ0WCcoyL2jMYD3e06B5IQBNFOex9XwQnaNr4zAEQYVfnHESehPgBlav1xokd4
7wHI1zIfpiLYtcx93eARLgP2u4NwdV9LE/zWyp1sV1yPo/SqQtCvLww2ocZllPDI
pMf5i9t2thAWxG4nkFP+PQMbAMuq/r42jvIEW0yaydvdPyiKFM/5VxOp1X8wzbsh
l8RdfON0sAjKgCamogMmtTchiu5OTRvrpsrIl0re9FLA6gqGCcZ1ya2rkcz0iha9
grOt7pDoQEjuEwizJIVL1MPjWrGY8jcmQ2wlNA/8+DtQ+nRwTchi/2mBzuBZ2QnK
cv38c5mdXuk3rQs+N0wsCPdGaHPamAqtSYFWa06B0xMj7jQxZN76GAtO3qz5prJu
2Au8Fg4jkRWuUs/ODybvYsw2UNwDnkmjMGKgdv7SRySvG1XzAJ/H/UB99vAkKtMu
dP+fjSa/zPpWbSlsJNbH2gqDx/Q9GKRzb9/+pSr0siL8ze7LCEvD81NzcGlMaJg6
uPD8YyILF4WTdeHv3wPb+yF9TVsNwpRoR8LstvsZo25y1G2zdMfGwRFNm9fzjfIP
46Cy60g7NrZsAB0wlsYcIh/TvvjPMjb7PnpxSXb9yYqXkFHr8qNucB+lwaFaGvqu
S2J7d0NDoeot/iPRoZDA5R3r+ge/OZC4rQAGvLANnuBEPE4AIyj4dcJiZdc7i/D8
0ISjkCnDyByKjohgytPKlwMeISNZZoh8OvVa7r66NnjMSZu2OLa6XJrDw8veXzUM
SCOoumzDgcZp1ILApZM9FpOZlfkDmtJ4XtmrEUibsTUy2yayBKyrL2XFNCRa9mCo
jIKiT6KUf11iyEO2YNQEis3bq/DGmR5URP6NWNkhpcX54X+BAb2jTgNHDsXygUpj
xpX8miTt7biOfWEQMogmzCH1Pk++tCvzGvtiS0BX7eOK/D2t90Emn8ViOKmJGyWi
FQd3tQyCVAfzzzX7IkYvPrjiEwdoFCt/9rlZNHLg/Inczu0u92B3IXnYKI5vYaLJ
aXi39iWw29ahw4cbAa9/hHig7HVP5NTWZWYxwfzDN8G6rtRdgwVHBDjEETjFQ4So
8uxSPPiaQfgKX0/mu/78ohhi9kq3OM/afzZia4kJnscK0OLxoyMYC72RsjA27HG4
FbAEzARPGj1A6SzR/LSMsv72YtsZPAOI5XufBPOm69lHTYUOnbIpKL+jV5CQLPp7
MPFkHomjHNCk3CdNbWcDfivHz0bRMjnGMvlisEm/f87c/Kd5meLoSfOL/3IRC3YM
ZGZzDgfjz+JlSGd53GIA2jZHYn9PUi9CTU65HU+N92CXoXyEHZqI8ui2g08WmeUi
JF0un5k2GVNwfPTKxelnnJ20HPrKTud+FvVBgRazTg2SSqdllFbqHGglVUrbJKNE
dO2+r8zuR8gEDURTKDpLYWKyrwqPCmSeVisKA4OHIAPz7LtRD5RAtuTiYZSkySaa
friB3cjQ3g//MAeLpqjrlgQo1CTTE4NoBhAAy4SC8CM+ouVM06u0vb6n7KFsj92y
2AbrpqpWWXzRB6x8MkcwPTyTDRPwubURzozm4yLzfoovM9MVnBUreK4yP42+7jIG
WnnkUdNxTbgHJKhWOMHxu0dEbwhOXwdN3np7JDkE5fX6ydUDvo0Y8gZTl/eUQGlY
vZUxQAq113lgfnw5NtQsuTS/9czInNfMP59IQDCKS2kegvH0L9yKsD0kd9aQJs7S
oK9ZBfMMo0p4GP3m50LSsdvoXa72R2SWCBOvlGs/J+y7EujCb9Me0ayA3GWzRlOY
b/+VUI/J8QjKe6bxCzlfXDIbqBSDW2+z3k0Ea0Bf6CQS1OdQUAZRXSZQayMxg7Mi
xArT9wINXBw5aKjoczDPll+sJp96ITYx4Q+S2l5m5uOYVdUm8iMhNnMVtU+E6Vxq
hXCnpojvukyw9LHrBPWxCoTKKgoA6vtnpY5zy6tCtNVW+2mYp5wyXwT3QxNLRM8C
w2vCL8KKv4ObpOKfNJ/h6TAh93G6XDeW+afsYZ6jLk0xa3sj7tfZ5dQy/GrB2oo7
Y/asFjpIol/xy/7pDZT0SznciBakNxHYgxnWJ/FSi2nU3LBsgeAL8JOUigcLIsk6
2E5HuXVa8MOmg9DXJUBYQk1FaS40I1s4duYgtxVyLpcohHI8N5cLc8/S+2LEpCir
OCgh30xXaAUjfMjaQkt6OfgjXj03hikAqcEWWIR7VlRh/in3IsLOcvHq+ClifAjl
kBB1GJXB8pWjgvWEL5crseUVzxanz1itFl8nmTrvgard4CmjFxou7FRVwKp5ZXp/
hUVcRAunsPLUSlHCuirH7yzYy4QiCDhvgD4zzTAG21Xhw6x56AFtjKUe0ZMC8sWk
tW0LRc12zpgS70Q2+tIG9hNNMQfxcTtMQ7Hb6ZCizDqG2K9ReGrgajJ0AhZJYUG4
bXURRhDn4B1deSEg5EI8vBxY7QitTPyKiDoUSTgCj2PLxpiCFOHSj2P2C4wFp8wp
+c40CV6OhZgQoSzHvlkbva8kGqmOrjqW61rolIWfNwZPaMUQgcZ0yXruXmTsnCkE
zvZTi7baRzHNERC9YaW/YlCl7LrkV0wxPal7+S9Co/cPZ+beQPokv11TOAnnwPRz
/ygu5hPJgF+HIzX7a1tQBXjNkhYVsvZCOlErKZAapcb+8HjbWls+j6EZ+5yfRaO1
geZ8l1mbg3Mlh1OJxeUzV2Gq9iyWaWenxmqh4c1Dw0GE1qzuJOkAH2tbXJKy2vHX
q701whqo/LydiO1O+QR9uqU+MpGDcqE4NyJSWO5CBd0FVLbEONlV3T9p8ohEl7hl
vYiucBXE8SnAl1KhYrdmy+Rv6OU+FFP/VVyQB7c7LNzSkxRq50zE+Jx8dusjF36+
UI1LvYFHpiTBV80WFQQc7zWuKL8UZA3SQB2EeSNMMfMUA1aRkb/UTlb/UFlFBCpi
jjlbkkIYYMyAPBiZOlq4Fs2NR2bued3WG9ygbYK1nEUfVoGDNi7wRAeOdvXKe6tF
Ohj/Fb2pydlmONKHV4nEnJ/IiAUwfOmuaZitEePMelKm+FVyobWkWGnEcxmfgA+m
y/8eYE2HYtq77VUOj0mpGx1z0y++Pt6FSnZOSCHQUw3Hq2/9aquNBbu0Uuc9e9MU
LTaVcB0TsHnGAa8BsL5GUmWSM9DzJj8QzWOi3LCGNqNcvxUZvCMYglZDOSwAJ1M7
iIt00gjev1zVXWhjmahCkQfUzslUaklmCy8iDJU5wtX6OOxDzG+G8zq0Ruo0segZ
JOV+uIssI5vQGBNECl8ru7TVMkPNEba6roawHR6BzMEyywBf2hm9wocQGbQabK+k
v7YbYPzZkgEyfDbkkChCl1SWK2RI7JmpiYgJjIXbesyvrdP46tlbG/VbVERCp8W0
3TDiGNRawQl8bHb189dbIgmT4SS73pkviiB8VO7P7jbweUNeYq4VIFh8ZyTd/rlW
GQ7bmBKPclfkm+fGDiyifgpov5Z4yI1ONMQDHgL7LoHL53Tgi7RUm3eELfE9wqU8
TMDJVz1PNLTgZVPPQ3VRiFNROkbU+x3QMCmxTX5z7GfHeqvEGTFOKB0THyiy7fVB
1YbvXwzIlWURkE64fm9F6NRoB258HR1WCXLtbVjq9UtspDoJB1j9eIvWZQUIJ2Bv
aLt+myYXIOTT3ycVcpji+dZkGaraQ4JrSfE85mDXxEJEyB/DbKtaEprf6YouyC3U
gQ8+0NWjEi8CCSwoZYrJc8rHYK2KxvdyC1WPd47BLn+JlbWBBTLLHfUsHFLMZpBE
MENWsQz8Wci4zkaHZHevdn+evdmhTj3NL4gHx2G/ve9mYJAfH0yQva+Pgvug+9UJ
dEfJznN9vSVXeYkv7tgCvBzvE839j/j2ubRxEb7Twf9Kseo5sM3T2IU6a9yXpzah
IgE5VhSKVr5m1vOyq+SoqKzEsfet4bQuSSV5X9KDHo0PgY8un3TzOOgjlm1JPK2/
y6Fyoey+jL/ktrVUFJfauBaftRLkQAN0tNR1dZPBYseapTkWpARcP/QCy3ekQqY8
YCf/LgfUZqkZ8y6l5+3Du52xlBJXoQKTrkpaJa+9WMZq/UB+PlMqaDYm80jRPhhB
OiyM/cXNf6m20BVn53IvG3GbJFfERu8uvD2KO4nq0SuzzYdjDMP/zmZgfgEYeFrq
jG7CJD9tNvA8gej5Jg/8wH0MMarnIJ6dSOwmK5S6nPz/y6C+ESkm9Hv5OK+AYyO2
k4BgW3AKZf9TpZwSBsgcrPrrCrPbkKqiXOIY4z/7WpSiOYyXUZGELiS5uAgDzTHX
cnnVSEt0PLAsWxx3Un0xXJzCSZVi33Knx5nUpk6wzD1PdArR2laYtYcj7JqP/ziX
RZRYorKgjDDFT1hWDM3X47TzUEksF6c9V6ko4IitYVaUJn4hzhuHSzrWzXVIDqgo
X6qVelv7DwpnB+Ke1suUQS5g3Ga02Yh+coOaHm4vQB3IfcqXiWplDLjXwJ+wJ4dk
kjUbbGmCTjesrs/pKNq/62ST9tGCqQFq4roouytEgP6ZWaUvGsQIuS3VMgJ63zJb
u/uAI942vgNMlQFwevJyY+SpNXbA649ZcXs5Iu0qhdFx51uAHeLAJXRmMDTGiBzF
22vMw0bHEIUSxsfMUy81dKVok7Y1k8VMkQYL/qgAOZwtkaTj/CnBqIaE8oSitICu
0T/iTL9GxJn8KspxTfBRw4kcfxPf8kv72rCj7koUvr8ekCnkDHAEIseaxCpgxWQA
9yah9vVKttuA5r2lnCeXk7WBTeu7rqDutkDRT5V1WFDMAry1gfK7mb7cvyOkcQ2N
h1GKeeRobK4eI2CcbgiO2Gemq8pZpOvsV5LtFN2PhHEBS44O37NAjRBIsFHxQuFd
lh2oUR+slmOWWfMI4/kXQL07g1Hx78uWKgEBkVmPYfg8dTORIpgqar8JXSzFARdI
FmTZrn8evzlIPc+IItAEV7CjfkO5ac2ooK7XToXC5CXg+k9r2yb9UG9bsNocnr9N
koH1DvaecZQLCkgNcGvhM73+ieoiVpqivDroX7AeXNEsTaceZswhk/UUgiMDff6u
HLN35m007bSZtwHjsxIftB0AzTeSoFSrhHQsZIRIH7QZdmhxYkPfUrAd1biROsYW
3j0uWLETaqXmZnCt6tjxISSBHQ7YYqq8XQQ6mkUo40M3NmRqLNfIgCuBb1GR6kYe
XSJD8J3vP0835RZyXiKn34QN2sV6oLXsiAWrWZwpcj4YyJtmksczANjFiiNcyW88
6J/OIhXCJWLKpBLKL8jnwFx2V3dy94otM9ozQ8oJexOzDo+RMjC3GD1WwWDPhz4R
BU6TPTRRXztg86zx03oLk7Eu+BMr+Qp9PDNTCwl6S/ole40H0IYHfJMzp+Xa7ZMr
qBIqKvwBDr7xv1O0HRtIzzeL/l5KAh+mjrSLR2qu0iOC8H7FEEAH9q3Na6LZsPrW
XKUGHS6gUAPJ4oEhxj+49Ul1mQENy4zxMa1EGY9ly/7Lp7m/3kMfbh72MMcec18m
GCM3B6AGHkdW+LumggaMi11i86lEsdBennyzQzpz8E+mXp+UEZTxlHryyyHH6PuH
amGIJTFpvp0ATsojDmdzzrdbcvapY3h7dfQHaUMKIiGuf/KdWPrvu2IVpWl7eQ6o
Q1laTt/dikv5cBqnmk4UQ+SXrXlgEw6TzOTnz32WRlYlpsZKUrCy/VB2HLaLwNMd
H1KHIFD4voFrGPt1YYiAODlVkLWE/XZioi7c4pswRJu6vJSRU7NP2Cj3/v9Zd+rJ
+HWlQBAXLsTqGLgwE1l5n/7mrSP9a9pAWk8WG+YCFKXSQHCApY4+tH/UasNOOxhw
HdLgATnUpyMAF6YqGyuYPbYSp0EXaQuHeJt8Dcvrl/nlxt23g0M6272pHQKB/IKQ
89CRMfRNcbayWmq3wAYDm9Ni+WkCacglVPa3n6LncEmioo1YI7zTkmWT3NMlj8gU
FWIGog623I11qsXd2jKRsmUCcnA6X+F9H9LqRLwh0akONSDKhjYZup1uU7O1Na2m
wqIgeYfoL2m7QI2ozhaqpnjYBvRIhkS5Ssz9+C/WhTxxB1JhWPHTPciR6l6GeCkb
t2kNnmo7LxsI4FkiuHapB9QNUGoxfBvbjR/JBySVluyz5UArLyM+7qGs2q1S9Eev
iUF/JQIjg3Ncb7uksWp6dKbsWoxsBTVVqZyNaiUGwi234XYLxVf7w1HAIH1/v+CY
qmLjtRBJZqI/MdYa506rNJkMJsq//XCQ87d/MCAGmCl8a2JWw6lLI2c3bftEDxMi
phLz5hj9uTFkl8sfRJo5Q6Q11ZNUx4ICzMmnnsyi5rI21McJklw6RLU7OGgEQ+SW
froqilZDwPPOvJ+nvDK3OSxeyYirKypygVaTkrsQv/FNEnFy4ENhmpBw0RFd46p3
022nlWEfCe2jPCb5IU8G+TnWTUZA/G6E+xTknQ/Qe7+18xUxoGPlePsj1rwv+gZz
8erhgAFvUjcBF1eWoUyISbl/u08wlk23t144ebYCiGkEP1eKMDYrR3/9M5rdMj4B
g4TMTl4ltFmsyy5GzoAhg3+0mT1ucbPTslyuBw1QOVwIDURD6sQVpuhwljJgtuVl
nivcc6bFOuq/yvCzO4MPydO0brCzxOjIULKwohSYngX1ftkox/SEnLVIA8gXuGWM
K1OcGalvoY3FrRjukbnof29CsfubrfJyqbmeJLoftgwkQ4qwvyCmiTL+KJ8X7svW
CSmMR8o17N79uwBjEymhliiU+Vwu7BzjKu7sWNz1AKUTKhGvpPYgXKT8lPuLvaJk
FRehtdAUgpRY78V3lehGtHgVHkMMimno5rM2fCf1DfIlXbPG4jBW6UEA+WRNl8cI
gOlI23/1f+CN2XNrT5qJVtY+KPJdIR5dUCY9W7Y3sFZMtn6z8bckOxZtGQXQGVu4
ETLZnN48jQoK1xg48jGf2A+ev2oMNcuxtJsW9wAFwXVJOm155pDgubPBOfaXLD5K
Zn8oA0vsJclCGSpAAwAbw95fC6wmI7+83AtwV9lD30Jn9Q7fX6W/fiSEseEWXbCd
7X5+vZTjxHZ9sWDpRdgvFo6fi0yrAupf63chqLpgxh4DUslG15PDyUIGfY6evdea
GvY4og7YZBvksVhQX9EqPUutWCYXm1Zm3zKXvbNMi1ilJJ4YhuIJwYlii6baDM6l
etrXRj2ltxmkNrt6UJNhMW1JgoEdz7+bf8OGvhRtmb7iXgy9Cj3COnh+QpiWqmHv
RsJi/JA3o+uUVONwPSA/3Or1NqlJWZgpGOpLrUkxZBMgsq0aEt/9cwI7aLlg8xbT
snxYi1N+buMLoQYJGBi8KYceiT68v0zPcEqUeh6Osn0pcX8GVIGCTzHRbb0exPQ2
uY1nlvAKvq4IKpcWx/8ohB/wsd4uae2kxM7wyJTQhb8soxduId6z7B/93F7+s9wZ
+4pD2WY3SGnNUt/T5IwJTUyuPQnbP71tjkNzp+FrOUmCgLQmTXv8JV4y2FgixuBC
JH5MEn9ctFt6FwjJUWMfWrx88zttV07LkLMRfb+Nxh9wfXzluTa0HkuBzNVTKsF5
p6Z5676YKSmp2qnZqb1VjRFUpoy6X+8wMnoIhC0ZED0AHUEG9Jbo2ZLz2GPkgiGU
uR0fR8gODbJGowUqnwiUMDpnVuMGhnozF4eCexFjSgOSQFdrnDC30MB6f+crbq2b
9eEgHnP5ma6P0hUETS8ghjGeQVXv529EABYBV+h18PWM9S5ihqX9d/bMEf7s6bt+
WrVdnU1wij9+pdKBzlVZWkj4uSY/pHDiKDsoa+cDn5T2SrAsQbVhYwf9Hpv4Rvt0
LBPoJHPuip/sjK6uSrfyy0uiekXwRhgWcz674cxZ8gy5Kr5gx/8p1wd1qGhVXXey
su9c5H895Qe8navmzP38tLpGxh44zIoCU86EjbhZG8+B0IoXBAfjSf2/MTlrZzS/
z234Xkwcin5jQk9mi2f0GJRnhHyFBkgXrg37DLVUTC+kGmdm6iutibNjocrUJBA9
uyBX57DE+v9g6K/71z36iYn+1oVNrz7YnyOg9TMDd8PNTYX5HdndpOeAhi9jZ0so
j5gFiWeVOpghw1nPgdDP+cv168pG6Os+QQiEOJBRv2adOvr5XNF+jeDfOHxC7Yv6
Rg35/NdXz9ySjDT4f3Y+P2pX1Ga65A6mL6bxODyDX7abLl5tXUo0+iOQM4D3v0KO
3xYstzumUGRgYIPj64OSHmr85r74tg1YHZkQet4pnUgbyDE6Ds3PzF8Ga5wtjNZX
weInminevZ61hq7ogJn9QUEOdyOjlqKEdhaiI+zMIwe1NPiWugWIshWo7inR97vl
iCuNF4N0e8n6asQnHAiJ0viK9HGmqwt4RqVd5S+i73lzEcvu8lRHnR32lIVYOo8P
XqRpGQjiqajErdvxclhoCZMkEP4Qek4vTNKVE0AcsR3naEh30GCBUSCVSmQKUDfH
8xvm7Iu418bqXLSlnsX+F0cWg/dX2HkSrunqcCAuWPTXLwDo6aQ8ok9CZkvu0m01
cS5/ZOmi1cernhIE5msGe8/MA0mE2B9jhKBew8CghxSZ/DuE7UXnzJXeC6V+m3Tk
X9WMgp8lSJHm4qR5bVqGv9UGmms5FlhjemCNvGEBWzPmNkzwpiapOTHnk+8EFkMq
bfCJ8Y7liJfulECJ2rbozLdWkhQDDBUoGqJzxyaJAAMdohgy+hnQj9PxVTCz8t5I
lqdxXR3Z8Z/r51efT7Q0mSeviOWScN4AOtKskzzm8IKDPQCRqwiWEts661OUlNp1
ZcI6bGU9wGcbNu9GADRkNFYMSqkXQTrMaGw+7ppoDp/KnobwRymQJP16e7xp4Rvz
JrYKEF3BbXg42ibTg8yy0cWeLKeGbXq7lUMezyEcZ3JcNAuVYwNiwJDyZlkJl+IL
bNZSwyOiHrlJH+eGUsFr6Gs67LoFym+Dac7i1Zi4VGhXe1ArySionpYEzWNLgnxc
DnZoY28fiY9zoSrCQ/PvGePW1+Rh+OKp21iGYCr/2bRA8bHjzG8XlOeov8+CkYhN
1eNB06hx4S1e5mV6hvOG5pVtIvuLECLB0nXoPwdnX/ngKqgnYhCBK/00q2GpBOC9
VP0l5gcjAp0+ekrBRp0nWCDN5iNoWlbZDOmbrI2j26CKRy0c2oGYB6VQfCSbP35i
D1RS5KGkVLOaUhMrJfYu6DYPC6gULtYopWcr6KJk6rkhGt8FDjT1y0cwa9y6QZn7
1JTEDpC8vTSh9dyxtXBoOkLN4q9trdhl5uElq0d8+dNy2D1HhgiSmFQYTqBPuQxF
bBSNOM4JboW9WTUfbGtBOdB5HUVmZ0eHxqjyyJApQSoI2ZZU8ofPxEQgV5V5GAfW
+OOZTZfvDk9bALLSIE0RjZfxkZfEcdghju4GiA/RW2sHAjLphGK0JBz8oS/JXgpe
pdFxRjPKXHQzoCHQ0BNPIGlA7zB53WHEr3zQY6TrqxlGYn6PU86a+s8MoV4fWjNC
Zf+zvU+Y9E+S0of9JAQvJvWelmIWZEEbhhk6ab2QaIlpsNq/hCdvax415W3BVWFo
rKsV5nr80tMVit5NyyljXvxA4Ocpf0GPsYQAMt1CKuqBLE9XWamYdw9h3RkFUm6j
Pgijk+x+TkLoJI6mdREJ/FBzWvs8Zm9TYQIfVcbDaPo5MxTGOBoBguWGePaZRLXc
GL+VSsk+luT0tolzBs+fN64cX4hZ9VPnVUPMxenjZ/lTR/raVtZxYMsW28opDcmr
SKCx9rpGhGBnnI4eTicwhDu9ohvTwTveyvcEe9PlPWnnOnLBrIF/q0l0cAZdYbY0
wSvwLbdxukukp7fDkZa+VPq7xsBx41Mel2Xc9o0RvAARybNyoq0p/Cl1LcMfiYPi
4pea8Co+NlC22g7+xiJJa9VS0t4pDnzqe8XenjBjy9zHenNaksza1Pqz4sXKd99U
1kYSz5FRGre7nBJfGLh674Ui/IStnZtJuUu22SWdej/r60QF+nTOOnuR5kdkTq+A
gs+XkeqP0CquwSHQuzwTPT8ezEtayTAr+Q+3AYz7YEhmi5AAEw6/Cx8kjDZ3jC/5
dcWQp3gyTLOHTSFQGNbTCV4ZuGwsNRDUqhTxN9/xeN/H+Ey/wzxTJkBIvqV77i5e
figBrXbAFNrbX10hBtrz6TLXw1sYe5qCezptrvi6ZK/7NPJG+qKtSNat512zHft7
3X/8ahshfyN/fl/141xVnu6NkmJiBl7kEfJ3EwpG7pcYF6FrizT2AaX50Eb7/A+m
mtk0RnvMVF9bRHhh57vkZVIGvKlbRTlXUjzr3xZo87+Kzzvd8gEN1hY9AnXc6Ltw
CYsl/pck2AjisoDZQkwxIccu8Cb7WAKokTy4v7210i03g3ffXKve/438AWlcS+vM
GxapfI2cL83lxJcIfn4y2boREOn1nog/73eo/V5x+N1tjAa7eLZ3SqJOam7Kv8mF
9vTZPv1+dvA47yfhqiYKBbyo+QJTa1amtD+RfwfOQHZ/o8P4ROKGY8T7Wt2u/R5K
CSHNmSLLVBo7EqJz1OoPbrnbHut1n1v6MACKIRiA0sM5Pmu9qRbb05nhOUgC9mRs
5nAdWDipb87nxCSL17UeFDNAWiZyDGz5jV3UIsmAjSZDV2XNU6ZePrz04v5Kw1rX
cJrcqVxSqxtrgUDGvL0D+Ke2pX3xu0GbftHsh7Tgsi2l9ovjsCjlWOCANEertOxr
EPmcfYwde9/td6rd9idCfF62jqhJyWnuUWd2L/v1+qst0cr/0sPXV/b2Z87V4ADJ
5SLj2lRZDlfMA7S6H1tySQfYovB/Ug3qohkdo99cTcVxgi0NjDEw+CZhP9ioTUn5
SLVaFpKDGdtzPMZsPNcYuu6R/yte0QzAiigoQTKcJMwW8yGd1BXVc3qOI1BU7cVA
wjB5ecr7AaCpz1pipFTHTYqrGVrRV4k0qeTKr577MRgvrGdwhpuCIk1lVXUCL4QN
82gB88rdvxdIlECiaAktfV9227gR/80svKPI5Xomjypaftnhedz8vV56fHvOL1zC
+Lu5h0BE2ww7F7fuWq3QBTansHR6CuvCEdSsy5/VHdYd53BHTOD0UuHa3UX23v/Y
vbZlk+Kl+ZmEqKH5r5U2RZ4a4Pl305lUEYUChHuIo3oxKV4nk4Zbi7w2m7m+hwVB
fMUGn44f5Wibbb0Zn+Eni42q0ah8YkLlb+QLKIERFYkmPGxtXyvmwe5h2/S48fJM
XEtGVn+qtvo7W1tLlPAwNXrGC2FY3NVn0WFdO2cNas6A3vJxn1EeCYtg3Dabr5bH
0gZamvaWgflDqT8FPjabC1v+oaJ8PoD53nBn5nL4WkwFMUpOdb6b06qWQ6DJZnQ5
NsViHWjrgyeU7L96XX7GNGU36z60kLn1RVNKq1AJIygzybZzVCk/VeST8N9Kyubu
k4tNQRNv0Ebmfp4FRztAssbVj+RC9KZUcYhBzpN+OikMQK7xx5ZlFuAwXAk2GJpH
CvZqmX1eu1wNKIBlA8OyTzsyRebLA9/PGMFXRhrfdiP4XH1RFg6xYQC7fwV/V2WY
GQpgr3KlRf8pbxmTJ39ZLjUsCyNFv+9aPlRMtPOUFofdzuNb4GVohA+YNRamRVCI
xaFcVBt6DbhrUWaM1ua4V3JeOegEde0ztJxMRc03oy+Ue0PaK7lqy7cSgv+7Su8m
rUrVhSxpJRCiWsK24WQ4D5yW7xHGlHxx+CaBO27YI9gVTQVPArkcqkZMMbporPHE
Ek47wTFT7HRqe1ef1f9wv4wcqclSZcp5EQx7er70l59xX6XZ0jAlvrYOGCHFAXfb
buNlQSOkqCUr1ME0HPVNKWuPs7hTYzaVjuosrF2SK2m9FkpmbY2Keoi1Gx+7VMoc
jPoIdpf5IdbvxFSi7RrA0+Ggy1kAzXdokredKclMJRvJ2q6scO2UEtuaa30nDnrs
Sfonh2tLM9nMwfweDwznX8xxyEVldJZVog90GxBdN8qYdjmOXCwlwVt8LLcFfnL8
x+g4hv8oqvHoEl8gsao8uUn7tOMizs/FHXPKG6v311zSXt2o4YWlRo+K7sTDloQO
HXOVTAs3Bo9WG//VYyE4Vi9vkEM7VmTJ87UljwXh9889YUx9blg+sPrS1WgD6+JU
lD7iDU17pRp8ttN19j5S6MevMjCSHysyxoFiQypjkbI+LqFhA+s5emrkf85v9V8r
o6Y4+jYx7eR08HTU4N4fyRL6BO/HlnY1/IrGsITb/M9OhMSYt3FeSi6NYY7S/J8b
f8W9kv5nz4x97WloRUYRX/NlZoqgwozdiw4FK0UBx7QIYri7zONJPs2A7X8hGdVy
c+hZVEDLcBtpCbt+A36jsvsKKEXsNi8aTxTvxnRDZBrp0rWFyhJab7eEIVHtbM7p
dbZZGME67iLRF4H6CaXBumzF9p3N70Vc/gFyLYZ7WT5F7ECeUoHs0knyu2QTMeUv
jXH5DW4gJEZdnozOQuIBwm8GbR65lgJNOhQC9DG3qbNyuOjd+pwa5XmaPVsHl3HB
WiLrljUMSviiLoPa8PKKkE+iNdA+BtssydCpEIc5TPCDEsSfEQmTUGWawn1w746g
2p+h0Wo161S4nAhDthbMFVnNYvmjqkjJdXQfLwVJpY1dwLk1Xx54i8asCuQ58Kn/
F5EMmHHwbEE61GttBakaQNL3+rByQ3j1JtdUf3GBfmGHva3/KFWFCOdoKJIw4a+O
lRk6Nyfkrm2nYUeuThuop45SPeO3T3L9QUpBClrVOVfBWTPRxKe2mfT3ZJSVDd7O
mEiAEi3bBJvVTJOpdp8DORcuG1eSYA2qHOp949fQgyNJw/yrbQmHZS4N8vfV2pVW
1f2ZKm5/7VYkYux20PoreBePwcSZvsWysN5AxTx7A0FirQnXiqMtJg4L4adgEv8u
4W2LAAAClHezq8TgTKctdRiYN7691dbvDRCAx2pNJ3pAyIdOaZwzGabJbUUxfyYp
eDVs6o6SLfulAUnHbflvc2mXmihmSWqd9oFZUR+6MMFF7ZFdjuNt2/7NIKqjhvlF
pTruthNMSPnJOojVEm+iOAXq0A/ue0CRuClRghAiFTAdSaKnFo9RExWl6QRNX53J
8DwmEBbsGPsdCb+bGDtYSTbeKSYXHDmOnwI1O7XU58jo33y0+2toxL6lIWPv/QYr
/q46iyAuiZHFI4Cs+hk4WrH5oZgoAgfG0LRBcaBdZsZ3WTtIeTRov6fMW/SJHzo5
ShnYg9hyJyzb9LhyELS1F3ywrFXomSFq4R2M2mQdlv4G9Il7rDewRA/dgLz7JmB4
091dpsRTwV/H9vKrplOH9pTu0aUD3sm5mxplxi2RUf6WIRi5sG/vx8qKbiUgrH8t
P9wsOgAIhAODG+OqX6l0/lPXl1961Ij5/eTCbl4klRfjsO9F5/ghbIs9JNi0AUz8
BIp1HBATKJucR/T73zCh5hO/jkCuMxMfYYbsP1Y8eFCddX141MLBUTJdl5VZJIZJ
fhGXIbCO2uhnXSS+S5EV1PV3S0DZ2a79LKN7vMyYsvhaZv15ysI0gZy+A6NVc/h7
vAO0KWzA0xL0GvzjRPWpNMBB8T1OxlfYOvFasXeGbEqXXetuoojISvH5Ax9J6ZNn
wtEO68/eR/1paEainrqTiANCWwFOnPIAW6A9a0Ipaw2urFkFBtNFl0LwPUOjLKfX
AyDQK5GUs9Yi2gwAjmA45wiHe8ZidFcbe2PUp4J+b3JnZTkmhg3BOo7nY1ZfWBSJ
Y9qyamEqdaigdt2YswaxwgB36lZKuUzQAUrtu4TZz258soium9yxCeklfYgOGjAQ
TbwY3m9icwi3+Hk40QiGXN5EosxnJ5vOcbWXk1nM04NEEYwJ2UCPdDs4BSwT0wC0
6NFAb1bMM/Ckh1qC7G/+lq0rrznT/BJVf0iy4n9tQV9jlQBstoVZA50ECoMP1u2V
Y84QibjSPhHnU0ljFjAZJRMc9E50/2rA9G9+bVF2upPFROxyz6dfbitCbrCENW/I
glCynG/+OvDh3YlYexjuybZFPN0mtKYh9QMHGWExXI+l/RZlt58BPxiTyJPQyl2b
zgf10iCQXP5zd8IzZE0CXbvR0178he981N4ob1k+UU86XngFMClltGGsKfk7fPoe
sQnyC4I5DOVkQRloBKK2AuczN0t5NV8/nyMm0BrwfcXYmERa2DYZSyUnRawljEF+
WvuVRifYFnG5jHnFtLk4hFrK0ZUNlEaxuUilDcElJSGdSp+i49pUovRe6/D3uink
U98VsZarjWqwW3ZiMvkk7Ab3KUFjsnxb/xZcEmq3mgqpuDKxZ6SJxOuEjkSTSWBN
nzA20sQuB9FhTKgh/SISblSe8xCROhhC01ZSliULlr3BLTTS7W+qpV3T1C52Wm8R
NDRXItdCpbtuKC8IMIa/ug5jhj6W1gqUtvdoRfQVlHJ3GyfZXD7OzxtCGe3ZO7Dx
m2DSvuHCj6+yHS5eB7OM54xq8TWnP25GYmU6Q8yCfyq6byD4xdJjerS7prjXBkVJ
dIT+g/PDWWFNkBAsyXXpjfWqinO2BPUWyQYG5MRA39seurTDg3Vvx044Pn5blCal
bg1WOl2P9QmBbtQrYzoU6aRHui598xFi74VlJAxb4HV0Rlq6GI52s0GySsBLTdox
bEN1HXaikJTFl4Fa4OuGtCUjW1zXDTqxoSw2HENPOgqJOIQg9rYEDhhBxkRO9kxR
E/Wqb1GZCoVYnG10/SFeky5GQMxhC7lX9fr840YFpb5tdJsFoTq+oJZ3mzO1mX2K
5iX6arh6poHCe1NNOd3+GCpMCeO84v4beeNhB9nwUjxv0rl+ve1QQlSkc8CPPhhe
jsHIuiy8XgTxbrvwh3VEIgBG35uin18OIiOgY3653eSm9rdKQnD3iLhqQCw2EkxZ
Q8w47V9fskIq3qwTjOqjKbHgGuYKULGzYWIHHR/5uqa4PfTvFyvCdzdN+K6Pf+Rn
5NcdT6BN7ImIgKZcBoicv6MU8wYVrS89E+eU41K9wXwIO/uNaD7X34jq28Ony2QQ
FlvuiHDFm6a/8qmvog9sxTJfDjdiEUawouNXcuBRG4vWOxzUP8z9oDrQjCrYe6Bv
09LwjMTGwoqwSGQfGN6vtWtnPpOvEtHkMaTIjZwRPzFwmX8Wx8l2eLzgIOz4zvTm
yA5Onj++7IY0cP6a7CefbkVChgfgOcXD34rWRAuvYAm6cNO5sm8gz6atIbkap3K8
JDVEXjHjZPF8LJruUVepd+jEDMYa3DWoWu55FjHJMJrHMYdmdECjD9vKNx9bdQBL
S6xkNRyPBSXytsahgWLgAKqhUqKT51LtiJDH6qM5xqTeNSxmnua7a58mNw6HGpUp
OuEvumkKEpAeshcROhKpsyUfHNcQAllL+WyTDT2YgEjs0ekNatICgE2hhAkUZrvN
n9D9I1LpIMImPinoOisCWyqh9scrzuwAFmi7kxPPM6poY8GKlnOgrIANjwKguHhy
+2VrLB0DoC3FQHG9y+CPMYnPWt+nrZAd4KskScHQ3Prp8SlLowNrCMr4qVln2KIz
VXpWdc4imbIi0BcWfWg+v6JwJWo+TMhzsNms0A7DPt/G7CNzmOrUK4C0mdXm+j/4
IW+/ndR3XeW86NWPydiy2O5zwbOzxP36tExIUeeVpYc11EBxWzD5HvhemkJ60m10
ybFg5j/totP5e/hGPGGIRdh5NBFShu51QBNzyWEllLrRi/AwTIwvw2KfU+rSaYSZ
S4eMs7M32RlJig/2U4Zd8s/Ng/YaTNxo8oOJzLkqT/9DhqsQGkozmadCNbsiwTXC
vR9d9FDwP7ZLboqJ8EaFT+ob1L8chFqizbH0+/0o+j4cRrjSegHAfNpOJnmFZoEK
XQSQtQRzfV1s25LBMMKlRc7DIKFCFwD1d8XMjyZJK29LITQG7bDnZH/27Q2/SL5z
eylEuKOW3pWsei8e88v3oc9MGfwoq/wFJreWovhVb/g3MgFob73ASxQ01VNBvomo
XUNeqmqOC/pN9yXEub6Eim9CpC+Ly7YX5AUidPQtRyxwkoWJpG/ruypaBf8HUyGC
c91Gv/xLIBaYUEFkd8ec38HAB6akzVdq6A+VHX7T0VbdBaj1ep+0IhX0CCHDZUFY
wR895ICFSeMBuKoIaTOmSJ89UtRvf5206cLQKM5K14D81B3Yq451bl1PBKYhV6Wh
3MAuRTe+osAnHJeRzUjmyFzKHO6+RLAM4K2g5k5mPP8r0KhjUANRgjUJzemasXKH
TDEPoaVGDPasy6k4PFI2lWauSmxgXnAnNPQJzCTdhDWUOSj9TBXsfqlto6OSHjef
IUDEI90Ip9GrEbV2U4O/LPCUU6w0Nwp4vTVv2ETYCcnkkobHntvKCqLBzlbVXiO8
ZfQJ1UDCXhLQWPVo1mVERJbAuSdXyGiDtJN+0U+tmqjtd335hRZklRjsLysQJ2sx
QzRIzu5PuuEp1o0+W8hhyy47ucelQxvRgEyqvp1TPUJ13t6gd4aaQG1hdjQwCp7Y
WM6Y7J528GPwx2SwTwuUi1cKJVDjadhTgLHtCuRfF2obneoHpFqFcqCYTgNBq+D/
sS900tmSFf808PQKVQ6cLARYyYpZSi/gRz4qTFMjmu1NZpMmtTqzll75vUw+w3iX
gfpf4CkDbpzaNfMwF9mC8KlD/7s4eKNS6LuSIXkkyJT27+MoBVGPYTHZ8bmQVHb6
UOeDOPLtw5kP/IGct0WBuEXqRhTqKmFibQQUc1oxp0YX1mFbu+nI2YrW+iLaxTvw
wZBH73ZD0MHzq4i6FrblHXfOmQET+sTg1eAz4p8r5bw2AFKU5X+QZnKUpoZQW2qa
mw1vieVUsUqLOqLJHogxufW9aLHUSzhq0AunTJ6rm1Rr1gM/rRV0N5psBsREjtYU
Uhx0+iK25DPH3UBrtFKAnko29b7BmP04tb+ReIQlQpwRth9Xz04LNL8t5jeS9qFX
OIS7DkXSSUcveCgA8uN3sIYzX/6aHCA1xBaOspRmQryzPVwlbm5OyJDW8JUP/MMy
tIILtlmGSK7/4OtymsZ99ZTsHAHiJTkv4B5Zkh6slXAky+YPkmB0XnfqlkMSaNRV
MONvuzwc1Q5pUVtMiJ5cLEnw7aEXTbS+wRFpImCfKoXai8mwbqglXs7Q99aXhcmq
o5OaqdK+oR4QIRESxgvJH1/DnfvyjeQUTpZrLC5U7pvClJ5CUSvpZBDMJg683pij
kWJZJoqSUSmiQxPvZywieCGdZviF7Z1G8GXazT6vWg8Btiv4UdWtH1MGG5kAm2Ka
3uwANkm02J7meVO5P+UKcUyLRjnew1N2HV3NquB3m7nnPViadDXPQUQbTU/9dnAS
HpiSxDEmi/f99wPkONPDNUWpv7PR20FyEhjoI2he5n2M/I4ETLAekKw5YRaaPTM2
uYGqWoQBYvrUDGttX9G+cueOjOksYfuZdn4MJ1scVulTkhImSWIbddy/gV0YXZuy
bXhgpK9wqd8yX6O94RrhO+PV1LK47JeDm/yCEY36WaY1Xd6fVAXRXIWghU2BlquL
T66n+BD+jPsMnMABxgyHQayMnpydvlZi9JfgJva54l3mRqN+fyjW9CqPvQYmeAhn
0BG1qogOLMCqo0d/S1sb1veG2BJg6h0Mlm8pi7gcKx8Gk8yj+eJqM3luFeR7jwmy
f+Rh3ZT50aRbmxnbjQpnnPq14sqbxJlJAdqworFxHUSohviirOqLd22Yz/wEOXvr
gqA2YqK+maWHbuDsR+Q1S6y6dqgrgK2PX4Nn4hbNMBKQo0B99zUIqYWVug/I5ZYX
/Nr02S+CiVE2HX5RUQPwpNUJ6BG0HcwuhVfNGZDmHR+JxgbFPkAbxXtkIfcm6KAL
pcwzrtzj2O9fKUgWSdBGQB2ywVIrWmVS7eH9j24+vzr0cik000LcYDsuEZo9G0OF
t4Nvjmm+9BZOdo4sWs7rQeCRLRCn+hZ0zc11f+vmMwVm73JEm1V0jp6heq4jaoEw
Xkp4dGPbc0PK3NJhZbwxorXsyJLAMSXha9K7X/xP6lRvvg1X5mlFdJFxrJcRFnLn
ciqhOBt8a3PtZc62JIsfzjquiiKfqE7XMz2C1B5/9NxtQ0k6RO/rFJ8ACTKayV8G
6aOLLLW7YHHKffPllCyv80+Q6Qp06/IuQj80pXvL9SFizdaM+KV7pz8SvbxwEak/
Fa96C9havG7BHvV9Y5LjzYr+G9t82mjyFccPnYLl4m++O2qhR/jMU4xB+R0XTFab
23Ex7cU3Rm3JrYk+FHYM6ZgRlXDyQXxJHy11GQ8NRVZP62ANe4tH+U1uW05xsyND
VyQcZ08WeWBCwnf3Eu9vT4m0CCz7icZnvB+h29AULMWP3l2ReRI5Ywtv6ofLr3Rx
HKrRPdyXd0S+Aw94CNup5tGOoekptmV5G2CdSiUXVQJxxk2PoGU9XZRsSGehjtIi
Xhcbhuz7wI5KZ1Eani0mZC+jpfNGPqhT29T6tJc/nZznH5M+xBP39FVXWkt0wQZS
JrB0mu8z/hhblwL08i6g1ANhgBxjso8OmWy1Shr+X/j7vS19ffkoGSwfPDPHsIOp
LPMLXZhpx1cAgnwcVVTkPjZR2XhxtEtURaK7/y/bUE/bsnWA1LHLUoEMfDSf0Ds9
8PS1tAsun6gRcnRBMNpVLxg0nN+rKqbl0T+kKfZknWg1YHzb65um9Z/5JVN7rf0l
nRvznwPU2rDbM721nT1mcDsgVWrFH+fFJaoXlidavHOPA9SF3/6s/HkZPUPUcIaj
i6rko5YAD0ZXCm2XCOEOzyWkC4Gu+BSSwsOr4LZCX5qAqLJuabU5wPT8oZghW+Of
Rf0fJBKiGVB0c6F4/+Hp585PaZJyL5epHTV1tjmlXnEJp5g07Q/KcvDaB9XgQ+Hp
A8In9HJ3I2w5Vvu5FiQ23n2k3d/C7E5/+s/aMJTFmIHBUr0gikUrbrWhnei+kn29
bqHE+7V6ZqlsLs11nxLsddt7lN2R0yaDKhbpbfJffCc+1ihaYlbEPE9ovWhOztKU
SnA2KzfyPLkKRYeM1uS/v1BHrCzGq9eDSG9GrPz6HAxnRVQaYM98XHLlA3YDX68u
JltcV40Jgitk+U26+iOlP6/uM6ZhYXl1OgTrJ6KNwck21vgI/5S3SH9L2tHESgrw
vPuGJe5zZjT13ThmZVdam7eb8QOwRlVPDcQKd0WyKz8UzQZxwar/AexlPE9O2/EK
jyRPjRT6H4hBSaWhyLFYt3q1a1FOJW+RfH3v9E7KKzz4XGq6ixk1keoQpoY7ciKQ
H7b0a59CZsUnXn/r6hMHzcyu7IGLj9lXzZqoNREaLKbjiAfu+/4+Z40OSN3jauDb
TKBIA8yHIF9UGO5EhPirr3MLScdYOQSlnDYRmfVUA7AP8AyOqe3TcSA4IjLqcHFP
yATsaqPjW8X50rZs0ZbobNz8stm9LZjaeEtpajdgXJ9u+4ZPz3hBmiuHdCVNoRMc
XQN6d2sVPtZAhFGhXDSQ6MoUnONqXXxFmSR8XnOa6xZOjs81OKtgwzO9uNSqqplv
LHZMyuCFaznGStyQXDhN9ePQIsQKVT9A2NwTToF6WAm/XRxP3J6MBNvkpo5nRQ0A
x/iSoE7+6S0kAf007PU5AdxId4yxZU/vGWXks/3EtDkqjOjv+PzvLAyW6OKBKefy
dFD7jJXmVLkREkzP7GQleVIwiAtXI7w+WuMBptIdVkqQw+YTpx3EFbfCZDDvq9LW
zxKkexNd/9X5RATGm6SIUQuMM4lfyAPmFer83yAb+6/U0O22oBpI5cKw7mWMfHON
yJ74/e8c2o26EHGpbpl1XLIYLa8nL30MZUBxDR/3ybbsPi3O6FzIHN1AgGj6MIqZ
jvI9GC4/b/cfMANhN7LqLEdsEhGJJ+IkzGF2XzRB6qdBYvU5HNRMyCPEvET4gCON
F0AHEzwjC3FnEvXJTJ81xbunAjdLo15HbQ06JZtVRKc78/P/e0Pn4CzTmSzz4KKK
h+dQ8jOMxvxG1sS0hHKuHgdNR6Ducn5n97zwiONJ3sLMQr7sN5Wi85FnKJvQvEbU
dwwWsYwF/oy0JIEyK4sQXPhlM5cEcIxS+Pus8a986UtcTQq1/V3SHjTAIAul0pSP
M4SodnZC4/uxUMBM2W+wt7xdhbJ5U3xoS03Lwlvsm/RIohdRKznW1EJPB28AT/w0
XiGJajR9LmsDKmrtQc4nv2VcrYlG7eqra9ZNLTCyX9sYBpC1lzoKLM54I7YSry4Z
N+S/G6wE+wCgkfBhioxCBjFRR2i2xHOM0jdA0/xvDaCB7Qd4TlB0HcKM8tO2Av4d
Y80HJzM+jVIrPYx1jF4inIHg7omkigzwgdWuT8NE/QEXt9y8S7RniCXkByteqXLO
l9ARDvnBs5N5CNh1fWCFKq+BCCJ5IZTNPO3sXX5/x49FWN2sHjGLSpzrZa9UKWBm
HmZ67vY6LQ77oYaoC1ls6y9lsVMLJTHVUeTk67kmV5ED2s2fx2T/NFdDPTx3DR4x
/Q1u9+yCxYikvLkUSGwYahA83Kw9zTYFGR7+eVI1A1ST6tfI1hhglGXzdYczkSan
0gTfQq/tKAmouP7KN/G/P9CBMYgvObvq4cj0AeTT00IBYMKdF7BOk7MGo1ducOQY
uXYtvQKpsZauQ9iPg8ukFp/pMMNlBoeggmEF3lTrOjgbEIUmxV0tR88C9AIH/RcZ
i90PRNifv+UG9G7Q9m4XnG5/tK27QPtD8ojfpmb57PWKvNP2CkhvI88HKFZmsuJl
XtFV/THJHVxzyDWCRCLtbMHzH7aFmIW9rQMPZljt4qkxuhSok4fjRWjmV+6LKlzT
oLvxAWI0f2xlT8FYEyQhgj0GWF4/1yQvnFzUIDsDu6+nPYeQDLthBO2QDHgCubVQ
/f+VxRfwL6//Wub8gaZCHUnuHAzDhF7gRC7Ex9Kpwt27B7Q0Py3NVLU9nP9ZMtx8
eDF/bk6ctgLruJXABW81EJ9kk7Ldq0ZWwz3xvU+XEUsYmthITRRx3H//2sglYzXY
Lypu5ffQvzFfbmWUBIZ4QCqcpetkDHDJeG6rqmxElIHcNX+8flI7yBVzAwc1HkRD
lsn03sgj+GyQQS0rIARzuA6lCEOoGziMy+xss8ki0LtG6if4nYRb6m6tJ+4P1KGI
V5IeCeyW/oJj9dz6CmB6FaqNeLF0xABlNga17pj6y7O2BM70CYbpy1S0qnFdUISr
HZwI9c+b9S+7GAU2nhaovUiNz5s7TM8a89wIa27fXv5Yv9sMIONio8aBaXuv55qg
elPD56X9k210i/QAHjljQ64nS6jMLMoNWUEi4nL6ue8yWzKEBPO87lQsm2Vfnd41
yko+Su0RWi9QX5pzmQqqXbdILaKZqZ/Z6BQGAbGUntOJNSgOh+A1cHo1FEYTkeuH
my8Ff9nD6Fs7SlT6ASRL5U61AOfFDqsYcRbxIgJBZY4rqgfn4XbsT7MI7NZp2Tsm
S8f37FskKFAnO9+EzJJpn9mx47bbCegQ4CG9QMhfmuYmHg/MzDFEhc6olmlTgztg
jSgpT+Btxcec1eYtYDq/9uggQt51zI2PMrjuUwlGQ4YJle7B8cILQvaw3qkJA1SP
1or0mh/gUKhqEArWfYSJEExCc530Bekh1HySxYNi/6hhej/lU9C4XRVJp3Vz0HzF
EjZHLJIkXj6NAfNxWaiqSVIpqWNLb7mncTZrJHkgGBVV1zzz/EbMajmLDDMts0bz
WX3Y8mwdBThL9/jwZwRuUEwnTFGEheLU8ZRwJ9kQvY4hur+xmVXxUPWDZG6F0RFW
Iq4ewkClptVk6Jk5+h7/ItroSGhbu0Tgpr6U0uh4ZvgGs1J4cPQYit0DdxVbugqX
JDz+aVi1p0Lw5+I+80KCe0XWtZIWbisUEGEaRGL9MMX8iY95qG7Bf1pb3Rhj3ntH
QBz9aDPM8bV9kjLn7s+XVCAvjCxwTSF2aAMn2eUWyFL8nxDS3ktWbhZGVZ9YKyiX
hSa5AT8c0g/WYKnvB8LdALVZ1NQX6NAs2MfYpI+/xaKiGwgsAlZ1rhurBOdNTuq3
9K5XkWHwh+ndtATYzHaVUSIy7s8Emz75dn/WwXzTdk2LomUQHFInv5JqDDC8ut2K
4Vh57Nuv08I41q0fFZQjL0q9viWTMyWU6L2klGDdFmfsQ3lNuUp0TOHFdmRJKv1F
vIW7zci/XrVe4TkRdfOApYwti8mmExoH0dG+OEo8CSO0QoLwq2XCN/CRw0jKeIv+
aT9fR7XF7mS7Sz5fdF8Rs/58JFyrnMqbnyTdZZbBwmsZuuzZE3EKEpvuhjH5UAxE
Xcu7tCFqBR5zkKlBverFshXTWl7SvdH/5nV0RpyI2vD/ahb9muQ08DvK+469ynOM
hrLfR+N+MBL2WcEqdfrtZXeErVtrDFFiggC4S8Vun1zoMlZbaxy3fJG6z6nYqNs9
EQyFgUy8de8nCHr+3BBfF0YItWT8nQfA5599tvxGHIMNRZQt4l9oEh//OEHyLdcI
SvDxh7sUon9yqKza1Q0RnFU6/4vPycQ2E/Ik1m9D2eEwAV2ZaUvhVH/R8MWjI7Vx
J5ipSo7JgJdZS9UEePeh+PIJcdFen/X3DTUoc9+mSiWbWyYlyE5Vq/AW65N9kM/q
rNuBqZJrMV0nLvZJ7tGf7VGS6Hy7Em0vwUVPI8qE2zyHPExBlCDaFfP1vYWNf2PZ
LcFc2NHqY3DcXEuONv5aDVP7xQdiyn7Rd0mA/3pCjvl22l9qsvBrs7ZOACcffh6i
o7QMMo2vUw+nXpRwSVjUWzYkK+2PcnG2Z14KWRbuxxrvAiQ8yLHd9PxzjpyZc7mU
6Ou09st6rDdvMvYMIbh4SEkn7fGsV7qyY2479NhvNH96ZmwEbA7k+3dYcNg+xgvt
IbKZI/eo1q0mWg/Dc8EdwvmRZZBSaOVBoNXq03ptbpsgBkFBPpSOrRaHOmeOctek
8Q6eLqNsXFz/KrLvYVHwLKohndvG9afBBkiEfQw0Nr6cPmv1dEeKkHI/Yt7OsVfh
68o7lyAM06d8AoDDnxJtUyB2OofrahAzMEMFLyya+fBtEK7qutSJOMMeuyOgBW9N
OfeuBfzK8jiBTmXcwv2hXwfl6YY6lIdgyznfarChiK18EMMlMzLdtenXkPGpuHvu
3TFT71OkvCpiPAl0yFU8Uqn1fmlOOsO35ImAz4lt1EmZNGJ3HnuUyk11D/RwIiKA
ZapOyCx7/VjHRzG3EuPhVnFij1J4Y+If7MZNFZDK7kXGI3ffrzafDVVcuxgjXVON
ql8PhD2HRH52xGDvtWJ1kfYN8jIrog+Uc9bK54whbm3wYZKzxLhtOJk/4MYRFDrQ
0m6LU3/Qy7RyOzKUNxIbdEf4JvAj4RHrOBviTO3e7E9BXQit5RWsePFqVH6seCnm
fjyDrvMHKu6OvCJ2VDJhewLVvL8BWxcpSllJsw3Ak0J0fPhKvxh6T984QtkmFj3O
0ljslr0tc/vw6FTJxTokNbaKfi9+EdF1ZQyc9w62VOhHAtX2YWto+LsfW4s434QV
Wy0j+RBkCyAkUFPXtmIrxKddM3SlWgslGMO8A9R+z+FJdE53G9JsXzn6PZyHSDdT
ftVIPIQopwcJw6oryUnurKkKl7be3DRMTO1M7sc/dJSajteeAyKVHOjveyKz4Ob4
r3wo9H0PivgaHdPYRj6BZiS6p9BdNLWLfW8S7dFZcHGwSQVCJpiWbVnK6QoAJU1Z
jJ1S6q24VXb9PRIfuR0GDDahp4YprBfMw7615x75o8RGEYX1GdBBj7V1PytLjCHz
w15AfCG5675gvAp0pWvrlIELsJASg+9qbkICs+slSVx7styL1l0edQv4Px/UyCPp
hasSRerRQd/jbDZAUBjS2VjTuR5XWILwNzJZODCdVknzQb+hU/3HDf+8UzW8lNPE
eQk/6cXq97fsd+OqELixUNiBjpfeK/exqPYkbKrP2V7dYFkhhfNdvgNeFJ8lLIq5
EXpR1KuePNwS2KCs1nZ+BICuD9kWxNznBl+JxdMTr2HxcpFoMTXEfmGeXbpTgFnm
3l+rf4+kcD6u4mf8l59ErhMxO4cy+MOIPRP/F3LUBNSHJVoJyRK8S2VR1DERKYy9
ssMAEiazVN/yjVFRj967vzseS06k/dFKK2etSDvMha82UAYPaBFmMLp2JCQ1WoJk
30YVqI35c5CcR5G1UHp824VsvLtHbGZL03PCxljlOTfssk1qvavDh//ALN0UppPp
KtINZfGbdhDtLc85rf1EFTOMWu3duXfCktJ++nYECgfiE50R7nmmFDe5ESkcBjcX
eGTSruz0epbCBTbK/nTHA7adMZhecUvLIetAJYlA4ukE7SwgcxWyTfXe3egqmIRn
TczEP1kZ1NdQOrB1XWPkqhZbhuPJEsly0+mXKlJn3ce4u0PBkmiH+5ut2BaF0H4d
jv/SQ9HwIzjAqags0NracD9nNej3v6S5XANPHvfUGazAAyhp7SmeoUZguX+MNseU
OObkyWwOBoQ8XKEPDeHFBZ0vllsaFtKyWLzATuf0s/TRL6rf1tDGz7HwDx4HlA1C
8d0fb7oI22Ttle++IySpLnHBpefeafZ3GCjbLLeR1HwsM10Wu6uL10ExkWzUk5yP
weKDQFsnqlcj+bt8inmdK5yWATbnpcV4kAfY32bDzszFr6IkWIuPPxqKWC0HAeJf
vxQEsPL3e3PSAZwj+YL+xKEVS7uCsmH/u0XOUrRj616s7AR9Qz8wGazFOjCOnB0Y
zBxtyouGuv2NyMcW2zBxrq3tTfF8r5zVdi+CdWYhw2QYJ/LiauIseRn39If0bkes
+UHDDNGAQtPE6THvO3FD7zn/uX/AOItxjXCAAPEwu/mLSldYYhUA2ojELOyZW/83
ObvLUby42vAdGjlPCEQj8SyGybniJDuHUkLhYsazmuhYvvfJhnQBf9vmii2XQqJB
r98rmpsTMpttKAqVMI1Uhns3/0CUwqTkPo0EgFIf/nKu+g5CcxERowghNomiRl1z
il9PQ+Xd8m2FJJqdaA5Anb2IEggHm8ODEwBxbiutHk+rlhtX5jg7PTyWFC48/Ryq
WfrgDLeush2eS30ud/ZcsU0dgWa0Mi1/k9EnGQbMrVV4vnwF+7Vy5CLdGgdScUsJ
oeGGNnWi+0zm07mRlsoAoKlWxKPv28mn2P1yC98NmbsNb9GE0yl3GsciSbTQYqVN
tuo7IkZPouYPsldizNfso1fWsbaFjkLPumZeDo7SAz35GK7TlZDER7twLTj2TUw/
Arr11bLQ2sDdJB9DO6FpLF8AS1+1OqBSmuxPiRTyn6flDTh44Oi+RETLtaEAI59W
sGqnqLE4xspaA/KhzKh/r2CJh7BZdtxeIVjeHEKayeNJKiyBHoK0ileBJpNwYuJ+
o5e+H7J6M6p1bkr1PQztZ32dl/fLN1L1O01Tv8Fiffho2qqUc8fF5HeGz4xHrogQ
SfEF7XI1KO8F9oDJeHZBGHbUPI5uSxfOuHVxAsp4IrvKOV8ulnIX3oxVGq9Be7Qz
KUYFTcdLhvN1hDHR6oDyEuebg2aTYIzJouTv9RZP+d4hEDjAXUqipUsx6IPtAS5O
g7npavxJ5l2PnOhVlcvBRdHwJj0vlM9cJ0lMEpOt4TAiYZf9qClXeLtz3/EChZiJ
TnCcOvRE5OzGN9si1gVao3u2VM0/zW8zaB+w7laHVsGlaKXdYtvktdHNmuD8acZn
CR5m4HFm3RgxcJguWN6SIA/iigFWHRd/sniJ0rQd68WXvNNgzkWG3LhdqgVdOWMc
XaMyItOKbhzmC+RLD6oX9PY+aW6h/7AcJH0wLBriE/YXkJlRyLJKTgXRYoriGAHJ
ZRAEMPqbVux8mibKS0G2RfOd0cp1RpSNYw9DT/JToMV2kg52WvBo8ydt/lGJsIfu
l4qg5LhVoMXcRdboj40ak6YmJodkp2Ivp7Ar5/Dol016H88UYz8MkU9RPyqb+Ibp
voUuLQMtre3Wzew9VDBC/6339raA4CYz4yNNE7P9AU5fvty8R1f4qwcT+kotd43H
YvdqAv9qLlpisIActTUmCA79Mmk9xvRx9sqEC/ae/rjs/MxHfKXfqT+E3lISkdQW
3EX1YuYUAcJLOGmPvctzDbGdcea+gOnfJUOrPdisJPAsIy4kBXpX2K8LL/o30dCV
7LVbJCA272DNsqhMjyyNbofDbIkwEczISqts7fVx7n3kask+4InstAAC+tu/W3Hr
9F2aVJ9/+cH0ZVGzpsmfTLfH+AiatbKPhkJZregpbMsKuK6Lj5tLPnYNcpN0t76D
bI+vUyB3CTnLzIU/cybYqGGucsUDEq6qOqYq34Q96wD6KNMpNqk75C+QoZjiOK3+
Ag+lo6nlBTGPcU5hpPOyTUVua7PEojaaLV+4bOrF/8rXaoZsOcixyyszAJoFRxyL
B6s2AWYV+XQ73D6SPscasndGSUaY927UT69EUORyuBOLe7Hj+3Xzg57VaA2zFqK1
7AiFddEHSTAFIwiu6fHB11xcMGoUYY63zhH0TkVJaab5ztVb+C+ra6NvIwasksaO
3obC2MmRkYdH183wcpw8OACZh4P/SbH4SEral7oGxYTKMER7/XslH/6EJtuoRMEI
S2yK/q5DLHTnHVeEPZVu/6CuTF+EICVrtJaXsw8BzjyhbpNsHIXXd98SqFfpvSt5
S2PtjgMASar3TBwxCfgZV+FjSHSSoUyu1Z3Ilx/t97p07Mr680UoV7goxNQzIoJM
hVA3HEbuOcqes0nD+whXfTT+24LhsVnyALC6x2Ly2zoiA5lHK6++grCO2ouJ3daZ
UON1dESMRnaHJ7NrhhfEsUnDQcD3+Giz7Iewv/8Wv9l5+eNqA25U8tm+G3V+cQo6
zBFGksHjUuTj4sSJvQ1KP3rlZzwsBlyt5YV9URhhK927OVpesXBgejOoPVxj1EJw
jGgcajK4N78tLgteBCF9mKx1p/ouMIDZIRx0JfzBsKpcdXNI2wuHpJaHLK2LzvPu
dyrgoYYy7XaCGdCdDNY2JL9JzhHi24uESKWn6pYRmvL8B0+0FuyYbQM6ncvtGNAd
+kbNyLGnUv/yzyzjWOYR7ItxmiK+zirusUiKuuX/09xeyqUIIcDoKXq4p9+v6GZi
3gKTEU/lLD6w25yZCbttmsobUPzNAKPyc1vR5xpnPE0GLXHsjng5gS0kY57PSFvJ
ydULexr4GibE5goK0WTNjBzUOystpSfzDlmo/y/iCCrMfEkZnDAwrWeUfOd5nFt8
IiuAqt4vzWvtNlXqay31f/KLVeRaqkUhRsfZ8EIlNX4QV3iTXHNcNL6il7mpPMKz
QgOJf7HP9SkUwpT+pBwbun8OeG4Gb+3X3Dk2BzoYfQUq0Gb59S7O7zzc9y9LFUFJ
109IcdlyV+M0RS3zOT57NUiNV8Y6XhcgNq0DpbQhASG8iQijsqU0wZldjS1r1zPt
eN+CXLrvWzprZyqshZJrAqvsJock19HQEwYfsXHv0n2tlizMJBNz76c8Tp8TMYHY
m3bjjR8uupnHJe4L1h2i1eXVrR/93BFw3wXKbBVFYMsIvF8WUnrPINuPZZBIADj8
Sw+4qv1Rp38ZBK5SMxoeFuq6CXdmCAtCFWxXbmNseshlHNy2iJ7Cht48sYt/wNqe
+U1GTjiMwmOnofSVZws2/V3weUr93cwy2qQS99Z8L6pEEeTFvgeqG8+47TjDyCfo
6PMBG9+47VtXxjeON8LRfCrq649inNzW1G6KwHE/W4zH3XaC0bTI1nbAgXIcfPyt
9k0ccXA1q00DhB/2C0bvrX9L8ZvB4SKdftP0uSy5ziAW3Du7ZKb73XlqD+cj+q4f
L4okj7B/fQBSQ73lNHAgcO6nya5MAetSd58+RXYkpa/SIcR47nYTIUJRinTqYtuJ
CJ41mv2w/mMdq7X1YqxoqS0s2WhxrdozEpuv7EdkxlnvLmQeKJ+d2XeosZNupAmA
04Bf6RVa+N4PlOZa+0vcDF6T/2HrYlrieroR6In76WqbgGvvkWQ8kuRbLucEYZYs
95FURHB90eHZploEZBVfSBs8Iktim/KeTydfk7FyX8BCAQo8+KK3LyQYV8n/TxAC
x4jSWgKbJFWy9GVh+vcpxUwy4uL6y9piJECwrwp0o1T0Z2rC/Y7zn+vomLQcLv5i
jhpL6GMSI749fwdxnpX/LeuhwmN8B919zwPymz/UVv7Kt9xjBVFo+arAyQMC00P1
LffXDYyTE4ofFhBcYyqcmwXZWmHFjtqvJ6uIMn5PPVcpFTQLnc/2KBmfyIuICTur
UfnWgLmSU7UCdB9RBHTFx8dZ9Y9cWSzH0EzIi/hpADJba3zOi0sFLzqRkCvPwIDO
4LdHw15eCi1HrxIcxv6dPjI4j+k3Pih0UzuTpEhT2+p5WpZM/evnge0huOQAU/rT
235kOqrTb1Wq13Ll5FK3ofKEPTJHpfFDwYME3fKulVGh8RIuD462O5PwICEiP8Tw
oamTlKNCYQbcGsPhscqMFoF3STId5BZvJ6PAnfya7ktVokUuubH//29Qjsk9v8CF
+EYEQTSHfPDMInyieDC1IbHWOvMPT+PoUcXyPh6KfmArK5HYFbingfyLHkXXZk+r
3DBA88TuxuvWR87DCcIRNJ02jegeT1VV6O9OASoKZuS+cDldSbv0NrOND69nHQ1O
xtKqg64mgJmcoWvo/N+KkO67PNkf+fwwxWPMyuDoCufdThFgW2vFzRr7QclMYhEE
7b5y5iLShn89MO04IFmbzsh0Q+O/4H5FC9NqjLyjBJn9H/IIQc7TS9X9sBGbHS/F
3r3AwaRsdZgYTvymad2K4tsDtRtKkgqDpNOv3ygnVEDYtuuYx5pXXQUe62a8wsE2
GgvQis6Iy840RJsvGDD2Ko3LWApBaNGcqbaHEodq3RziOjUqpc35HJl6jhUPCXmy
URE5WKjh5oDeJVLjXgW1Jx6Kl4AB1B/8g+H3YvnlAwgmTeOBFpDbCVeM5mnGmtYt
KlJG0AMredgKDK4em9l/6Jl4oXzF2WMJbdjtcbRo2adVhlJjBU3ES+mzhPLMOd4K
Ul93JnMj/Wi78PvnfYoJJVStfliF0+LKAPSwYA8S9FmpX3kYQNlTe6B5kn/zXGe9
L8Sgx6RWr7Gu0P2gUQW6bmHhDjHWBib7AP1ATORs4oV4s97uP6Xs7Vdn2fO1ZykF
DFBMNFqFqBcb/8OmRgY+RQ0JNbEcFvrdiNHeQn97xGcgkCbPg1WNao2XsJFuLPk9
yEfBT2IxDrO1RzG/fDIOjJuIQsjFCVDxXzsm9JEYsnkZ4gIHeBsyBqPzH8CB2t6l
iw+a+cvJ0BacYCxI4lLVMmNLzptL3Kc0cPSpL2cmJ0Ot2jlbOBbjIWHOA2JrSD+q
Fflyy0JpyR3nuvy+eBjGSzKcslB20AfU05FS/+6G4+JSNIEdS5be4fu5cj7hKPbl
w+bb2tkG6Rr4DZYyU4CMoP8tMeKJWF/pfwi1uBdMKjycPo1CLiazu6f2b43udISD
UkKiBue9V9EAVF07DEo0bocKqLJnm6tAkxNYJ6Kv4uwEyT4ilhCphRWNKfvXoPHn
kEofLdLCyY8IJS7UKEOn1zbnrnLDW+/3Uii6nh+luIuAK3uC0V4MjlJLnuAYMytg
YxSIBiwUzZAfXHODFw1K9uh/7XgwreUDrCd2C7cpsukLaTvuLe3qK8QD3ZJA5RTU
Avwk83y/tvU/5XJKGe5eQ4UdFMys6eZfog8wuQIWmtFKOckf9SdUq2BAwU2MK+MN
sSbtSWFg0TloNoe1oqomvZFPf54OMCZdKGO6Ot03tXFly5id4JgKW6u/xtxiZdJK
Kqd7Q9YqXXWyWVzOKIiWI4yDnsPhW1Ws27FVWGCr0xc6ddJiTCW+n4ktrl6LCeFP
5CMfjT0P8E9rTxxsgLaQQzI876g6EVmmIjYx0hgpVM0VKCvHhzg4ltmUno/gB2p6
npocqGq64q9mnE9+hwuoNiOaxA0m6B12C56B2m4ZQXvKSWxKdaz0rjCP3tsV13Vv
K9EOnFwl0Pf3Nr7uo0eMKdgtdGpeBa2o532ldVJKWmWh8E7gOOBaMHewVNEgJsj7
tHl5pkPxcTvlGSuWPVKwx/s0A0SBzhjMmapFr5ltKsaOK7mwQj+XTiD6lCuK6dLl
7J08tcjma7jDCFTxolAJyy4e/oaLbYrP7HfAdpALzfsObCoF5zUvk2BwcKplMRc+
B2386EGS3oLoHHh0sb19CF1qKlPEh8Zn+VYJSfP7hYzhU725Ue6i8V1l82HEai5o
3ZbkQ+3hVwQfJ1C34oflg+1JG1CnWsDn4qo87lZOEawRQ9Nne2NriG4xaneuOp+G
MAC7OTx74X7lN7kST9pD4eu/K5SSD7qqLgP+gFBMv70AQBF1K0Yye/UppSTPUB10
lfdi/KdLgNVG7C5wJyOOtcBtoK3PvNYnZxAZEWqskTDrpe0WSAHR1kljOnk0JcvH
Z66k1HI7RsEOyELDwSQpSVzcT7slUycF6n/Hcy6h+t+furTeXCqyzd78k3JChKl9
jfVOV9AhvhVDVEpMLQ+eqr2tVDivzyxoTpoLhycQxR2NukOFp4PREPdXHUZhduOA
ZJJqygN80vmXDjWUr5YNy1FhTBXCxAv/oFCwcRPaeUwoGJYFvqmYjWZ88Sp9qsAl
1UcX40HSkjs/fpVp/4Bg48WgYfw69OAAwgcolR8dVQr74sKAw4+MQ5Jh9YgNDPGe
32ck8YLTuW3m30cDBmQiIcHO1U/+2JQlulUqrgQcjvimk2ZVvmr+uxVB6hKnhgDW
xMwTW4IZv4HL9CwdEn+8XZrGUx1VNThW/laijHxJAnzpH5RvR0t+4dDtl0i4Lsau
Ou1ANPofdiPvD802rZ1wONw9BN5A0yu3nZpSPvVR2JC4CVeLLFPUJch6O0QuMMm0
9Dih0IhwYfvWX0GNY3aPaJyGp6rgVHEmEoNj5Z8fJXZUe2H/AbdHVpZAUXU6nzL0
WCVr3u68hjq+YjT8WbU4pdXKakNk9vLUEQRtGdOTUTwJDeKhdDUTqMkQTFsZmlWm
UBdFaTIdm8yLKkAZYXvDQFFTGS4LVaytQd20ANGx2VdPaEBbCducRUnGckkM+zDx
Axm35Epz0inCDyxHh9RuMj9PKr1inofKw25AqBNTgHQjadZPLb/wTluc/mPPSdry
MJggPzcorhf/mMtgwuMxFW/7i9iG9JyT8u2/4nEPAs0rvFl41NMPN5ghOtmFNNW9
wPeDPtq2BtJlvxEQ8ehEAeloNtiRR2tCEySEdoOEf8vV989zShV6wFV1hYMCbGmX
JfkOcw//sXSuhpSzLXNngQYRIWm3KIcrKi/Bvg9jUyE5nweoN/jAeQzhiDXGFx2x
MEkCrZfwqZ1oPRBgxWA11vfYms9iS+O+D0c2OsSzUA3rDb0zIMZcbiBMe6vgHeA7
jivEcgWM8Wl2vaLVUqwt4FDls6lQzrLpzcFXw7c+t9fgL40YuncgtLxrq08sCL/b
hm6pNUBMuL9ivqCaGLlc6R7I2wh6HRd4u3v8GCnrFW8oG45Chq7kUsfABqrUhXdk
HF8X4+Cdy3NsRMrXTl0YrJPpr5dPb0x6u6q5xu5aaPIMXX4i2UnKwNqGEYHhZiSb
kzxjKxaBudEx2QrkgKDIrtpMrhLITMDO6nEIoUK/tv3RRxffEx9R+GvoncVuYAiu
EXC47WC7vAqD7M9fvTqqqYtKbL+xgUeY/ONo8fxcpc2mEQ1iAcHpudE3uw6ZWz9r
DIZA95mYtQ2ML2/5jFgUL10qZ9e3LRmbRfVcVDWPfxebiVWiYWB4Jupa6SkgeGjt
HA8yxeTAkRxIymcifTA0sa56K9KyZggWjf5PCWmTmsv59nzdRE1CIZR/yk26r4RI
tx1togpLvNsJGAZ7RUcBrTn5JgoBdHWCEbyghx4biL6Awt3oW4t+MhNj5hM4JCoq
lvMi6Ehne+ZUlzC4WOWf8bNd+vSuOWaLholEP9+VNIw8brrmUABTgW+fiZGcUzX5
ud1zKnTIilo9R+i76rj6FbKxOiyziUubtg0ixyvVYtFNIFHrJWg2k0JM8jQk5NJm
d0cfUkZcQqs6/BoqKOVmG0SqzFvXa0E9bp8o5ZmBwB4dhEyck76dU0NnADa2TIn0
KrJrIny5AO5JfYWErWGzCkjl5/w20lAJg5SFWYkON1kr8WtQ7XVpqIqL85DXKoYF
qyVA/TJDUwDicN2TqnttHGNZNA5kvA7sjnSglyWqWFIbqc1/L1dQqZ4YYXsUodPN
lwPgLKsEv7jruWLZ2dQPWnU9QFiXSS5HdHGYyIgqPh9SFEwF21bxa6dn+IO3fqzQ
5BbPutiZTnpERiSMTNkIhUuEL3geBNbbdkTe50LiPB55H6x0mQin2mVrfr7woqOZ
vLqujz1Rm3spCmVZkYSnQEszh+po6GRpQqQzH2z5k7gAzkzApweSXXf+eDTDCYfw
CE34dklEubab/tBN7YSUAzmLlUv5OFVasKjckwOuK2qErtCZB7GchpNlgGaZTYJf
JgaX2wD/++440tgmDtIRjffZonXfCcSfnZPhKe6tYodCmtL+G8XyUmyuX5+vf6Ui
q67Ld3RFR0k3o9vrFtE7ZmaZTB2WLCjfaiVkwjYleqO4VEMLtj7XtylmINs8HibZ
vgWOFX8StQdpr+DBRv+ha67On9oFrEj5g0qte4vcWpKJ3vGZYup/juBHTHgvF5BQ
Wp6sOmljaKKYKSEif5lr1GTTP0JJZF84KR8f15gRrgj+yNySb7r1SBK42pProI0e
tsYhjn+C3vTA7FOExqI3aufGc+oo/QorDaDI3TUpx8ZceYTDoV2OsKhXEE4feGMY
EIN0vypPlDZx241zadg3o5lgbtPKO2rjjJZifZKO4+12lD4p6EVwVbWsipacL3Jl
1ffR+OajH2fC1n953Sav0+Qi4lwFL3vm14PhsURRwgNnLrnQOA9U3cPJpfyCKu8/
BTae1+NGXkmLhyZ+gUWqqT2lLbc4vU0J0geKtdUVbCo9VYU3+kRz6RKuZebU+SJR
zBjuSPKhYTliXsU4WuU7ktNRt0I5vuTKhWjQ0SpT87bqv0Btp3IdlfA2FpuTBr6+
3y6lC/bS5BL5FnzDh/KLdG7IHR3dFrrFQZSy/ELxD9vQBagGdhrzQD4hyCMlg0IY
B2U1ma9caRB/ia7FDvrNHG+/Kn1jvBSeyLoN23jciPY/u8F4eOxkecuAyZFybbEM
rdEcFjhfiiohS7ZgKpA6LZUQjtUb5YMyikOwgshwxpmuHoVgb1sFIQIMSjAf8A+S
DQhnbexGnThybExz2QntoJyAnQbGa2wrIN0lSo8ha4E3YKfMoKzV/SRaazVcWcnv
Vq5kCq9NkdYSAVDXsipoZqfdbiTQAHCNkR45uBwmPIAt43sI1boHaEzXE0Ru3rfb
T/WKFb5WAsKvImNKjzPuQA+ecWp0hPPPWFp+1EMEysl6QfqdAXIaEYfsIjHziW/4
aVzTTr8HO4UOXqTeEDBQPfwKg4QNIUiZAGN4MJs/+WTORng79tdIGuABP6Btv5NT
GBzkL09zurHdtFsXEq8abRDPo8oKo8vEWS8DveWXaOqpPpmcrEWtJmljxA/A8/8C
cOnP92P/GbTRW+w6NTyABMP7eljU8CynIjLXd4XifFn7pROYDcTrX/KK3Je3jExN
1bxguz8eI26L/KdpNlD316mSRnoEwnG9z8imsiyyx5EE/tqlHyryuZPsdZqqMGEc
4shSnaKFlK10wI9mtdKwxwQzN1hSnJW3kv6dh4cox1iYyVTR42ZISgkNEZk9ozXi
JD3b14G2KdGsoStQJ2IImLABTpgUl9yNyieTxj2BPbMug1DI309ufueJLS9l2EW7
E8Pp8s3JBOVbzotQTVfQVHQYGaEn2yo1Iqe9uVtS+Y1gi1bO2WMgp1eOAcrlwyUa
cppnzS4sywevSYAa8ZGSW8LNqr4Sk2OXxLHJGXE91ezX21xEolLhby80MSAYfugb
tH0JcIIBAGFSC/bIw1xix6+Rm9AfL3Lnl6OJyc/FYXPGtoffpYLZ8y1jYxKYOnqF
voq15rWzgZkQgqTaVdDZMvIRryFGbweSToBHXKr2FsqawWv+0k7+2bXwwY+b6D0p
EQt3sZGe2F9yT9kqukcUKONqUwCn9DaYKnBdcedE9nECXPe94fhT9l0/J2DoyF/I
6mW24x0xRl9u5ucdcNODvCoIPW5AZIsk+jApKFFzLPySZ9p/5p2crWKMI8+yg09J
CrslV62mXXrVoGsIbxgeKyfQEg2Z/1b0/YBLrQUmV2I0GlPP20mUVgh1NGjjGwBY
rG/ITjDRnl2izxff6DI5rBiViKutC/3ZbFTZ75VRCOOJTwbISOZrx91czaiWlG/Q
lGCGpo4Xql0zvkVgozpXZ3ERH5M+XECQduKHaCu3RApB/R4qdzo2MHd5tzi86qug
k5VtYIQ8rPIUaTkhVQVZoO9v7ZCaAB6WXUU6JhuU/if6GiAu2IgLUW6FAp0rIBy+
srMoinBdGqE91pw0vype1XTF229m4VCBlkVUWjF31QgihHJf99I1n/xYA8OA2Q7c
ewavXaHsUUdU4dOHvK9H2k62AEQYMHMmHBERWNihZmo4yUQ2oGUxvbp+kAC4vltp
7rPFkhtWTip05EQQ7txt1qGIqG5L7ehrzySXR7k1ONbpU0Ol5PNZCfTIWGAEmapW
61gEofNr/6EMi1ZXdt34hpSKRxBp38LDk0Faos3icDL8s9jcTGn3lDOVK13JkdU6
oZml13vfBXcpFNoJBYuMMlmQVybyVWczdRUnxt+C1RxST71GdxBHgxOrjqOcqZwS
oowlyaHtfPvYBe7SZ0v77qNbeX1r90iTq2+THdLhHcrEc7II4J/SlqoHOk2znVMq
pV+kaIXwQYM4GLtbb1M1SjPmMcx8lpMgDIg9sSjpXvNthAIz9VME+gxwR3dWBsLs
EaWzF7upVs2Q4fKve18dXtAQ8PaXDzBf1oLtW/Z4gq1dBHrEtGRELX+7974mfLDB
0dS4BeFitiN5ze4u8fTSVQ0zMQySmF/3NcHyWU88UHCGGcxkEi3pmupFBj+mpnKb
XPcDzxPW1ZZQVRv58Aro3Y6Zj5di0YNzfKkDYULqqlGbI8YlBny+5XwoQsVA0lsT
rBYApjUQn+FOn6ccKAH0NuvQSqc5skuDIIDrHnbEGovwnM3w74xbdrNq4q/CLBg6
20u5BkicUj8rnnOQJ2vZuCyjTu89fzAA+8X+RDMRFDdXSpTCMIG4HrQah5e4o+iG
qziQfd5mdih1Ee+vmPAiuNv2muwk+GPH4lsZCDJz0Z1IWJwsm0aF5cX7s/J6kLM2
02mjhUQ7TbByAT7+PciV+FbiSgmC/MnmIyOSGj+sAX1NMXW/I49YNqqkUJIN26tx
IGmEZd/EsLhRLkRU3rqdzU9bY6fFZK5GTyZ96MH5OFbcwmWJPCOaX1PKHT1ZqdJ3
2UmN2BvFKHEGCe8i3I/4hjGNpdIo4v1xU3DcI4tGPuRQd6ZFt4sHV/L0OK9GaQeC
7gQ+BjffE1wnmG3nNHAzvl4G4lqwZY+mfqrdIaP2crZQKnogUJQa9X5DzAeZHTlN
Ht6yuZQMzIlR8ZX0XPm8vp5wt7TQrYHYB0sre/xIluD09gImFmLKfBVHzeJPFZdY
/IVFGE+qwHLNRhdZ2BxkClOid+PG8oJ5xDJrkHS2eYs14gRMe1z7EQziE8ZDi1/+
PCQpNDYdDKAlV0hjfowqNl/o6oIHLwaAhXNbhRNk2VvUEmCmdC4zYNY1B7qKzYHf
Obix+R4ECoTDDAnejbRB+9PD2G91EENGk4Z5jUfg1Ghv2iBodtDbItQ07yKKHTTW
UJMukZa+t/CbXWc3dOebrWocrFu31EBf1cEXPXv5A7e/dTq/t+AtLQqarQa0olZ5
Svmu8zCPkTwcPJ+T0W1YiqdU7TEhbC/U84RXBPynbW/d1Z1IpfhTJorryfBVnT27
SbvUlqHggJsyp9soAY0h9nwVvTMlO1/MutXBnxOCOvuZaeZsG4lTXXo0YuOPDBRW
PmR67noLImUctPfVbm4PuYV0nfUdajrzNjFStaq8r/3m2tK/C13vvsMrN+MsIVoP
ZMx6iKwPRhNc+MhVjYKUVPA8J4UDUSwmeYlXucNJZWFp1cCvhFIlNfCdWyXlxf28
sYkKQi0gYU3LICIotasr7umYZkXqL5Pgqx7EkcKRygBqp/F7yK9+ufaD/oWXdXGp
k7c6zv9SnfdypK3o1nTWH10oQAotlKoMSEaT/YKTy0V3x0VjDUTWQV0UAXMwgtrA
TCLWjVZWCh6CCW9A5hrYmPAcEJYxHlyMSffnHuZqvi//l8QQAvMajb01+v4jlnPg
TVg88vElUe9IvFKbJ1W3Yxh38TBDOiGUOTakzZGPvo1AuL2UChjPojRxg0Mg4AMl
h9AExXUlAaw3YZ87cDHrnIsTnA77YaynAuFFTiWrJUAlhn4yaZ4LBeZ9jOeRQJn1
8BODz96A/30iT0uTnG5bZOK28lVoQhYh3jLTBXFSOHRhwp+lMPkQwFK6GeQkWFsR
tM/Znck/B8EqgVjD6ypeMGlMV+SU4pLkI6AjCaH2sbbgsSwjaKf2eJjHJcJ/5qyG
9zag6kL5FrmlXXbF1TT1EH1Vf8v3EZkSe9GmgKfvPSk1BfvC4Mqut1QXLJZf5jmy
mFFNc7Za1tV0gv834cb5cMeSs7n62zVH1OZQ1A+cpeNoNonbU3G8/T1cr670mjHV
6fYYpl4URzvvuq00l0YMxMHpJ1Tz+yBW9YTdB/YHslFN8V1Qxh9OERFFSY04Aqlv
ippuTKuXK5lqnGPSZ5As7CHbmOiLULPzsditZkIDJHR62WQFOEihMggEEBdks0tA
gI8wcSMVLWvCoiD1lROD9V3fiKeyYRAtbLmWcFvtwE7yqmAf86sX/BZAaNXjiWxd
/bL3iB//Nmx5DJvqZLWlcp18U+ao0BnMmCLY10ipHiEF/hkIc1eSWRqtZZDNKaPw
O9/iz71JUWZxgRa3snVgnFxA/c2Q39gL/DWgNVAGrM93PnNWLMVRAgPj3kh5+mLw
AH3Vk+oMm6lXsP5y1ry0soH5qttCErr25fp3cdb9davlv4iYOiJjiAKPLxl2OHyy
ZkrSwwDSyPEhe2nphGFE+2wR2gPUG1gip4hwmax2yQq0/9Rs8c9mSHfqzIdQlbAM
e4ac50Tp2Stzo+WnJKcMHGe8aqTJfj6jmb4TrrzdH/fgo0wJVA/seIzMg9yLylnd
iLsJ5h5avZUhmToGK3q3viZh8lcp6UMERSA/frWMy9D6oC0Sl4paDjjbGPz0+nr9
ULmzd8DhscqT6QGxpD+8CtbcZRoTHtCiBlnq5aZS9z9aGJlQ5Y5LH2iUgihJpSqm
Ihq07cHT+Lg1juPzRx7tyH5sWZW9nxt9yDlbNGXFwqefukp11jBGI1dR7VOLdamM
VWP/2LlXOdM15QJecpnqwzxQdhuBT8TYDOXCY/WedngYRA2iabHG5ypPY5eomre/
Y63WwTg9X1GuCtao917aHyj99gLzm1H7vXbxyCgdWzAJkq/i1uO6kCMRlnyCw4BJ
cJm6Wl3yQjnCqcf2wsJFdSK7TDcJEo4CGokzk7Nd15ROl3nO2sG2cN7e3aWtEmkU
cUBoZcQwXlo5USQm4aR+gr+Buifm/5ZClWgEvM2rhEi9VVeL+VCjqWcP1KTrhhUl
21qG9xQ2EshaN0fufd1TL9PZQanNPMBmVaqgKhdLrMbEYw/VSYZa0H2/SDvanMSh
QCM87q6WaIO8axLef4xlxJXhVLcENRfJzR+7SwFGnPycxO+LZ1r/v/jNr6Yyj+pr
p2JI0rdSfll2cr0pWUMI9nicC1/+xCvrdm+yhdJnsLMxgRhlrU19yoFh6VGnH35y
SaVXGPj6BOBRhm1/Jjf+4yOuMyy5PkEmMZRx1lN6fim0aJNnXBtwdNqHIyL/cECl
KUUVKof0jH9nM01bOd0oFyk8he7nMX7aclmuF+1jpOitwPRfUQAiUowuk+BnWwTJ
ZK0qhR6aerzlobBO6iVaarGgvtygWliZXiPwp16PYR/zpdk4RD0mAXLTh+eKxq0+
24r3nvykm6E9v5FidvxmrIsa3wlw28Qgr0mawRoPvV7nauXJycAs8uLGKHxVfGaY
n7LyiGfFPZwd6Fqzb1McUO0nSbifdoWo4c4V0R/SRbAmrFW9oQU2prGvof9bPil8
Mj+qOArZjcbJcU+GgvQY+HBBcmRBGfrBHJP2O3S3/lWl79lelrVv2tM/jO9SUUwP
AbO2ryhyuYiEQ+0RzDBR+C7a5P2v3ktJJcuy1vcvLbP8LSnPJe9AsZnEyhtqUHdC
kIVua4QPIOj87D8tWipD6U3x1zQAc8faZPbUR0GYmuwlkKcCgFihF1/cmNYfM8q8
yqZAq+zc+Q8unYbfxSXjzgQoDuQIdeIZI4QvyQdC4vIvlqhaioIBmDMU62W6CuWv
hMT8pmYErwswdLJQyTCJAYF10oFjDtXwm9S2g6tGfs413Nk9EQvgHLAy3QRU3FGs
UJTJjHuJBoAq6hjJi/5ulV16KKZcdBkJru+aSW/sSoKxjCYeXIf2MzwOVQcNKWvh
w1uSrhjhif1azmMSrMlamJ8QsOSmZPFrqx4H8Vlv58zx/t1iho8BQ6NME0MzxR1E
sXBql2dpRyqeiG88ozcT5/y325wcbv01th8cGiwjbgMD/UzGHk7WxwB45ZtLfOWb
cWnT6/DKxK9ZOavvrd14jyfwAno0ND0NQk+MWLmA4E38gIdWkWS9Avw/KH1hOv5X
fC4co0rSI+mg0LHDkBeuy+NdmL/uSpU6cFUlaq3MNlXfgX5W5Gz5PbJmLQq0asy9
9J6wDdW+YVt5DhZ+nq5mHng41PAU22RfcIhx9BEL8ZGSSpGiOUmkeGEULZStRp7O
NqlqXyWjboQVulzQpIUqio64XESKiDScIQLFxgpTFbWMZMKCOmr3pjRTXWbIQjfV
a1mN19kmQFjJGuNvYPn1Na+e7ttVOaCede4eMYh9LUtMm2RHdPkKKC5SsQnIfHwG
iIF/W5SGjnSmiE1MuUU2HkU4FKQlbEO+eaHW7s5AoMqPsIpyKHcDHmmlWkqcUb9l
5cBo4x8hoqkGIqRGGFHZMU/0ooyPSvw3MdHhVtbveDCezIIOPQbC+n+Jskx9uag2
pUx4a3b0fowQd/+NPxffypAQI7WQ5a9MjV9BA1lEJdMjUU6qcEqfgSB6IO8vwnOq
gklbCs5gHrQBeSjuT5yoJBydUi4+gweIDsJ/I3o4pGGk4bKmeFqMxAO9dWY3UCZy
D7NHqTwW6c2e4Zd5WjyP1BeAViAK6cnwqMH4t9XNwPAErGo5R+TGsVGC8Qug0QEm
uBJ+muIKk5ITS7vg8KFZxCEynZRl52c2wrd3u7dgIs3JElslb167ihrSX//rLwOE
QED3o7QvzgJvI5L32t90bPnriIqbUIFcoCh+gIVC9h4torioQhywhIPb+NeG3syK
PN6neAy25hjkIA43Py8CJrvHc1auD4DtovE6q34Br5zyG8AXDSejrdmqQYfkn5/A
f9k1yxunjITZjxVyqziO5cnWkP6OIjCfvAqhWr1IvJcXHLdQrqUby6sONnGzl/WR
BXj7DSuIDNgEjaY2jP3K4Jfy5h1Rrx36UYBj5HQsNWmi2lQQfq6oqV9bIwnzVD/2
Z0F7Kk+3QMQkHGBeAGWuQcxr4T5ZFh5GL4hmtkbCkhj8mw3cGHGRWquk2sOTOTlo
M23VOiqbefE+wg8rFxoSdoq/uCl3fZJAh1393XEqj9Lpufgxuf3705tVlmCvxDp5
00wzXMfTSFb/DO9yF3BcmGrBI8hzt9x3ft5VbidExfnSewkFKHoAYa1elyJHm5jK
3mu8TeoDMetiwl8E2IRoQfQf+nNasNvHWP5OydGCt6qeb21DRqWycm6GBKwEjnYM
i50CVa7MZ0Mtfvb6B4aNukbVlMPriRSq/1tZlGRQG19pDY57wSvzAh4FSqxayYsv
Q+QxdLP9VC403D/AF4d+Y2j7iUfn2LbG401+e38lKjsAtjajS7VpyPxQP5Q0xRkk
JFhK2jerp6V6AQvR6SEy3hgSfiLi2Ili0Iwy6aUtOFsIb+jSpYNFPBn0Kpa9THbQ
qPRx0JKCw60f58EmRZ2irGEXn4Exvc0oMF+RSsYSZyAeObkL7L7g2nbLKflk30st
7SKenSI9W1zkxLN/qcFMWQLFxAcKqpPDBbxfTHdSMGtWsRZRCxFPVpj6lE7Djwvx
+XjLmhV9ixlrSbsRDal0ESRh7tHSVI+cn/b4YKcTfHhI4pCv3hg0P3oYrj+OXhL2
CyskE/owNZ7T8IPPvExIViW/IXiletHOskANSLI6x390vrfYRUDSWzPUnkhHGCd8
buBZP04hWOAeSvCAyyI/drQ7QPSCELyteTqH3YFg1N8+nWc4FpECjlBEzWrzi7qc
0qakpawLQigcY3cCdsaHqEV4Y+joBlmnOeWYofa3mi67iPC0WyTlGabhwYdZsERZ
3bkFg6Q0xj2kLVVM4ezlvJJHYBJdo/FSOZGZmwVcfOJs3Zkt2uG/jlCT+Mb4NhVL
Lc3awDaBhZXP9nqBqOCWB8Wx5jylMU8xK+zyq0RzJbwWDsOoOOy4wz0RgNyqs4r1
j7osbtfqF30rFakKt7HKoPOLJvDuHW/UAQkpekrv0joEQGiYSEsJPnwcNHCuDmVl
m4akWpwUtLw13wXzzXrVpzmA62dCh9zFphac8ymapGtKUHGnjFdExuK9Nsu4YL5+
DvIEtE8wtfabQfZNTBHinQH3l0y9tHnIppaigG51frfIU2MMlwc5PY40vfEpfen8
cyL7VIqEmRu4wIx3zfQos8GDCGDfveq46ngMbgaCRmtmQJQnKT7ewEUdNfZFAEX5
APKwPK5aaUhq7FNjSBykSE2KVBgRMMo0QrbG00numhTFRFOD+NiamjMRBRSEhckF
AzlwICCwQkW2Xx52o42askFdYvO4SizE2RONGoIpSHhyLj/J+DoAmEoln9kgHMfh
GOYEWtB/LQnyOOorgy2HuFY2ZmXhr4aL2jrxCGq9E34cCKGDtGtIX8JhqoUC4072
ZMYnwOYjNfmVuLu/IXZiCosYmSAWfZ/P2TNCCJ5WPVWYM3cZVHLp8UbLKUbjwveE
f5+d8iDOxHqD3dFIB8VD5Dmu5LvlvuErobCSLpQ7HCU=
`protect end_protected