`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79KRMqfN1CY396i18KXVzLP3
AtV8fZkBIM0v525LE4mEt9+6ozD0UU/UcBYn4J96vibR6dhDiKcTn4B5o9kpsOxw
ioeMLGB5V05cY59psY7TKXznLqx+u6EDysfzP0FIRSZOcnGWbBlWUXQZWHkFzjc3
xKicfDuj0E0D5mMhWEaHnQ7QCa9cUJIoJzHNiSpb/pL9Y7U048moSa1wkWbFngG3
DijkalfTVCDmSfG1Yp+PGyH1Wd1cUDyOeSJI+ezKkt1QFKAFaQeZLj73vYUCo2Fu
r7lh7DlsWWF4vxlad2nmIMxz1FOjUR2KmuSYJS9pdEnu0UL/qHLv9a4wMvgX5EAX
ScMuR8109K5UBwncVksLhvGJXcnSRJdD/vQbNjnzBXlHIvOcZcyXbkcuAktrYjOe
XWAvYXWVcAJk3qJfyEVlTe/WIs/lgaIT/qXhBeGB8G6acSl9Ixht4H8ImcRN+dgc
EtyDYu9CXwffULcMDNBbEzzdEcktVHSXcOvdHNKGtd8SXlNvd3/c1ZTYAfcIuMaP
YJUv5TYDVJwcTm2hstpzYy/ZlhEMyuRzKmDc2k+K9t32PRYKkaKMHBwwcE8E8vE2
/n6B3+v3rfeHnzwmk3JFdBxO5NHs7ZziV+ivQkU6MMIzcYDC0QZDIjck1YLF/cmm
1+suhQp1E1ivqWrU8IhqI6lVD7NVd5Vv63erdfIjMtqrs3LQyC40aCbdO/iE9DiE
WvQxjoZsipiyh7IPH1ph37Wb7H0dEzYo/O2pA+TF8z84BZc81HNPFSAig5vmWmeq
vmyg7SdN2Tbdlrxt7Kg3sZJP9tvS8gvIa1BQgz9WXun8/1Xu6yeUc6x/TUrd9o87
yIFu8w8XwGs3Y5HfRsCAgQlSfVmRAJRI1xqooGa87hm9wU4VoUA+uu2L5PbZMO0z
/P8E0eTvS3zT7vqsLAoTnX6C18Zn+glyu93UVaEMhDdaUZycv67U26D5CKX+aeVV
NkGqvQJzVwgOcCNpjeTOAnkd3mv+YGkPFKu0RQscC+ZLFkT0Mqk8HV/mwABb4fQE
gAxjBHZqLI/H/jar0kygGmjZVzduwbsxGpTcYN912pO6lKif31fn838RQSLO25Ne
Dty4gFztIeczU2krWfgBhs55pGE93/rfCZqB+URxbQgop901j70t4Ht2hk7eWAjf
a68oTGQe2ysExs7qIn6B/cKE1WIYTPINo3XPedWoL7jxS1Yuph5UEdQDOALRqNQu
ikpK9ZgfdSc7IqajOgHPb+dH01kClcZ0qrUDvL3SZqKNpDIMg8Hup+c+Xj6ri/U9
+1TwekEO03UvZQdo5+9+8kqDVW7nw45vuLnp2LuS71xXJwF5rY6vc/lhT3HPnZh0
8VzGzDDaJQ5PSekCXLZh3PDSPe5rKCq6OhRKryykduPGwo7c62tpQWNqANYGmy64
+phDUea7q67x+jyqQMu9UfKl+q4TSl+3GSaooGulP+SX2KgTlGXdpnNPDm7lTGaH
ohWCrLz6VELy1L07HiRr4ge1eQSlS12pdxqXDEx2/Da/2kl0DwarBZboes4g3RU+
PF3WoSXRdy8quk6mDFwjeideEWBsrF2ULQ2NX+xH2pwMMIHMBYi09p6GGCLJpRZj
ngX6XgP7iIeNB0kUa1gJMYq4mYX2xbhr0cT2lhaICKuhR3Z4DztVBLFAT7xPF/2D
GpsTAMYkg8N3FZ0FxkqlvrKDqGB24/X0U9MOry9+/VBDimHSczFxRVe0p1SGGo87
vjL1S1sI9LEFXzgCrR5YbEaeqjWbi0UnfR+iK6EBL7jCchdKFJDpYqy2/qsl/q+V
rAsKiYQDX6E+eryNoEtB1z73rCwE0vZ2UKelWyGBXYOozov6ux6Eg9zcd2Ha5WwH
3eXJ7ymVmTudzo5X8QX7uDK7BOom7Q8bQRbnh+wRoBaEXl2RKfAADvPdvpULDEj6
tJz20DcoGb+JXVOEjHhZQENYB0ACBVQMXOAKsoJMomNRvMTqyFhcXIFgt7iOd5aE
2N7ImRoJIIlS4ICcXWT1QGyuPRbraxti+faTKtw0gNeMbBrij7ci9Q0DBQWhHXOF
cGB2bZ9qtBCj4NMwAO0VubIytfosWbkU3fidTqvCTOu2ChAfYgOHerRn6rQSGKwg
j7ybROy64gYRJjDYPCCkcCT4GJH8Cn6vI+KmRkgDrW+D80NeTnFh15EimC8ZnqBE
Pt9tY2j3Z/CsoXSxSDVbYNWDMlheUQj4DaWsDDTw90GI28KME8XzkJQKiF4Uyvqh
/Ejue/ktfdgIURHiU1EXQx72poYdpNxf4MRJ1F/F5gWkaLMcAYgJVNO3w34DP92w
n2Xnfr7gZCgrVTMFEjjDM//ULqcoC4ivMlYkdzGr8ofkMOaBlyHyf2gjWkI9/zAi
d0SVPd+rTun+SMGLkqJGtLlCjSbNPjQvfoLd790NQbnheVWCLjvNh41whn5yNIhN
xUZitJZfCXLoz3xrgIdOxU+bapYjoisO+iPxMpwhFF9Ng3kX58wpZ9biTqOc9HWE
Xo43Hkb523bZ+dLzrEJDhKJpvxvbFJ2Sf/Uu0JL6/ULmIVTcH+xNHXJmLDCzVYDC
8J888OwI8Cyl94BrHS/i2FGCMDBl7CPOw4Xk9apByXIhGXLXLjRMsvDcUC0Pxuy7
h4WS68ixoc5xU0mTtw//kgX+cnj+CwS1qUN5C6mp59diiDc2hAVfat7XoIcNxW5L
Tg3nylVTXv8GMlXZsh3fec53UXWQ2YaVg5gtyIwR8GZKOwH1pp6zuJrCf0KR/NFe
+xSeaktPizF7CCDVE+rg3U2j/aJpoD2Giluf6OztVw62QcatSNwa14g+bnBIMG5m
tz/77/yTBGn64xe24jOB+W1TXcuiMeltxai780hfSf1SNUGJttZjB2wMRqprapRf
cBZ0XSX4oRH7rWwn3MEWHDloIHwO+62EPQUmcIOe1ifMLKmR1knihyBpC9opYC8j
ICtMnfaK90y/Hb26b5+Ghpu6W5O3X+5SWFKlFmB0WJIOlzca3rNxTRrq6aEoPNDv
l/xwxipctmQ7J00AsC+MVW5/6F3VjD9bULr0UvLDAoOCqwE9ucB0aIM36KU+oFPr
1Cei0v9f1KdWxQELkHdhbdHr3d/W0TJLk7+s9EonKs73Z0TZ88ZgRsjZfFHVCKoC
JC4ZAyyzqhh2cdmn5Q+Np9eZL1jIg51BzS3k8Sx/ahWjB7K+OHuFtMH66Ngg8X2s
/oMWnpyeX8IFsN9ndceyiFVTTyeh+wmVYJDGpc8zz93bV5TQ9NGYAAneARWvqw/+
Ng+BC2Bohx6X6EvcYarwunTQ7CaAWxQBzpjY5ud7F3WmJN03YU0h1WyDqAtets/Z
e8GjmwmRTW5fI0eEGGkwdrBtJws3HxlwAni0g4zP+ThCxPYXpYJWthZoVMHCrJVk
TBM04kiKUk/zSQpr+u8pGKEPPD08Pt5qYKXKMeoA6DBGyr2cRRsfvH3Tvx+/U6H4
2NGiI5Kp54iAJzGUaqdw4aeuKGeGz/r8rMZcI/faI8+lBJAPW7j2Iijg/A1lp7dg
IILyrpm9/si0aqJvGLMjoDlVIJ6DUY90uOpPaM6dkvSbmPMc/4RYie9x3aLC1zYu
9DIwBSTsXwJTquG8XDkM9NX9R/DawOgJtN/tB7GfawcBiklbIAi9Nh+Isl1wjejp
jYGRKg+CZKnLNKigZBmMojs7LIOdD1xPYHh7q+zf1u7Gr9tl9eikXw6A5AeSq23e
NtUsEtQsLV/zR1S4MZrH/LJOh7ny3tLIcJyxTZnEJCopnqOGRgQ2oAjrGJBa/VA+
KlsEIPwvgIeP12CO1WreEUQQ/5sM+TKLdqwgDYMuUfJL8B/mLBcGIAr1ATA+YYsR
1ZF78QWDPPsKNETxFnYdqx3C1v+fcAfAPWF1JM9ViJ2QTWDAYR/Nu2T3ZTDf3PFk
2mYKnN8RxZVgcymHaFm9Qmeul+rkhX1tdCA6vBD1XF8FHNtFyROKXFnD4zKB048N
wpz6Lcpf0pz5xhMYeupr2GLBIbtoRAJArFwtLa7GDuA9t6KsoNO4hzpbUQZehFjX
yhnP0hwLZioixq5ntREJRAL1DhZb1aMVP6A9im/i1Jp69ODhcrADL0FVPISug7QJ
zuXwzldp2pcIf2drnaQUwpXwsiWLKXDI7eMCXQ4LqP3tOeE77KYqk0FHMxD7iMhm
2pHuohvfsXv67PKcPrqeC3kNSSgFh093kVPqlcni20JzHBXv012oBKVGHiy2/5Xh
unJ6JVabrqWudmzmBmIhmWvo5ilqz1+NLiUgbizj/6muRqDFmPQTv/3eKP8Vh52f
B/g57l6WAvpDsLUgU2MXq0lDsRFl/O3y2ubEXX/qzsw3og5VrxL3IGzBQ/Lol3z9
XwjdvHVQTgZMWRMsD2AkdSmKeDBvlSE235mLR/1nde/RGqBGyB0HW0lysNyjIdD5
QhByEA3PyIc4u6dL1GOLcKE9Sf19w0gv2Xz3Wrn2kvGtxoQMs5dyaGC17UyHBR+t
tTCSKpqP3+dJxdoO7xPCbaUvU5oPi32/5XwYlA7XhjcAHUSPnVrvLtA6+sQVZijg
YccrX8xgGWdOXSzEE7ltXtmNWiCiJsWcOICBJ0p3RPaxpSw2klY10uOYoPBUOOo/
bTbgTZooPnVTBohlo+0mwI16CghY5U9g7eiq5QlP+f9W9IoIeEP096tdMlvAK1G+
uO96PjD2T6cx86uuIRv0BZozN8Y/zg2DKDzrInvpEZ1KHPJVE1UEvmf9YdmabqxR
Jc9Kfz+HJ0iWlPCxqmYh84KF5TGoDJrY97hfuNQ5RmBjiCMViWovpd2rSOjPv4+T
ncm79gcHX9CqTuViCrQbzKmYW4dSVfrvvL8jLMV79VPBipfzY1bn4sIphmDlt8Tu
NQjjfv+QRUDpU5nSAiPTJlEx5/sLaDn8zvnE29+yFaTXbg1Hg7edYyV2xVpJlXHH
l5N+rN1MZ89gcsWHpSjrpizZCtBR8gub/CxwaI2rxTkApT2Hdej/jVK3L3bUtBK2
FFW/N+zH7f/I4ZZKJrT61ZoclbxmVxBxmtsMoSq53hgntY7BF7W1UhaSsmQ1oyEV
TssvZmYxzxYEfy3F1AvgyAqSKsIQpCmEQVDHPqN65onZdKTbQlkcgGqxwRvUhhGD
rxBKb1rT2aQZjbp65sLYelhCTUUKdGne73TdB5lz7jRlrC41QUuv7W133MuRvY+U
7u8R2+B9tnaIh38MmwD/NItRRkTIo0nJ/n+ehDtoZ6Tqq9GVPhfjmp/AOoyatoer
Q+DF0Zl7nUzhlV0sw6PUXgpCMRbxHpwAHRtUozSoxvPiEW6zql7f2r45RnTGBfhL
WmrT4DuKzozyafky5LifeF+VyXpnfzZbRDAbSLuYZyFmaiHVP0tnBNqoSB8vWgMs
Wwhd9fIBnWGBiZpIt20h7Skvra53Psi4qgdKfAAPSnN3im8QRLVwQZUJox8PVnlE
hdPhB6HE7dJLLljYCwMNwWbq2RlLUTtVq0rANuYtzDzdmPIAVYX5KhvmoOPv9yVC
MljWqe9a+7qKfjddMIEu07UMakbcW+qUqs6IPEb3oMh7Id5QEHpwVHYw0hxxjaAc
MWJ/zFTjcHihfmfLWF1VFe5xzsWvUYIbUxR/tMRJQjnJ0YtKrImDKUQxJz48WLKg
XNwloSYJxk1CDVl4pKTyQqSbG6sEwolax5qw3yMAnQCD/SvqVRy1ayCEGoOrH9+K
LesoDWvn2fwoSH03kjMqScRe0i+VWF2rpo56DIFGT9bSEAfZyhavNAlrdrYsz6is
qvByCn3wKYb8fZZQ0tplWisCwildrh4dvIP2+DiTXNII/i/w7uuJ5lDaWcf+igLk
DSqq6sOqIT9rJnMYfVJObkBr1c6LAxzod5SgcruL5MIamKX/YU7URG4tP082p5R1
vOelHjwDvU1OOWz5Jp95AK9cWx1ZR5fwTah1jrbhfsPYHPeWlma8xigp2IEHRwrA
kBI+8bixxm+V+AQ0JauZGnKbH2vH5+6ZNESX4zOSVJg1xqLX5wL8TGvTXgR8D1QQ
FXy8sBOEuWGtjGvaEpSVG3rNPQuyrtd5BTkk3s6jCGCVD1MX4egirJkVb+aUTbDq
MlPIebmvywFgKC0ZSu31SQWyrKlvP0ogezLTaMK9DIXkWuIXyNhn99jtWD7uSkmy
aOWM82eq5DRWWm59i3AOtgNZ6TumGq3h0nUwzSoJQz9q75vbYJj5uo9nyuTkZqDw
vLoaWmUI27CEtvEEaP4TSN1mh2wXTAj+5viYTgtVMrCclstf65wK2Jjh2IOY7Ru/
vR0OHYyxkCy0XosJwopduRUxvJG9AxFTwr++1wSGB8V55tsNfcTiUjPH2QIzLb32
soyQqkzs/YSPzVFLQC1M2SScjAsf5uszemVvPXsGVIheEPPw6IUsNewsvXvnKUeQ
1A1Icqbs6qucjHPJSfyGi1Hb8wAjL0WL+nnA9wp08w7RYeCDw7xh9Lf8lqbINoVz
oLhaXAjGaQBGp4Hsw/5mxJsS/tzk2Hk5epV3T/hlY0TontQFoNeTDZxZWmDNz0RU
Fma1ClOi8GZ/Wl/ZuD5kcyj/XQLfV5cdo2blV3Tba4at5r2LgrQ8YSV/bTCJUmyx
ooo1YyTqzVbW+//wkBQjdUi3KHpDmt0dlsjGDMvdEJuTq1B/AtJE098rkNqLr0ZE
j6qB6j5t0ngsvt7OgT8a+MUIv+nXZmx8lkv9WCuB4ZaNf4xCH3yUBOd4OhIn1TGg
PdLtz6jhtOa9FoVdWYRkF8xK1N0df2Jk/DfmaU1zZq3H2cfY/wLQ4rIkkoJIPpyM
POq0xYNcAjOnRBJajjXKOCAX2IRmWfX8A5W1UUJ5czDdEFv2oZSi+bf/dDswa5ym
llidrx/1w2c58i60xE7H5NHmt1r8ll9LibmcAMzgRpqkmTOuPcJlPyDttAZfZzv9
Vg8RLW6oLgzZPZTAvRkbdNhH56ThjdUl09ZEMGvqLqLZ4DY7y61Y0gB3pWoSRl7D
IxynnXLWw8RWStv2VZL+02CxcJj4tpeeZhwRgaOrKGONTGRQRmeDocj7G7vDsB59
dgHAVztVrXx24UHffG7w+BOiKat/5HBrUw81rkQoVwKO+/4D7rfgJ01m2R1iyBJO
immwkIM7rA3CYhtiE3AZAhYHBZNueONwWLXvFQtDLCt/9QMpV12gdToR9gydfln3
vzC/sW3OAgsBicOcGi4SfvCSvt/n+V+/hAezDoraqUf2hSnFtlHhf5K8eImOSzaI
GKcnBBJw2wJNsZvMwV9D/8D4Nx0hzp0r4lZzCJ38r1FOJm0M8a9RVqSQa5rx5eeV
EhzBTR82MLZBbGCNAzbRC9kxi4haP53UEgbJyjBUqsXk7zYqLH1uO6QGtaxkNa4V
OfuPYud6v7GgrCbRBEjTjM7rwCSC96idxeG7zjFo/cPYsIChs6blnGDjgDooGRpS
qmhypSJBChr/xQnhp7c6pqaXeyh4fXeLuieRZuxzkBY6nTe8mc2kBs84aDPil5Wy
fVg3eRx2HyxjEX6h1cPbfsHFOXFEekgVgjAqhWS4zHEvDQFUdf01EBQ2GkqsFcdw
agtU8OpdkI4+iVxvy0YN/18llLqz01mg248UbNpFFnTA19v5YhTpJ8OvS7O2WoZ6
lOz9EtljL4OAWh/XBv4gKGsK+u0lKIowhw5jy5DcEgSqKMg68M3JtnnlW8NUPmCP
S1TfSdVhNB8V+pdd/ElFvqozyaU/XZjhiSv3uB+2bMPMXwSOaRtM+vjplRMCXFCA
S1+soPlUHyilViCMW1cYzWOPjLVIWA8wn+2fc0NKVIIZv9Jx2JGJ5rsIAoS+HGQH
NHwjdU/WdKXJksZ+/AY/3fBqrfio9Iim5Jzd8X0AJ08kMyQ19N4aNJ3oxt1MLCRJ
vV2/ho2VqBVCYxRqQ7raGq3FksNtYScwRPA413rC2HHA7M50CmTGwcsxf8pj9j5w
NGoD1XbvXVTt8MN3G5NaZDkeFOk2NCrbddBsNoEM50IBOUCIntqp21yx5bh/ppk8
cx+zhnYRfuVkcP9UZaGMGdHhOnV7DjpV/YFT+86ZUyt+exgpaG6vsnkz04XB4aFI
YmirQBITozzhl8HkDcJCztCQL26AbBerMxa9csw9b1lwDFvS1Z2E5lPGt2iiJ4s3
5VxB1mx0RzA4mjV4BAJMVHx0LOWR+0o6RD8evj9AvMBLYwC7Vo59MzbAIDTGH3Pc
exXqAefCTX0YtVDI8GpOyHBf0A4VvXVXQEunzX3W+1uVCyQHnDYLXwIVIs1kn0mX
NxweUq400Ntt40Sj6VLnOWGPrbb3LkLs6H9a5b78r2ZIYz8lc4G1xqi68Z8FHy9j
wwOVYPIqly/PR6mabhVUVdTDrWB+XPG4tqDLs0sxiNjh9RQPoasdKtJq+6BP7Pk2
o3grz7DqA6z4t7NNMlmln7SlDwAgCNXx2p5I8SrIYoyEgg3Cwg8BxuWR+F7QFUjQ
XSy4s5UxzMmTYSkxprVy4hjqWIluQQ7u2ROxvg6RD3YXAvSs4ni5Sm5mrDLhBEx8
87aS+TeGiwSq3bAHiOMyWfNgRFfx+Z3Wp9vs1ljKUogNWUGoaUullbCzNsCgKNBl
iN7T7sl43yA+gIqzsMPWC0lyWggIfl13yadqOTTzSdCV4S4MisVt0C5xgURhDYkd
vH0iM0SJCNtBUFViR8YIcML89HeKUKQ8YFPWGgH/OiLqlmpLCLebp72CRgfiVZi9
9hb3FkJY8h7JByktfunfBRaaWaHcAgXy5PFhHj1BnXTF1hmpxN0khg7z+pP+QyFq
feOtNceQW7tpLLZwP5qV1/2enJ4OSRPBx2FOaTapvKmobmYoDIBhH47EZXooWH/C
tRfcconmzzDKyawfjN8HCxleRD+CReGkP9qt3jslJ+FIbCxnpvSM9sPYUZJPfLmV
C1DoDpLMBmqDTe/SJrowKJCkJRlR/dobZ/jmdV2UPvzOrmBaifxCcZC5TnistzlB
gGi679hcA9oO2tOoTBk134qtV3jlg4AqyqFvwnwioddrUSFohEgVzVJ7DW94/3n8
zRo06V2bHemMKRcRgk05tPSufExBDv1+0cxn7e7HKQES7mWswRqz7zag9FkRK3sb
2jUerTGKWyWM8gGWU9+WERnIBJ7zsnBtbYbI6kmj8m+eJSsNoYYz+P4UQ/dWncnv
vYHE8b+Nny+kDqAaOyzxR+iacVaAKp8yMhNilCU+xZO8gAO5JJjynjHPAua0r1Vz
I1rBROgd1HWWbQVDihxXh635Fwetw+ok8ggaX7n9BAP+UyVLym6/Z2cRm3Y/hXH4
183Ut0MLElxB6Oq54FKgX9PjK6YbzZzIuhgRgKBt09COfzH/e4EaBbffX7Wc0YEz
qJU+XqvOn1+hAZGsMyOK2jIO1jVr5NrFlPw8r1Iap3FMsYj0YU+Ksj4bfKW4vHJ6
hZlO2zYnZYZe6zsN8liMI1bFO2Zj9AfY5sk8phRaRt8KGil5dR5xHTbvpovEi+M4
g/6VRYT4MRswbsAFDRVChzRi6JrbuGJjZGaIWsbejM1zn8CypaYA65hoLTJjncmq
zAC8cUxf1iAT9yTkZktVF+6vaQLiAIcd2Xmd+pK0WzEPByynu/QVIcfci47/h0Fc
Js3sEcKn0TlYSL4fJ3uOPlbuy1it0+i48BurLrDDlqOJH7CJOkAai3yhXxr6YTKv
hIpZ/iCesnZYrjkW3YlMKkqPDkSBOgXfGq50IlUa0w9wG3jrlnr2USEzjTWVQFVW
8rZYRvNOTJnlCxSTPWKq/8uh2Q6SElkWJEAi5YhMvZrOxiHHpYvXQGbWpJblD4RH
duwVwYnuq0hrwCaeZYQNCR+BVKYxq0ZDuBWsB+Mi6i07TCfC3NMSP2yr31mtnZxj
bURrgWQEDVKNi2Q+re9Ixy4g5i0J5/ARJWsvH6S0uUzaC0wHuFTzIsr6GXc8ku9K
h1xA8UwZ+eDIUDV7oRYWVYh4RQimHrvKT0iCqqgAQgTuSxisA3o2v7JSW0y9u0L9
rzVGE3mBCFlsPdgBjBSZzLoaVeQyQrMFmUgs6DWJVzI4/QQkyMZn0055BA88Nz1d
E8OyHl+QeuVdq7HK5DaxNwhgy8dYAuP50dOuJHF7fQ8B6yR7JLh40mH7a2wGo5LZ
H7XD+aZfmsBFJG4iLSL3XU59BXmqvHXqBMJZK8nZ5J798h23ZqQqy5aK1MMImCZc
BWoAHFWuou8/O0NrB6nBtmH5jLMF1kDls90odTfVpUFi3F3mynLj958Mru96+4l3
NE8w7Br4a3NJkYn3+FwroXE2MIEaNiOHr1Y9eMV2YZ4ICcgd1v57e1vXXjfTa6tF
UEAhHO/DnRgXggx1Fp15NMB4AgZE0+G2TuWQe0XBBVNiWh0lT906YATM4CxM+4/H
FWoLQjvSzUPT9A8NFd1JdI+9haTgAnwdHucWKN/o+IMnTQmlErt2qwT35Lb3THat
w5l3YoZse86Z6h+93A+wgllcdr4Fzhec6XpgQOIf9+lDS3FQjal47AgSAZWdakH4
lJrtZeeNthoihgp05CCxGlK0kLTW7V/E3K+5bLDd5V2gzdbKeBnqpRxDumiRf/bX
A31AykxdvUrUZPcHLTnw8Q82sXvaEg+nAw+vYMn4/mL+ega95CeJe+7TpF0lb8ds
0TjdxR89p1ep1Rh/FsqmdOab9R28jHZAjKALGn2CiQb66S5NumvhEJXil47RoK3Q
m8JCdmjKVF0u3tGh6Jkle+lWil9N+5fHlsQf+se+RhzmQ6OkXiwmZcVsS7spS8+R
26xEAw19Ve5w5P/EvuW23DDDpzQqx8sWaBzwAj1tHCo94xAp9KMLbtsPBjgpV4Lw
7FyhLqdTJYxbrRBsNZaSNKixzTLUAsioGuXBGwvUz301m2QrSDsyrjwBnjCDkPS8
GgPn2M3wnv1SmfDe3LG0eiBIal9Tb68OZwAWBcXqH8S73Gy3SC2/7v8vlGVhcWWx
HWXeu2kedsQIjhzzdSkq+U58nAsrv6CwH7daQoE3Wilore+tKijnpmerq181wexb
vpB6IF/AJiLtSsEVuxGlEomqW/HdJ4J5BIjCsV65hw9zQo1qmieqPZtJOF6vqj4f
CRkAMCZG205jWatiYSCu+H4ojbLQ0Jym0GHGKqbOohk475bdBLBdrmzoIj7vLZTh
uDB4hhuPh027fi2BrpZcg9EyfY03Es6Wh2qEbYLgkTabJnaJnmrgnNK2GkgO6NR2
Lb7PyTzAyxVMnSyFj45/1oOBlHDJMFsdnxIdP/bmCd7IFuqwkNnEgnIsTVUXlYf0
rHtRJNRJN9ugludocmmgwUtuqjGajFkoDKR3m677wq6c1Q4wTPtRQ4htjXH8Kx6y
MpqRairpS9R9rksMGDjxjl4bKbbD41rzzCx4hxGghH7fuEafsv0c7IlGHqDIQGbP
4NVXHuPk/FtjZsgcAWzRmlO9dLOwMe9IK4kl4zf/R7kjYmvloZIFGmahN+cToi/V
1VXGupVqRti2+g+S3Goioq8BEpXJiQfSLJmNCoh/W1GRdvhgHWsVu6+HZPvYiSCC
RhbD6TYSwsYtKpVKO+Cwvi7QW0gt43BVebKUkfuaQQUdNNYZX/wX0PMiU7Remb4n
O+Aqng1fzfMTrMiyMEEpuEv7QOYrUeztZRFSLYAgR47k9dHGdyGTlJ57tOysqUBF
jQjMpiUqLOtbHwD8ysDRa2n27iX2QjT3JahUyBlYceKwyzH28URfDJAaDbNgaME/
ZJixYfd28/hveCjeT2baUuH20kwDwTH0g7bWqZ0B3Vr4xjEKPiF+HLnXzPVlKuCA
TAaTZ/VywAOgj/V8aUzVDdjyMwWapiq1T1VIAz3HV3c8i9vYLjTi7byR0ewHSbRk
W3Rx70SqK1+lTAlHmOnfcFEDJ1Oj5HkIYa+8mMuwfi6vjQzkcDh8jef+MZdR2pti
VE5iFaAYZP/LDEOcKjH8dBuVmG9TCyLlvRRacobSY3140rlosaHoLU52OvJNFJfI
aDFQ2PXH8G75ckwd+L4obutdDh2DGW8F6guXFgmO4ZgdX2ejbuFD7Y64IU0Ux/tG
qWtbVXfMOjAL2Swh4hOVzplHxaDJz/+5GyoTbSTyFm4XQAtyvGgAZJtwRT0n41W5
BwfSq0mpw78BWUkPKqi7kTuVi2N9g2dlErYMW/1mHOcPWqi+LEYIkpzaVqyiX22B
CEE+xmw4DcpQhOZ663Xa4WLD2jO2KILwgc7JAnhqhK4jOsvwo/XTIYVBW68fmGXo
IxTO369Et7IyguY4K1IgwC+NYO/BZcg7yw7md8I2e+kC6blq4dpOCqJpTuQmG1Ad
DJYkaDS6zx12NMngWzPLI07x9tXL7LEQXvAqfZqzIqVk8FAAnz+5MDN9eQAHhIoS
QriJbQ/yYuWSteD2Vc6WZbtSvN+zHZbxbbaWjeJ+yadDUcX+TNgpn89vCWxpAN+5
DrB9PtVNxwVmhkswM7BA7mGUv9GgjtFTIvPBmKnk6vBxx+coAWD3z0ETmDpLLNP8
aFjdWXz1oj4hgkz5DIQwfcga/ol+9faRTTcHtRps8nDprK8cHd1/UcVjwfOe1Kss
XwqQ9ibIfOOJyCwaofpSv+ny7NTh0z+S7egi+9jk9dV4zKFo9AGLJGMoQu1GxKLH
mMEXNnfbjAgC3ytfDBy6M0Y9kKk57Qk8wR80n/rZe5sHVDnNToNEvhr2UiaYFcjh
tiMLxfmjMvBH2eE9urgWCr3Wq5mOraW8LoJMhWFLd4PciGEHW3m8n52izIWryPYw
TqQ3oX7SSQ+o47lPq8RWjhC4iYovgeS5MDOYu9pqR/9SD2AXqwjb5Bz0sWxdIVD+
N4pgp0Vanya06UhCGXCneE1uwVi/wzeh+j44B86qT+Pr9h9B5Qs+Xn2YcVRLRehH
83/3cz+cL1TXu9mIldVsTNaxIKzDQit66byohsk36fqEeCdeXXsao8X0RoJdtXmJ
Jev6T3I0q0HGmsP1CC9jT7enlS9P8bJvf989Nlz+FG+aHho1VD0fGgUw0qsAM36Z
+QlkByWMcotLSGB2oeAHtkmd4pF65uO0c+OwZMfYcVo85hDZTTHwrUC4DhJYDkbt
Ie/g8d16aOAPkND2C+UqBqVGgCOIZLzF2CKQ56j55fIAF/CJDvYjnHeCNtASn9Rx
Eq/0yc7ZbVOfIK8LNtNE2+jrFO/tmUKJzxU04AxyMKjk29ZS+g0wNWT5VB70irVQ
VPvf4HaPcNMkAUSR+KvVFVAUNtHtoerlKh32ePaIXP+yVgfhTIGLzNjluKjDD2HO
dihvPSo6+lGvNsY0YinNs1i7WGN/Xgkf90dJ+Cf7qicyfaoXUMBATAgRt13AmA5b
5ogkmUbblbgR5Vc+tURUPBvbpcfJ9NWKEoD9x3kDyq2pO9YBHzooqf3wmnylCIik
fQ8G4gvx//AZl6Nhs4LxZS88YB5IpgMvfYNA180Ru6mfJG61mkqwtMY3l+nobtnb
FApL7zvew/3RvBBlJNhAihjmFoGb/shm7xsRke/VpDiqo0l3BcqfK3CXCQEoen5V
wtSAdIGcyUgC+QYcliBMGGFBY2k8EoL/AMGq6cxkBMrnnDLmxvAwPjgckZfaHaSV
uLyVhKu3mHkug13wdCPltRsqokNuXapi3/wkys/0sHU0h2F21HjZd4hsTzjPrDfM
2o6ij0X7XP/QyjszQyTpVRvmLNvaQBVbDboshqzkP+iVKNpegDRMssuSgbuEap2e
KIz8WAZcreiTgtBhlNKr6HjqefrbW2hD1PVI3WpsQufU2JpvR8dt6mB9OsTcA83v
V2jHCGU2ivw0yXJ2OK9mbhBKAN6807AjDneZrBmHBkFLerlKxlj/1q9z77MAJ0Uy
pIYNgtGO0VniNb3qx03mIvoBwpapGN94/khVX7YxFem1JTU0uxczif5QWFQVsAox
Kro5FmXOCl7DuqgWtPXG1aaaxb8r6XVpdBA4Dr4cc7omheeuXjzOPk0IjmrILkxt
5gIWQBkbEyKo27ePh0bL3tgjBzbmkZ8y3N6Nmammo1KHgAw304Kx9FNsKaXg1fKR
/4DLocerKOX2Nxrmz3CUa3YTFj6wB3kPxfJCwwthGgY5oXyZgsWcdfWocntzyHZM
xOLOIeNz1U9TS+FJM2J/FJsIClylUhP80cGqGpn5Ji9aPZQsoHTswM37CrpRLtFs
Qpu65b9cxm8AWH+BGG9izdYpWXg7EVwA20HgbRe6/B5fDDOl77oxs8P8MvxB6Y5x
iUlniXef1DMy8c1/pKd8NlPciOvQHbDuIqcGWgsGCYAPgUNgI+l/dj54NgKcEleG
d43w3MiUBu1Q0WpvwP1kgHc40bHKBfo3uRYW+9HnIxSsRiFFTyzWU8LNuOwu3e2R
Nfo7nY0KEi3QWqhyO8kOeujQr5MkYXdDJW5kNo/ZdzTerV4Rx8f7cfiiw2exUsPm
baUgyoiZ0nA6QSC5f+5Pj/02AyU3OylDWzOQGxCHTrMmBiNNUUSPixrXa9DeUoJA
eUBGn80KzTctzvDdePWoxVm/lCFILDUoQ4puXSBteW1e86NWA/gJeiuCKV2XvSnT
FaeJGum1NXhk2+izZFot7jMYwT5bRr4fzLV+XacXEXelQIFZbpPRpi38D0Ha8yTB
C23vdoDkiKXCxis9QdYsRM2t533nSy8eLEbBhN91tZ+wgeWgza3H9ZS6YfZdIheX
2wvN5p6D1I4voU5Vku4ukiS9x4bFesBwPUBkc5q/fzljSAPpYrhQE5vBIFmXiGql
eMQxNdwecKNhnV1jl34AJDEeFFN8wEkVBTnOSkCMmXcKErzDOncSZ4V7yPGRxAMO
42wVeoCp9v2u7bGanXgJXC3pfbd4YjR4F+VTzJpTXw3g0K0eunu2jTp+sD4rCiVX
kB5d8z5shOmQyxCQjvu+WIwRD2voBmbQUzrdwwU75PDqLKoJHjJ0j7VMJq3KqwCZ
pFmqMK7F9jMcSy8DaarJXDVjWx1VbankdeK7V3T9qobvcbDffz4rhhqg78Bvuafn
sCfUyaMi99Kyr+Vha/y9a+INZKJ6nW2FxqLEzpC7o0y7v1ONCRtNOG7RnhZjwZeB
YK1gVhjkkhMlmE5qVgJ+s0JGlrMoo3tYNfbguccNKvH4nZMV8RLFYI5ULWjutX0w
rHvBLzLh3wmO8Rfm9U6PbXNQQ6GvEp6dKv6k5gnlbIfb1IjyA+lHyZKRWQciZiJb
Tso3SyQu3ZUb6osDvKq0JhloRR/6JXjkr/DF1uN1RJmVYuZZSZZOWa3m2uZUjcba
+r476guQQzmb/aNY1RHtqSZ8a22TzSOte6vNnGHsoMXUolQ0YoCQQbT8/q0jKTla
8oQAHID5wQCEBwJBi5TQCfFUphOSv2cuXqfmzn88NsQHikV8V/pgCUZGqD6ZCxjp
n4T3U/eEC/P/ieKQO0KnnAFUD3oavBoD8YieX+Ae+5+p1f5zlFojIY4i76oZcluK
kn0dKFcXzkN6RNVjNngaZFo/ErJ/6QHPT7/8TjmQLUSAVvWdWx/muMQavoF95Jlw
a+O+69dhfJHRt5VvXTZksYcIcn5paEqMxkeL8aNEm3iJT2zFxR8u9+oTy9Lw391d
NjcEkfqgt8eymSkkg5uSNSn1Kcy2uO3EUlUGg08xD3Pgf7ryQpZZxUYOlYcnCgop
3jAG6+lEfaGcyofLBEvAovP8HDw2t3LhAcZCTyI6WJCivXNU8czKslToRXHfmCCZ
MQ58jcsHgSvE1eK/bt/IPJcKsB+J8/vwV+iIhjIDg5uH2Aq0QEEpKfG7IpuC9nA3
gMooW6dffExa6gHxrGqYxcgQsR3mml1cWM2AVOq6cCO1UxjT90lwmVzifwDpP2ww
2+tVT4SulxLAfHSv59cGcLWDH4LeGaYjKUPq7TLVfIw/KHoYUXzAWDnX8a7dwuLa
QDsA0wmbRswFm8uQ6tLHdqp1YsrOydXeekcabrPNAVLr82zS6uHg/PlWvexYHJD8
DcFvgZwG50o+bZRVMLMp5hJu6sg63rOcKPZJTZOU8vQ4rMfPLffKIfR6mk5LrYoG
Dbgtt6bEwMzAQVuc6jBKLA==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aYEGshOCBNLOAFPz/YVL0JC7/e3ORytFJCo0DgZmCMCJ
ka/OQenECggJlHxdfJ0Tq+iWvsSDG28J1fT10cR6nuFFrhjW9bnWqnMqjJToWbY0
wWs+o5WcOSvlR/gGqM9eZblFol+yrTsy217ZIhFBJQ6U7c4XCX2E8YW0/cGSWkhH
OmNPmvA2xbDoqFiPj937hmYUiqPe95LPcbzfC7T2FA40cVELDghdXYF1PMrVjIQI
bkaTvMdJztDvqRdfhFeO11Q0vgY+I3RneQwKN3u3bidFQgL4h5vSfG7g/P9EHDCa
0DcVWytVIwi8RPPj7j5VxM28gc5bUOqmho8TBLn4am9RLqYhoFK+SEkLt1d+FYLI
QfekQYGRVh7OjzrhxDE6Eyx+UQLVITzmBYxPyahnDyZUT/W6mfDawqDEF+uHS4QX
UmUWYVkTDl6JefYn3hdsZ7qLgbt1uVtpQl+vfRX5QzufvL7frNgeoRWet0sq8ASl
ed6x2LYpaCdqEO7H3usSLOe+Xed8G/M8XrX3Tmm+EucvMymG4NyQKqROZb1/CBb1
4ZormsFRs/RWDknAbbWwx4btLWLD2iPCL4d0BdCaEvk8JPP++Lq7DeNO1+mV1m4M
E5NmaPnsRLMp42jOnYu0fd7dAeK7EqOPlBXOh4+CL9ATHOTXjaPjjiw5JxZhCk7x
yrNBRSFh5p+0X6YVZglLDM0z+1G2fK9eiodOiQ+JpNn4lPWKgZFyV1dsUaO4tF5Q
aXUH734MDPhi+gRfPmqYDO58p/ylEQYQ3sgqrcB4U2MTR3u/E12Gsgo2yvoDXcke
6LMKyDYQ3NJSD5YU5FqaHxBf4sZaAgH0ijuh9r9lJKsSoG2znfPRB3rfYLDc1L/l
HokYaxj57MhRrK8+Yv+SDhBkz4Dnwh7YArehwaY+6iTF90Papnb3BHRyncmc5aDB
DWkBbL9J/U/j7HlhXoYx8kFYNvXa/fX3DzlI27kivZg9m8qQq6r5Iz4LGWk8Xk4Z
O96+FOA8GeIXt2L8CLFpCF7+8LoUCWlxwbvR84TM4GEFgKG9kH41/ivLGxJpRDKD
L+oNUk9hpqJ+kYYEV/byON2xKkc/WQ637Q8bWQQ0ZfM1Fs1DKkKBRKw89SYc5i3Y
Alxvvljjn9hqoevoD3TErB0FMyvON4aykoYtSRYhk7+S1IItR72JcbRhXDOPBh8a
ZKad+UZmyoU3AUMJI5eP/etoyoea0+82WFWudKgYJaP+0a6n/54i3rD1Dh7IJkIE
4lBxZ4vDslmEVS/yggVlcYJuMS7+WJX6nb8WJeyiJ3abFHKlTcznIfYHEgdX1xrQ
KOJbGl2jiyoETinYX/tNCWwBTEizQWphp1WgfSgTWut/DISKYJPM1LLPn7xViEdr
0y59j8Za2/45M/NzBwbhCPWA+YxoWsGa1bjYvn49Foily6m7bNj+Ao0n5b4Fpt3m
harHLsNzCsDHcMZG5ZWuJo5+IkL8KP3+8nHhLZ8ucM4ekomOGA/xTN63H6fIro9E
sJ9zr6GLboSuwvQftwhQHSfoKpm945M0swH9k1pKhioSHFIrPJMOZVuLUmGneuII
pQ6n9VtvukMjNweGx02R30u6Jv1AyNgqD1OEKbp3r1sqja8lsKrr9qlG0/hkYCU7
+c7PSRzUiFyRo40AqDI3C0dMW4o9rNVBBBqVUcoeFVgx8e8BZrTBr7YPnXOgGHoD
zShpEXOQRdjE6iEZqyrD2pVN41fbkzWA7UlHBm2FxdxA/45aVpD+lDP4eTn0hRmm
0XdhSCz9dIjTJc6V2N3uEn3d1xVPoQaSYbY08gO7cmhh9Knu6cSDrKZpRFgwgk42
d55sO8SG4kDFfxpLyV+w9jzbIvSNryFfBnP/R45+P+m9Hu0MhQ4XWe0jnVLg4V0j
r42pdKmdDx07QI3yt8HhEqjehG9NbbKEh+b6+o4lrzfnXoVe6XOQy46cLQUkp/4a
zOJp5+v9Xj5EjfGdX5ea6/ydZYOk0x2gOv8DfkAzi0fl+lZkxG8cvEWxN7d83GR6
70eQ3rLJPtZol1G37V6Ivy99ipT5GVuGyR/WyOCs3ad740ZAaVw0GV1HK2po+ZdB
7pvtmoWTGRkIU7JXgIO0e1cDRZcZUjsjMDNJmbGWyHpklaSg/q+QdjmdhDygHry+
p3Yb1GZXtpV2PopazAO1We2oxJ1Gvc5SO6Zxo66TcXggjCS49eli7DE5KjBlFVsl
SBIcoQ3egIqRVxCJofyGNibRTab51mOC8311yk6nOxO+GvALUOWsJ7hbgQ+LVK+W
CQ7Qh+5S1X38iyQG4mafuWvMGweqveSXMr72XsiJ5EjdOOTWxICDVJ/rb/zvjMNW
xr0p6NEzKmMaTtl7qWrN7+lPTgAezwP6kR4yk3vpvKCvxagptdte2gnLVmqOy0fx
HUqRAujciitLyXANdgyDoHKvqGnoyr3lUFbidzbYWrA1UoXqo9T9L4oJ/7sv+xf2
icUSe669mpw1hXmcDOGhOyPs/PIhy3BudXeMuhiNx6XHUs29wGpmAz5ySOLmGgW+
WJd11rhTOxw70KqF2CQTp3Jf6+jQte+6jnQOG3VATRsj4PvG+zXYJNfsMgUpUBzf
HLNfAc1j33fZS3gxFmU4xrs1zpkhV2I6alux6Bn6KjlyvfIyJpRHhc3MkvHT8Lpn
lCLnrSAgKd55V7fDhRpbzJSpGi8MqKYUbqWTsIgaCwDR28Icius+lenVRhTvPLUI
vnlLvyUpfxeFbyLKabes/qwh0iRwDUz9jW2+EbYKeP3fBF6GaaaWh+iRN8TXMGHg
BTKChF7qL6VT69Azls7OrmnE9WYzBu7fm+IoLqTmlhVtMUK6rAyuEQUvkzKra8eQ
ELtlYJ+XMJ3dvICJ8knG2GoF+wkSiIDBrtX3OS/44XwoJGtpFwVctKM3TQPj3RvW
P0ybe4/DU4XwCWlfM+2/KKnyimAtCJ2/oL0O9XRpkOxlEEIvCNAZVGHOAhjdl+MQ
8GzqblRe13T/BIftVtDtMqWNS38Dm23YrnCvFOVUKNdxXkX8l/O6ulh+kSX7d9Z7
FUZcyHWIcSF3pjRQLbI12jfMldlPZbDQ0zfA52MHQU3E+JhX+f/9+7Btxsbynrmo
YnlhQxaG/Te+NG2qHFrihcIj6D8XjMlCfcLcdkEYq1+1kWg5rLd4cLy3dkojfF+R
uEZcwQU97xURMlh2MnUH/4M+8O1WH6kRrylmvCIAeio8HIiVxyfkFOQyVIMECPJu
Y5Q8hGVpwOq7z0BkkluZmZVo+pIejBansWZWC8bJF8WKsP6m87/qeghsG/71fPgk
W0XZc+dOgjbAe2J5GLKO3Ngct3LUzfkWwuHQjkp5SCLhbyo4W5edfnSTT+HpGrG1
YBSjC52PRR3XvA7B1BpyaPRh1P+ES56Fy3TbbKtlPnWfamDJlsa1e4Q0PSemqNM6
c+BE6rutlfwopYO0f8kIzbSzZIPutW3Iyc4KpObeaR3KrHDdYSsUCyFY0C9qVKwz
gxgi2tsOtfmmiHY4jdAN+Qpgk/2uC8kgPyUcNn8PYLkAiUpPV9RYFMOMj1cNjCUP
EmjJhaWvMLZuqNUI/s1bIJTlIwblh1Y8msQTuAH9eduo9Tyz0avS9f8LwgXqDspz
cJ3ySpcL0Th/yhq6Gt5ZqMZ5+Ru3dp8g2jGCDA6En8Vr0NWtGee83FVKFQglFuKN
naQXPO4Ba0jLMk5pKXed1rXDpuS40Fm29XclOf268gm68U85qlqLK87gcFDpRaf/
vMOahXqdc6eHlcqS2XtAtcWhWGRZ2HaAy3Ldy4TlLT5eBuq2LYdiY5Kt9aBlA260
UXyEQSZ7WUuW98QuWNcUass8cbQpeaBClHV0NSDLxe1lDls8s9UbVE+wIIsSlZ4r
tqtAAbeVCS2tZ4ZHO6uUQqtWlxWQYA4pHjdH4v5eId2bM71TGKbsShADDaOBqo1n
Flu1d/rcS3C7Upor0VBXb1pmTUH2Nofh0p3x3Z72BxFQTORtqywe5UxisQWKIfWi
Z9a9OW6AWrL5+j4Zxxms0FtYG/mubWEVJ070NWEvTwFDWJoGP/yzGan9rC+xvFSa
rtLA+nemFTWKxcTrV4YpWXV9xvdk8Ls/ROZy8ichTP8uLjRxPCdSPt7JdtaIUu6Z
/Mxon7z6OGpM3gp8xwDezrFHlxBqm3gB4MWVQ0agoX/rMHjZ4X/Xz0uxTbN5XDzY
uL6+zFFA8/4QOUmjIDZHCfbxNExZfkcTcLZd78UInVEzYxsY7zRJV3Q4eyRBRAev
7cqM4uWPq8ORGIUhMd1n3GEZ8gbRaRrHBAgE/Jbdv145jfTlM2WKn62g0pBvNFFi
hrG1Rd7gdY0HjZtJPNk4oUG+AdfPSQytMtXNZTRsBQDvMnf5cxIDYhfFXhljKGcQ
Pla4/Zy3VIyUQr3mB0QgJd3YwasaYDGdNFGtA2jW0TgTJn7IrdRMODfiFpoZp83R
CDT2rm1A0GhzLPCq0qG+eL0zNzHsxQHiPN1EoYEr7/hSE13Uz4ogRWLcBblnBsSX
24EoYpWm9MYAwEwUHj553DaLbBcXKx9TrROwFgIlNBeNsooRo+QB8IU+zw7g+8WS
KxqFcyCLAhQDhoxJY++lUwaQ73LhqI3/7eoxUtrMTwZm2zJh/EqvcMkAb+EXWmZ5
J3FnDEN/bCzFswxRYlr+jvlwmYv6N+BACQ5iW3MYrW1+si3s6BfDeOvgSXtpoYec
SrP7RBLE1m0Ptaji2Mz9l2JMYeVVPZNxe0SnB+j5A1sbl0Hea9NVpi7GXb8r9txN
gPHFPxK5dmc3HAdvNUhjvnnV/dA9WvxPvh3iCkL+ELn64XENIAlKwxKP8L5PCc0B
PF7e4PpjvNC8VSIN6znTBZyivmaAulDadvrR4WEVR4HYWMoZ0tQm4uu24Hedm6o0
SASPhFTkJ3+agAUt5Ko6fTFVSA3aZpWL+4PJtFgc8A0ZQPxw5FRAzLChOvxL+OsV
/dZuIKAm3sPTdEThxWBRnmFckRy1cqFDFPU2WJaU2uxuB/Q8oyxjIlXZkvkfv4Ga
H50AT+A8I7ByuGes1KCIIwiTT0f87c+3QdwitHdVoJOkCV8/Mub87VyPxIyhi1s5
JxcpgCCrF6IIHsJAuJh4kFeWwTzREyP6qvmbXeTxeEBY/R/xO1s+PaWsGftlv2GT
XQ/UU5M4tzkyG/0A48zjZpZ4ObHaX1yFDo37ZfbRIJ9j/Wbx5CMIMw1JGBO0DaZ0
2BXXoZI8vOf5AXo1dF/M5CYIWk59ZeCTxdxHU5ztRKrhwz7+boi18z/JB1ilIl0S
DQOknJJ8mhfFefG328+EZhKCIqmhlMr2Ad3mYvpSsjv2RIdUETp0bO5QabxvOBf0
wDADcwMM5x76Z5OoQvecBw717V8KtFlAbNrbBVR8lX/22KJyCe9t7wbjxMdIwcTu
3YnfYwr0Bj3SkEv4sUmd6G/mVDnL5lrMU7bRFQTUw16ox2ncuWO1cxhFkT+9OsGG
uiQMDq0J9hlqVEwUrklXmiKmqCJJ7as5CBaNzfj41ws79KgBccbnk6pzgkwTOYkN
1aZ6cufS9jyXN3XpbFXuMARzQK8iPfNyjhzkYGxIB9t1J9pAaLABc6Mfk1pR7fE+
0Y8pUNJ9HrnKUYFC6d8y5P3K3km45dkHOgt88jcJZNNKg4fOrQJFM/oiDx1L1kLF
4UkR7LWZk+CkqtcDHV99aiwES4CxRPDxQ+UdcXWkYOyOJqWOoIn9pOg6GYxtKGgW
njysb/lBrw3WsJBMYCNT9CdXURqZXc2wkZf8H6UQjpimUchvnU/SOBF8spfrYbvO
xoTKBRZfK5ZD7CptXZBJUbf5juwJ3JiINC55Hzy96o1N/B9n3S06sG5CY/vMbJdP
3tKkuIemtUxJ682s7Ga2FL0tpvfBKlVIA9FAcOubsHg3X4XxLh4fIhjtXmIdc/Hv
ayu6VBzIk+S4j3BbOvhAVYAu4+jGSh+y7wp5tcNZK+JDLkyowrnIHcN2xHfoR7is
7bmwuM8hbNCL/tJ1R1FqFBVORo/fw3kloqCETmQ4613fF1O7QrYy0wyQX4O577ff
mYGpXn1iLFnyO/LCZpqLqriUYxlLobviZdSUKED2oREhKS2+hn5pX8qP1eOrsuq9
LwATo7rXRTQpCvNg7fB/Vjm3sTRKx+sQYH0Fp3vYp2acLEFHS1LMF66rHeNHNCKI
61gtfjUGZPdZQe0CGoT2nStcRVDy0rEhikv+ys74WV+BCf9wepxDX+CIJS4OFQMC
jIYvj00aJC0HhhVEU9RkZRzbVfNTSlOSp+OtPRPv7Lgr4WigtDnalgJPWF0N7XlW
FI+VtJPMpaXVPw4fAtlNwPk0hwBJXk8DXN/vVlY0cMCAkmHni31qhwDiIV89Uzki
1bai5VRYkKvnbVB51DYovGwwIKpXmhxYhpjRrVXwj3WupJwZHjeN+QXC78Lc0DTu
NmS7dtwIvNJktbMWuSjWDwE2bhp6v+jcjqOGfO262cbyW/AByX2arStJQyUzCPdY
mdab8iuzo9rE1wuMAE9cfSLj/kS/VPmVHjGPx9v4ZoX+VN5dqYcm7vEzZ3Ma/n92
qeJvSwt+RnnRxAzhGBIeHGd30n2/U4tHv1FAPNQk20bOUcy/0C1qVPSiic0RZhrW
5ITqTGlal0CP5fvnr9kNyxP97TgNatfufkgUCit1cG5owCaBahg7ksxQ8uD6lbht
COiLzPOYRUYMicVi7EbXGy0+w5jDroDxd2VtNU7wsvrQ1y2Vf/F9iRxnf82nipFG
4bbp1vy1EVR9sMn5zvxGO6MDdvrvmYlau3UcuktPZM4zL3xjumVfhmYODgImuGnw
3WNEtYhu8xEOhHsJih3UdokmKsEfr3qHStyntZSYcqtsESR1NXs6wn5Ay2air6Ju
9IXzUT6s5GfkBSERj8WnXC/SZerXk9cHcQNsHSGfNpdBqL90iw4EoUD1Yjhu51jl
FD75owATSunM6V8O1IqhqY40t7xI27z/ErzSECVR4WeNbqP/iGgme26Sft+ieTSG
ft1p4rnXu8IeYtTd422Mu18w47v0uzePorFf6dvValPdLycC8sf/cI2hHQiYKgCL
SAlJafPK0fgMY9P6T4YhPFFCc8ZX2SBS4l5hej4NH9RGEowddx9Yyd9MvLkQkJ2/
eZUaxvm3p7W19wCwQbCsT9H8L9L3w6A+fslLbIk2S/4aHSD/T8V1VlVnXiBI/uyF
B4DZxeJuAHPFCURtRswkCW3+5IMxX+JvV6BT7wtHs50mUIvQhGiWF2y5yNoYfJxi
GHyIcezugm9dhVQT5VtF8U6luwoW5SXWbBtyZ59Opi7pT+BxjXoVl9s5EDmXg/7D
Cku5n1mrLbEWgwGtc/wRD+SqmVulglzZVB8dbqJDWFCuMiwIu3c7qgCVOrY++D91
aYY9gClUzdpAw/Th/oz0YERnbFbMtZJtsNSu1cGurRerKhFGmYvdNYs2+CKftqsd
NjMvOmcADqSo/r4aK5nnm8B6OVvT6rd/WekB9MO5jJNzbWv8lu78+GsQ75irFZAw
7O8VLiqz5maMSB43b2ctAJJ0AO1MlUdkQ5IWim4CPvnxz4wnY8wvWn4XoyzO+qhY
BcpU/nmyCYffnNFdYqMEkrlvbPB8UinAEQl2CYyMz9tQBzFDfV2h3l1CBBHapWnr
CoZS/jsOabd9Dcfdnhekb43tRPYV4yiywxYD1hKLrQenCT/CMi4Gz3DnsypBry+0
dCXJ0i36tSBtuNiTI1GptBqBZmCCoPIfVfh+Ssls4O/vkSafNCDAxzHcxR3FuXcw
V2gCQry/uwzl6ilDzLLw2U7vmG/GhfPG7hjI4xOtlug1P94pWad9Jzl7C+0g7ccA
yBhyn44oGB0XdbGAuPBgFGntY/ib5yVJSfJG4elNfHVxsU0l1aJQNuDvGfZGgG+d
k2swsFM317QTF+038T9i94S8yWAhWrkBnjVTT9fr7SLmH+GCPRFj5Zycqq7RZ5lV
SB7eXpceZQW/YAY5stKAdu/spuyT21hZgDzTlazqYeTWy6ajuyejFy3hDUNWVTQZ
znA7xyoFyoLsIU/PEwzvAsZnGpHEN+sskKohSIn+UhRHHwhnnH3j2kZyWO+qxnqz
X8ApgcHqbXeCN+tATAxqnw48lN4A5pc2wGgaaA4LpEj0hxLW8q4lobaiuWDjjPrX
2ZUV3CU7eA4lET5p/Npla59jNT93v3Qi78z3UNp9/6Db92KSH3q6wsyp0LT7Sk04
pOg/+MY5lAbDdxJUaj1pKXKgvR3M40BAw6bt1g7SqplqBWyIVJvvw2E3AMVS2Tam
o9cTomSIV+7yEomOjlRRCuYQcmaAh6oaoRrN3TqZG9Fo9bVeyIIMA4Ud57RQJzdv
Z46sq+LU3Hjwb16oxXidq7F8N2lK18OUwN5/n/f/SAgIVMjdRg3gUcaDrAS/tWyL
q2bzeLDUmHnE0cTmdTIUwMcFS4UE66z4aiQHxpOvzWcbL7UhA92rKFmvySEY205w
9ot/j/pUeV6jCmCG1tcKdOPjhwmgcYPcruzZeSQD3fN669u4WFPaGBsxuUnm9moO
uCHzk5ATu04wWSvYH6ztAcFBj2YYDApYqv8AxT7VvQNi/Gk7/Ux1W6Dycovx8ylC
ry5u6lTWi6YQl2rzkOa7EWyPljJgmLvJid6vuFvsSpsemwSG561lz7W5yjblwCWd
aSbsOlEEyJx5txpApdJNMRCEG2p8e51CSMEfLrabeVn01cnPbzj5XPjxS5fhFIKm
l+Ls9cOzqbYNdY6DXWWPTmYMhAU/sWZephQw4fRLBZcuP2gKfOaV0mgUgOqkTysz
RTC/R+xpU5LFRGfsIH330rORrDBvD6rtxSJwn+Zh5EyKGtNZnqZAes73BzzcbluZ
9rpUifVifKoVGsu+x+rxvCTOvkAtazNuChdh/QCCMBKuTOuAcdykf6Ii13LtdVSB
5B+ew+L0kDrWcYx0h0+lY8WKH7ckJ0NqCpq8xglg/RXADDOSEc5opF385GHBLHMN
JLIHZaMnf46//PNhALQ8bySOALDXQBdJn1XsvMqL/XpupxU8/zZ0leU9M/adieSU
Pj4V3X538T1lSUU7ljteh8no+FGK7NVM4I6I9moO5zinH/YpOGhv7bFhLstIyLTv
Rk8N8/0dbbZ8VEQ2B1jSo4rIQolffeZ6qRuU97NWG3dzkwHD3jHv86/2DIWptqKr
e+mhmGfjmTch9rGoFuv5xYa33x763233rossZaLIJ+meyS2eLCTv2B+5KGhKBVNb
sMEdiANa+41jO5j/m1NJhVsXemEsGKRgqpG3y5yKaMhWkm03UNW+CHtL5L1nyEUO
G0ST16v4bIdAiEIJWHY3gqFdEPXvoTxy+UAvCth6XmvmwI++A1QjcQzVUvUoFD3e
vrauFFyOvAbscBhKbNH8FKvlpR+8WjFk7zduRVcjd0wuHlIJGXzzfVj67mVCZ3FH
s3P82ZfZ8BR1/e9is7z2MiHc90XP4m5ffLfUIL6wTTPDmRw1EULeDgz2QYiqcAco
NgX1xRIQpF2c9grjd7N9w9TcxzVvVRBm5vAeeOGFhXP/npGYINxHWII2xhq6HTM1
936W3jFNq2IyLmrYDRlfLliNGC2lHnYon3nU9CRO1L5uoA5fSVLK7DkyxVHj+5yE
xBbPiZshZoxV3zRWT0sfw8TzYAQzkbsbEjLmK7VoD/Cp/ay5jrHhkEJja8QvvHeA
G9k7z6/tiefk7WX0Tf8iSGljLzuQvr15su6/bI72E+O3RrcqN1xWuCfkNKIvaMIf
Q7XiyV1bZpbc6INV16m5rKpnM2IMFaitSOHHvsJ8PeNkX2I1en8BFUw+N/pFhvf4
EB8UsGRL9wd81YJes+ejfdf8jdCapGcn57KgiCGPS+HqMtHinKqX3+WK2GSRgA94
+9qvNZw+DiqRaXBc5U8b0NOrRYdZEDsLPMdWD0YVpVx81xjJrpcNzhrLFis4RY8T
EW9HaIR7RVOJRhV34a/ET5ht0AoFvUoogBRPT56Tbte3puhukGHhKtZ5GnIUtXE0
hgQk7xm+qltJJA25ceWXN+LZRusqy8OLFXkIQsDEXaVwJPx4A61Xx6udP/nknkfS
ZYF1k8blsdUu+sXfM+/LsUjR/JNWGUABmHB4Ddj8gyhhBl6CI+06pSrF6VZqs1uY
mY068/X7jO1/IZKFe2d1I2LVNI4Hfv8sInj6ZJhV7DBZwmZjR18jaoiFMAfkQcwi
bRZ6FpK60d7u9MqCbKJ0wJmzCeJZ5FRARGJn/f30EVtcj5Df7n0vETUZuhfUzJEI
IeQFzIqzkgFInO5FuTcABVStvblFb0UuI2eyq/uQwjbrIK9XAEr2I9L4q83vJGTv
WXuOcZMZX++Hp/jURIjVZfzMjGH0cO03jG3QeYo6LDIiVd0lpABC1fpoFvQyVqSX
iogTxQBQtnU0TcUc6qf4dhK4R6xsjdHiNrdLE7Gzn9DxjCf+SuO5UM+fOcLeD7Es
Cwkk93sMdbpCurpBeMU+9khwmgpk1qWC/h2bbCxUh3GgkgTGylJ7gPwmCLaJ2Mwi
XsWeI8ygqAAZP+Wxbpi/0oTxziICfvq9duPtcWzrK5xZTdh2e+3xHdo0pmfq9eb+
U7aYkCO/fbhEjqbSe8KlB4mbzBRdCigXkH9pzWDPTSZCp/kpwn1gW6gAKRYasO8U
JOhVaWczCyh7opmKM3kKJmRdQ0flMdyclLfLnFZtPF3tq/kDbgSepFCOPrhDd7eN
GPnx86XHnXHP/Ib06FoIJhK2lNwB9G+S7+v0Q2PZdGyAFfxYWwnoTl35JnEeDg6q
+akcY+kiCoIAJoUJcu+/crinEOGxB+Z2fSxsTl4jKQ3jWD19J380DuknMl2U8RgK
MVSldBmV74dDwN7+flK9W0ukA2gvpbyugrocVLHjvhK75SV+j2Ml8Ze0tF/yxyPQ
mhZ6erSR6tGqMwcSTRvSslw3BOcKM1coXVUF6G8DIebUNbhOmHaS5TwrLignegWM
ODTQyVqK7mFx8cSUefeUMB0WRYAIBctkE4ZVAY2oP6x4vBklB5Rdxw9+TeLkZj7H
rPKGDUT9IXq1jGosOOOU5xo65pr9i00uArF5JbIEEoQsYO+gqq4ggEjU5MRLjouo
Oe4PMLfZ8PgKxBAz6MTDuavvRR7zmQ+o86hYvbuOH+d/LzT/7Hh1Q8ixfWRRfRMr
MnkjgSk9IfiphV02z2iHH04WtWWgED+kC13mthnUfbobERjyLdn9SOtjeHbARCak
btdgXnq4Olzf/iwPKL+lQIUrN/nNeYU1EkUjOqLh9Rvj9qpwt0RRxH7OUnC0SSxF
r5sveOGzB0AVWGhDowSGzIGiFbr2WBrmd650BFmVXBsYq7E6GOW5eZhZpX/Yqf+o
wh3J0neme8AaZa9OCqwk34OPF5QIZp/NjZCM46BBin/m5+CvB4fm8IhsRzr0Pu2o
/2j3Dxyt33uDtRmOFjd+28BYzXmFf1izA7j80vkiu09mMkhteijiyoB7IWFKKFF8
50rrad8/XDLxcrjM3vmCuHWny8JwnkXOdufPjwnRIL/F3yZJwD1t3+kPYy4/EPSz
v9N6MgCo2OviHk7JRPoet6rjzwdvxXOr/r1G2LLkrYlY4bIYAQcJYyQKtRG7bCOm
xtOOLbnjLtb7wumwTfo9jf/EtBhOPe51hocL3mReXid0QBJWhDLhJ5xLDUKT0uCy
JedNrgqbJFuusiYlZE3+YMtgP+ZOaDLRIQW81XuxyYuTmDogEdrgPEyvl4EVeueO
VoKfbzS6I55/FRAEKWiK5jlWuvZwqlOsT9SSpaniAJO3qMkoJHJuF1D8AN/lbm6d
d9EZWdqSSN79vZxIOji3zTCqKq2h/EnARkddEcSRx4b2VnWvx5nzxxl9hesEEEnK
gHr5NgzrfBkFD9tLQALn5NgIEa8F2mREmyIMAZ3dPuDWvaDmnd7GVdPjLPVisqn6
8ZJ3AdkVSkYqB404pvBwDwgNvGfK1IhWcbgMvmxGav0B9mrYebmWfpBWiPWCKaQf
DhhSiS1FX1LrjUFX3nz8pDnaJ5WSZW95bqr/yBb/YyX8sI719uBU2b/ISaLg+Z6t
i2MuqtrCUQSXnE0V2afvolPuDkf49shFFe3VP1aJujQaCwNr/PzET51PrMofm4UO
gY+gB6VCqDvKevYIn7+WA5LDK6oWtiTBiZQgP0uI5/NNj+r4IF9eQMy33AYziBZT
WnSaPF35p22GTJgv45WWL7+YQZPvfOjj8UBO+i2zH1af7NSCq9Ev0I/7Y7DgIX8c
8xeRBVz+glOXUyOK+E5N2LU9rqo5aAuHJ9YqnbsQ0Zu7NtbgNSQBq7YFfzSzsQl/
6gCzX2JfU0mM4p1+Vn6xecPOxIGKppklfDLQwSeValW/zuHe+WQOU4buz1c7ISSL
ioEI/LuJ0EqoFqxbkUW97UKBq/bLEuzwGO5w/t1IiBFYYAgm3qjKvQw2tHsXQEe3
I9H/OwkQkSztcCWKbK6DSX9qfsbMwLI02hl/mVXDE4fQ5xJO7R6JCdfh7AuZGsh8
wE/t0MDs+LFgLrlRh92EG7r2n3MNMz9cCVaAygrY5CE5IJRixhnQ7DZnF8pQrcs6
gmNcQ4aZuyxYD8t+Gh/UMC071BpiOuA3MCveFcOiUgTHNVCg4rFGhTxziCeSx/mk
4y2f+oHeGPTBqpTAAH8A7HEqr9YQ7Ji4P32JMjBZUhd77tkf+UI4wy5UIKCum1iO
YpTr9uIzS2Eui2anL8bQkCc7AD9BK3VKeluMkL40y088l+uBVmNT5/IDujVjMT64
rn/74XtwN+51a5GcKFQYZeZf2G97vMbOlt7Sp8vkLZ/3tYcntQUroQLj3aV3l1QJ
jjZ1XDrQI7IV7qKVfdryf6ScB0izM9gy2NcxLUdTOagP2blf6zFNiR6EOTJOMzsw
jRtkHh+Zu9WkurypMJfbmAK226wC3nyss28sdGYzEc1f38dBzZ5CFeZyXkNXfasl
52g87PfB/kCsNa/DQIzywSKlzTm/Bd/CIsp1hii8JFSZ/e2wvMPlzeKyfCcg9iEp
M46KBfTQlcSCbcOXaqHYbCT6q4IZq8Dj9i22qsNCT8drFwTI+Xw1OFnyr0g+tVAd
0WtaFTyHaYkkkT666cA5m21xjvs2dE4FyLphmJwXoRGn/q6AXn4jEzPY2eFWQFlo
4rucsiGU70swFwW4JwaYNRdYDplHGgv1Qm0qn2340zbHD5HBuZhopixKQGLvKADL
UKgelltE7Zzo1QJYXsRFL30dcfgf7UN0q7WbfEX02FvezJImDc+H1lYK2KiOQbOx
aRmmzBtL4k4F+qJUPk93c0eJsp0H03cmNKFkIqZdl3P/tqZB+fRUz9OcWpHtk5vC
WOszCTnMLLRrPUQQbv9np8Izivme0sGJL9EW3zMWXiPGD1L9ek+TKfSQIYYK1j5P
KljrsTOr4TVksv7kCUvO0t2+kX1RmhfjfLrXnw5BVGSHd/8mxOCwBql6RoQYeLQt
PyVMhqltCRYmC+xjkR2n8AtKKzEoHVdTJw4R83A6Jby97mqeCOlbQRrQLdD6RuDB
4sxRebHYU5mi7BMDxmRgO+d8+1m+R9pHKFZA1WkhwW4BRIKVnGeytVt3VqPta2qT
vJgqLHsep6/HXGFY70nlSy2g8atuU+OtRJY0k+Pu+bGonmbw4P2Gj7yLVDQocA3g
mMDgmRzjA+uifA5pzJlf5ob8F2HH0LBMRnfZgu4U1VWn1Nbe+4haAO8yuHvuL85f
6lEc4vmqtpWR1CYgmM9DSG+asUIv7HkqmmSC/JRlpqc7DFHcfTRbbP3Gz+bbSWgU
6ZH9yRxkSrBJVYWGz+P7OVlbuB6q5OymOVu2pp31ZVuv11/NXRhyGRrQpBhnRz53
kfZn8Zad/rPne0MtDBH0PwfUOGBb2+VoTL6CsJtLxFxzq0xNZWBhZoASjDadThU+
mM43CfKfNz63arOjWu16mP2uL9ZKU+o4Rntmqh/BWm/eYXO45aIgY+hD+j/XTsk0
IoUL0DD2WINDJzKvGXaUV2HBBlKqVQ1jjhDbI9gnoPw9ITfS0317MNiE5Cfk4uSj
x08+eep4OXnjdKGhv106tr6Nz7emZ9n2ukoWhNx+QB/nkNRuPYdLn2Wsgb+sdxyq
RnL8Q1Yp6OwoZo7y/lh4zcYHY5NQEDT1RLD0PierbngVUrOLx7W8x4UZ2XdBXqfr
J3tzgXRYp4h7LFVjh0iJBrnX9gYtoCJJgTW1BXSBw4QPR+MJ10UIUM2Tl0tFb+rj
vY13BZNU9wz9RhEivvnoisekcfZlG3uit56fCVQSAX3KH0tCltMk4STMwNpQHmO1
huivmQhTX9L7QgD/3ABepWRq19qwlDtMn+Mx7D1ApRekTPEoT0c8wQhU9TpcC0Jh
NSIAV6pKTo9gzy/ffzzSrlX4CJkB3KlvegI+dj7LhBW8wTPlkJhupSDCkxULrazj
ljBBkbKynrcOpXI8aTPr5c1S8IEqUyhIX1DAihPqSqAxqkmHsrRMUzFIxQgvc9MO
9vfCEmMRiLNtYIKOwQL9JjfYZaxtkUsToKSpRakj88ePNN0+HZmGH+0CUoKfOyh4
eiYkc8N/BTmckRI+LV7X6iRYy1+ieiebfT6sZUTOgl4Aiy/3zsQaqq/THscZIwgy
fKKQXAqKvnjp15odd3TxdDS42ZIub13cwMe57RnXMUEXl6Qv2Ans2M86fuR+1JF2
trj7SYLRpEZKLN2JL5SkbI2gi4EuPMh52EeY5a5jF0l7SYHZDYmnWh2Ey4n/zfpl
77/yzdz3ChvFwvG9k6JTzdLzSxasu/AllcC1LRzrh3OpnGUSs3af0UOJNPmzcUyU
UbZYqdA/AJI3EvnDJakR4zC2nalF0TWo/EGh9bFs2Fptm+gzAG8J4n62BoHvwB0n
PanVKZdUF3GVG5IERMCVzOKU+c+74Xyyv6eeFEyxjAfrHR2rbK9180/4JWc13fc8
sDCGsWsPWuZLZxy8RUu/i1tDfKz017IsPe3KLytl0cjMzMAjOa1Hab591hA1mG8+
hfVXwFGbZNx/G4PJKiubzUbNknG0ESDq6oorMlOL9n4+dwzNNZPmP6sZib1/2ARc
9moftQ9+e4hazwaPqUv1cOsC1pl/OyYB3QjjINjkBbk7VtkekeT2C99+rZxUIWEa
JZe89SY6cUCc53ezB8vyryBNwQJateJPt5k4bpfCepMtgvaOxs6iH4UrHntYNyUH
5RasAWtDdxNe5GN+KMk6gw9YgWm2twg8xZOXtH6BA37lYg44DhgQbVWNW+PzInHh
C1xS1BYFZokHF4SAPOhh3Bjqiv6jpowBhttrqYuHpWqvg05k0ZT9wBRjBlFZ+wVV
FcueNdLTCffMN0sDlpDEDoNOSq0JofN3SdY1UB0h5GuhXn4jsT6su99GN3xaOGaH
swqD1AM/0yoJfIpClnieEuPVbfVysdwE8ERq9Pqs+r7jPwz8EkkiAnadv8XmGftg
W7AjF5DHVLMzH5V6KwULX0iShXETtr94pVEaR9XtAHyMDF8/RyO5Y4IBexHdRLZm
+dOqD1Nq/91nbdBHZWfxWTM+jo84x3FYhBKSue9jA8NfN9ivBhfVh1uoFNyv04SW
ycq89YY6Jt7CddlvEck89SRMsQbeiWo3VMb7wBgc6zvlM5v6jOD6etgGu32ayVq/
4vTjnFzcXTC/zOcZmm+HMk8T/UtU/W7YuKIMMlkzEYt7Znujj5Gq2V11QzcqOpLR
KIcbPV1DLGpc1C5Q9+/KzqSgAcKWuT3hvmL/BlNOFPMZEncOIzAi1SvVJiKaxIBx
r2XIIjLmiowWav0XeXGgzF9HoVCrX3PrSr+QdADEWSseDvLwGLmwaqT3fmsQ2OBF
OvSEvydzIeh1fkqafoh54EgFyO1f/Wd3BK3lQZWJLkeKqnr1gGvHUJTcZBXD5g2q
Bsbvgs/ehO7uFGk1xSzA65nV045Tmwm6uOBCj++cRebnWm60fJGQc3t1SinOaPCf
L+Id1YpI+DkSP6fIcm6nKiOAeD/PFm9tqbqj9uh+f6PxTuucQQ13UPZZZ+QQV0TR
dpDe9CG0rpyCE/4ulcrZPA==
>>>>>>> main
`protect end_protected