`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
8aCqQ2oUxf3QHZjuYP1t5OjsxBy/GOS+iraSqP+jOUUqJHNSRnXv2WxIb3CUWZqg
IQb885eLT1c+iwjnK40Sbp3d/I47Q2pq+zjtXwRVFkM1qKMdPIMrpZ9AMX7MuMsl
aztacOPLs2V2iTdwjuTLquFeXNlbR/HagebbLw2PQUMb9r+IHZIcZfYgB1bDBg2e
8CU0gCOnBaHvzqLPRSrVFWH/BZN9u5b7umT3L12Q/7tUMxQ8MOUg1Uda72gll5Ii
CGXBzRS1bqKtkYCmFgWFx0+3CpaenxbDxjvd1Bqm+70ohU6JdBZdeBiLqkDXv97+
wJBhrH428qlpKRkjr2V5TgdtpPraQp5whqm0qrgJuspvDENaHSYT6LGi4owcyJOV
D+bj57qIPBghm9tAWVePRZ757zZynD0qrmcPgAUo4ayUrJivhW4gbmp5+NoMspvh
HC84nk2n5n1jHK+1SJtrduZjyhfrZHF9bf/dZV+tgsbfdWXjiQMwUMVzYqAvtupY
ZsScEFFc4JQO+xo2qzx4N9iqTYm19/kY3FMrcc9rLhY/3To9VqyUREqxxBkY2YIj
i8ldT9CWJSbFniS2uo8YUityuOXB2dtwUDwAkn3bTFdqQTEg2CWaL/V9Jtas9bI9
bum3k40tyhrlbh0n3k7vqJMuv4gNGurjEmcBOs2la7U0GPvVHVKJAJrZd2jXF19w
jgR3VDZly/GsQgA6PGip0ZaNHzs2f3w5kwphLb9LhwjFVlf7G+gDMfeYiIcQ3V64
E4R0nEuhOGGr4mlCTMNP6YrWfy5zqd+44/HvJjtWVjRTaGMS13iIrbSHkpJC5AlT
4jMzBQ0nt3vq8kWT97PhDsfm6/NjvJwafHkDm7X23klA4Me1F2dKpSLu4pkei2Li
C6kE9/vzu3q99xlK2mxZz7dNpRaYByq2+ZWpysJf4UQluX/rKzZzrNM0HLUKHa3B
SsGTdkyT0RZN5URdMLZwE8LNe6cSTgDIIYAqm0vgX4jYMwOXPgW1o/v3CLCGdbP+
sbayULcXEBzMAPJio6IrQ0gGRhgbpMeqZ+p73+wBbZEyAcqeOs5zTpFiRQl2cNue
rBJ6CQbRm4ZVmYH4nQWytkUVIHcjpLtvXoMlLqkp5xa4CFDlk8AgKhLxce5cqwnr
O5ylQBnH2aQha1m54fqO9EqgjGpnU+rf319ArFe+dQRhAyuX1koLvWn6OagYVCPA
aANI5ZQ96X1HsBr0c8Lwd9dFnJPYVkWpXO60TKT/tor/OrwEngqYLuWXJBX/Nt+k
vY63MBtlDsTB+fO7h8zRCwLqdobBZEtvCgJiaH/zwtKg8DjRexY1ZFT741VFZj6Y
bz/pOe5UJ1eehj5FUGsezwAeerAPNJQkwx1FClp4hAeC+Nynrg2g4ezctTrpDYqI
5xhCCdsKFvdgc8fRwo5nbuxFev8/C5QpOvCEr/CIAfnos13XYw1auGR+s0UjuX8C
jW/d4C1CAAy4jPy8E+gq8dWaB/go7/+ohitY3MqMKH+DgXSqJNtjKgParCqzyOw3
HeOWFXEbvTFSf8ta0VVdki3L4KZGOu8p8LnUIL9PoSCcvI9CJqGjXHRLS6dIi0q5
04uTVFJmLxd0QM4JlZYS6mE36pTBzu496SxLSNBsoLjssmhcQF82j+h3RsUBySI4
WK0KU3JeDW+MOz/vbq5DEheT3WK0WpC+yNS/SNwEsKUZ4Zw6e+BJwyTo3wDyHX3J
AoQUAQ/RJVdtDOjd2CQ4vL/h5dScgciamLgJSWwwjIQCcra8v+9vZqppsAAMnmo9
hwG54oHNGIeJaPaLOtW+NznQN5gpl75YAVRgZoEPFxJpbrSUpG0Nz3fL15ad1ay3
9JgnR963olwWWMD40DOoKh8JCKWelVV5ZrdQM6Aa6csI3M0rH6d+w4W5PVcxjowd
QDG+dnFDGvZmv6DP0kCnA3G6WZM/ifz2vcfggLSWENPz83VoyhQw9ueiaTHu6t18
t5ZmybU7Ak0UWezWQ/fze6PzAQAX7MPqwueYtfUpTEpJ8MooMwIXyCOQKniN0USE
daaruI1LbkilPYrb8jmo6xOCUgAtgnlnVennMX1hHsN7Gr3LDjOnyysJ0MBMqeUw
BvVxa/d87W6ErFL49R+X6Dm6eXaHCNDnhSjzDnw1ZigiJl6rxHXr53warLxpyJ5+
zOo+510Jb0k008tgN7DNfqC9l2FbNrfbRxetwjigEN/gurxq96KrsZDC8O8edAw9
rVxisREU1kuzlJogXa+k3RDPlMzwDknHHO+alVZYeYxNkmBQCprehgx9M+A+eYEy
E/Y/nFEcMhcv6Hiv6Upmzj/hBaA07ff0hGL4U8e9I/PwrjmT3BGtnZ7YJJqoMMPr
98ICVBxaPjIOKNZK5SjWzXhNALEf6xn7pfH6nX3v8E+BWSvwavBQgPJNpS5ENex1
zpEjIo5IJGyOmrbcny3LtqZFJgnI7mbTUfPJGuTmPQLG32ENYEFThT7xV36LYvXu
nCy5vYDZ8YDHBAmA/bdqU1Cl+wFG02GL6Przf3PR02Q9lVFj7eAQ0TRDecNYoNra
qFMk2vs0e1fOLXN93tHTgr9eBs+tOIeATPisM2KTeB3Ciz9gikR0V/ddziJ5Lp7l
PK/JsAhLA+1Oy9IsuznElo0+m7tlyh0aMhDiGYT6mCzFCFiwx7f6vQOMCGR+E1ln
IVZLDw39dYF54YjusiTde8eToPrf8Oyq452bDCxJH7MYFyOLBVVd64Imv+OnO3Cu
dPjvw4j32CxoG8dr3B+dd5Qwi/sY2kTV6Y/5OhtCOJA0aaOLI58pRuW62tJPDvZJ
b/cZDSMrPVzl7HgaC6qreqVkVxL8yVLTUvQk1ONXahrzjWfrFQFNiBhWub7o7TFQ
jf3j+wIh8x/OwNBg/++8nshxDPkWd1dPydSLjf9bN3JhIJTvcCknq25j8vuX/OQV
/fDRUyb5/BKrcNNKIVQCyzz3L4wl/OTO6tu3tCuB1dVdgZBtCCzFVvKx+d6X0NI5
PVoTcp/rPxnXOJTkLy6zwsdmEbZ+YrhZIFCVz0w7br2bzFo5yLj06BqjxEA/I6N8
15Otw+VLkcWEbcPCpfrlHTgyXpQ3e6hvLGL3Y89/SZ7V/yiSnFwpdCoS2DrsHEQr
b9UncYSXGsT45vJFZyOsfW61Gj6S4OroK+u5DFIfmrO+mIiIyEvWeG82bLBWs+6P
w8RSYiyTItHaU/pY0zbXeBaL56K7wwilvjKWlwIeX7ptcjisj9ABya9pwzRGdBrG
toeVI3uJDgfcBxAzEDQJ/3fc6OVwrK3BLJ4ulxnogVOZ1yoBZneIhynwtmwy5uFk
mg8lYWEudG9huTSQhq7F2w//Haq/f4HN+WiDCQFs/hMWzxEQviQVQANWcm2RleqK
xIDQPPTMwlUw0hyfsb44dnmYztEdLPRX+R2IVvelPfY1rUTjF0Y6Cksdk/LWbuYl
cqH+Xt53GcLn4j02PzQrr8we6L2rP3UHRsfSRl0CgYSQPwe83ZHYDBn2jxykcPbr
qLGXF+WixkpCeOazqPogbHTmu2KWcqz5Ma0Hz2+1DXL9BqxGthHAIGhQ1gFzOIsL
sIS5jQVPzR4iahwfXNG4lU+i8CesbpzZ6rsuxAXoOVP8sdGBXvNL9GVR2QStmb13
XNrc+SnBJgBsPxaK37/T2v1YPSIOc6I8Fxd11wY8AR2WKA7uVATR2Gtf8vo6rKXD
N7u1SUIp8vH3164AfvvpThVM2sg8xyCNoXKI6in49UkSlJBQF+Arrx0opkDI5DJr
/EMekloqgZA2D5bw5jABRRK9zn91nkdTsCn8wfjMeXukoE2s3WgFILJgt5kUilBl
zkaqz34KCXQWE75oLpTJotKb8f0VC4Gj8hqsHPGvWiYcERKGB+phXmqzKJ2Khu9s
esvBmMVOgZyPHaiyX5ebC21wolWflfNB7eFUMQHequ0fffwkqzCQWvWr74Imhpn9
/HOAT0WA+TFkahWxTytuQuPY0JUTUXG9cfmUrDJcW1GVcIvfFd9APdoAPvHzs9iW
4xjGLwVEc4bcGFhy6cdL/0L4iUMcWn3UiYCSAbW/3SP7Lse4lxK8+4Ou+fJ3UKEL
UiRZiE4Xt111SNYMbM89usEbP8i8KW5nD+5TTvD9dnlf54kPSU36BSM2qSGMIQUL
4dBRmtjXJOXB5R1VpvcD2arrOPlu3uATraMxYDrROwmWCnZsiv83j+S0qqzkGKSw
aQeQ3ExXYrixmL/95SbLcuAHOVttHcrOJPoR2B5L0fh61508QzAJSUEQWjwtwlrZ
ZMBsySip4PuYsfezns7XSS5IguIcLzTbs/w02or002/ahMaG9G50hcMyeeoP9x1e
+h25QjU7P1kdETgKexXprN9fNteGnXN31zzMDCFMrkOR9bYAGXvVm8mEv7Smdmbc
6trggrldvGBSTmABPhC2lUZTbupxrR5Jx5IYvthF5C5vi+BxR+u7CgwqfDGH7E/b
5nwOk5J/MavDPJXMjSBFwR2/0vsrg3iPltvS9uJCB7B5sXgSJPpLRMjxzODyfi8s
Q/LoGrWxErowthEZG1FkyuC9d6nBzBDpiR7hzE/qAcgjaCX4FquoL2k99z4aHw66
JZiBGq2osBHMi5yuRq5Zh0kTFWRqkp2MPq7z3Ly7MuixdtsZzHfOHICYH3Z++uux
8dTy+lnZSU4hzqpy5r6ZhYMWgf9PuV4AmMNyqFNTCSewomPMc5MkJp8pPPV7Y8BX
2nqzOBzNiXUvYh5VT+mOBwZhAM3TEXbBaqtnrFk2edX4zmf/yvHM7wt5nH/uKMXk
2Nu7yiqJMyXriLBAlzqeuZe60tesTvZr+FzhH11yyXI195arOFI9D+PJ2AmOA9/y
ENDg1rxEn2c+vwKR3QGRwK3jXXfYhUKPED8qKw3j7XA8CqrvAT8HZ5PirI2LuaPn
SPqijEPdVAtExh948uB1JO4rkNCCtRjXqwhor+ih3KXoQRDpB6KjE6Zrdk5I9lcI
wY0HKOwwLaoH6xL1FkJTew04nNAphAakS7JL20tiyzzwtagmJ0LKneH9hZhtJUOW
lyx5s450+3Hn4HzWjzysViH1Hgtc+MwhoO5lIguUfdvRkfTXdEpurxKAzGUCi+4C
tNQyWvOcXiCZxFJK7jdallA/V8MTuEWRqt5vst5jFkqkSDsY2SGDBxT5emLoMzlm
Mq2TVoMe/U+SIiCVazznra1fufHJc3GpKtBoeYrJglDGjEKsqQub3Bfe/WKIFmPh
a/DQdAUJXi/b5pg/PsNnp+Cj99ddGqmnhbYBIq8CgypGtqItqOi09qNodR6Dbnt0
TME6jQeJXwvo4EeLPDseXdswL05Earq0AIokGUs5yfGBrsQ1naNdouBS2pARXV3I
Wtxbwjs/V/o3FoqGqByg+0FcEpECjXXXpoG7uAugnHLDj9GSvd+9SXBKBbKHAuyj
Xmu/RhW9wM2VSMPmMZhXeGkn3ELYxCkAeckH6Pzj9QH703Mwd9Q0itL3UxU7U9dC
D5TZUjzSfYWtiMjEuwEz/Gpmod3bQ6n8+xhQ/sovI+D/oZ1PVYfExDZGtkazFn4m
FKJgXmY8DxHh4QCXxyVgzjL1m1H6NA9VD5y5N36mYYVQb302bVE9Hye8SEqYGFjK
qnnIj4mycLQkby4PpAuEe4gnCfNs7fY2rp8DLh7aPLxItgfjjDihSNM1ca1+gxGt
X2GIM/T2TLMSQ9VYkHSdGUBwNoiDyCbXmTJZXhLrZnpgMm8v0GwaGQBQuF85Aa05
9jw7J6iwnpshgAQyxG7ZTajQ5u4oxgN5nM4jh9p9C+OEkWMBz9kZJg8uvDizcJwK
WzmJ62E6Qfmw3Jkou5DwkWno3vsvpi4k/3S2wHAXA+j/Wx4xEmqTaSVfBq1KW/KL
uUx+H4ofvgYmX9A9Tvc2Ccm4M9s067c7MiaasZrTNKjS1JFC7lrbs60l1O5PNroc
UMn+x2JPyE4tOR0QoWND0gacG3jtgme5PzVNxDCEsATgQKkBBGhMYaZP23V1DLRd
abO0GHEPiSWecPMSlmsAwaJuFvUnn0+MLf9Se+dRlVqI0CeEljZbq7p0mXNZTZx+
oI/oErDJYqpMYmcntNI/AGgluQO5pO5vCOU5S2HPZLwa+2KWjI2pqqTDEDFzHC8c
BwXIBL6P6Lej+UZCE6z7R7B9cK7GqPhJ29hGkWQqlcUSOmvTRt8tkWG/dw+nl2oa
uHWgRLM1bal1bsjcoixhCrJQDF5vXvnzKfKJS+IO1oiuzDA/I+zDOrRwVXpnXgaZ
j8rdOiEtgEtMQ6RW5hVrDJYfWiMG/qyLESRbefrioW5P4CEFSpfJRjBuQtj6FFKo
IsoIYdmo1ZKRlVrrX+tyB7OrhzJSav7hL11rBpZ9By/RZATZLrEvqVu2NyhUMq9W
Q4L3vD1Yfi0IfJFKlO2U/puZ/a0S0Vj0yvgvYfzCJ8ssFmV8ThsR1xbH2h7GuaOh
4zqXjshaiexpYPvqN8u9DKecRBaNLLMbmru9fBi1ifY4d8raN/A1DeR7GB8zr/06
4LADuR9aJ1mcpaECGqnuvXGrGkiSaQ9Bbl9eAMBy7Baun9Z3/DoS9l50B2xCFp0q
9UTWrqGh+0fyZhQZKHc5+O3EK1DX6au67gEcAe/yfYGV5uDlZuDeXfauy7cqzoYP
Pt5AzK7TvshsQVeY7AZL85e4NiU5KkHqfBnSEVDIHGonCX08IFNd3N3Al+rdHUaD
7uS5xEKwSGENsV2YjI+Wg0k4bSmj3/4yGNW2Gu0br0Js8UNR7V+V5RV6puiciTSj
DDSYLr6NZopeSjO0acEclDq3oypN4GNcXqYW77bfwhC7vu+unS6x+Pshb/49UMY9
FZyGLFtHRjEsB1ifwbqPto8KAzQfagT5e038mOl4E15iKhnIpKRdkuCtWSTcAjMr
D8FtHTMTgMoMt1O7Sbvzn1i2r1648UnXc/dT2JVKY49J/kAbKCHtrRffxOwTMN+Q
JGYlbDEn3hitHNZK7EXX7/FZS64C5V+2cZw9wgW3XMqm141r+VKBClCjjtZ4iMaA
p/uWq/CYLtRV+2gb0IgQ9jy9pKD6NN0yp7iaGN76Oe8=
`protect end_protected