`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemKORsCE2vXewM+8rgGeNC/65p4uFaCkBXs7//dzKcQ3O
7EW+JHZ0cPiN7sYcC3YpkGDC6hkSKhWAl5MkaPvYlGJfvJc2jZArtWHnXNYCtJme
MmvKe5ErzuFshZgVVxytQldRmcX23Ki2PeVKa6HgGOOwfTlXPFQZ7GmzWdwY8aEp
coEQWJSKVjd2+sdfdJ7lPtuYanpVV2lXb/bCliNDmuZG7UtBV0oU9hw2ZTN6E/q9
eAZ8sxQ8dEZ2ZLIrhyuF2BsstHsmgaktde69jUdUTSKVPob4ZwTc4SvYK484ygpR
iWunZw4uUt14VVYmpJEktsFWhTYTruL2uxbq/B5eduN/mOXmiF7IGvEWSptnhB/G
Eb62pB9vPto1bD2R/8yFyR3pH17oNGaXr29pEgk3eh9Le5EshCW446radZaDf9vl
lxUDykjHoQ9kA3a+pfY8z3AVq4X9KkBq+PfOxR8ZNF6jt9rwn3PO/ygq669YwRg5
EUaZCKdQmho67N0hxDeDEENa6tHRubo5m65mmCa+F6cMeWau1TV1suGjAJ0RBFS6
D4A73C2LEbO6N/Xyyi2npMP5SFv6bzXi3up6ZMs/5v2+Fbo+G9zoGIlxCXPq2T5R
jRPvkmhSLZwBvFuwnnu4tvGU+32aARwmh+pB6eQeoX3rRlcZUCdMbTPu7qYxU1qf
WgQNk20zp8i2wloMR2ZFpYGrMYHltXFLLa8gQLhwUWB2muix92kLJBIOAlYW5MTE
PI4ZN9gghlgpKhYOaqIOJE7IR5Ngoc6999LdYW9zDNPzmN0agceKrlBfhdTHaH/m
CYgO2L852Z+Ztev7VqLaQtyUl4QpZzlkV9GfEIrVJBqGIpX5ix34KpeQO2v5LVFg
SPkNtOQYTq7MuQJZxSSkPwdMST0T+m4TTHZCXx+7TmrbU1W7s98XNK8YuYEbH2ja
Xq6DRbqC+iOAhOjW2vgq/8sXoXhy8WdOKSjxfrlOHgLCRIP7Kby07FL2ZN41iEDY
d9jNpniysK6vjh7vfx9eqjXz5Ssb/GP+9S7kRBhNzZGx7wfPcj29izkPKm7L2Q9z
qH/1zZM7LkIOA/vugCvdtet5g1DQKKykJn18C+Sgzx0xbwA3PF8C38JWwaDehfo4
xDS1eEiTIjRU0ab2i+q9kJlJZrqNHXB5lb0DJwRKAVTHA6+ipKEuLZ0Quetvzrt4
njFGJxhBgmIXJotualA9Oc62e2WXVeO7KincaUQeg+8L3k4d0mIXvr3jsi9ZgEJu
lixR9z4z6A+DzcGFjcn5PfrxezWC1lS42ougXmf4ZWoigRl52ThbL/A/TKJYzprv
fKkbyk+PsLX7h8tVQteFoDKyIPQbaN0OrIfsMBaMKDSXSJkEg9MGmvczINWUZN+Z
wOl+iuscp/AvqiTM6mfMuiXV8P2MRDfGw+B7NokPGS9RGf9LvPkVq3Ftsc0ADD6Q
cnJVG8SGtOHs6SzNunFWhe7qOEpZqnqcroeIjdrlXZUtOnrzTI/L7uSwIResDSVb
Zi0a5IaEJ1jG2y7SUubfNGoYbFXYle/m8mMI4Yn8zaxe54mC91JE6EqsNUZX4CPF
1+gBhIEdqxMTxFEu/cVRj/OTrOkXV+x9DxLYY6uOdOiUCYXMJYLXTLNLS5z/bxTi
wVnBV8Hi5V9KErtIEa6nQouWEB29iFabEUiWAwygUG3c7XwJQkuC3my3tjTBJS2+
Ip2CZRCGp3c8mhVJ4HpOQXWb+28RPI+PwdAcZeIm6Mn3scdyovv54vNzrA6SRcN6
5WsDIhYO7Q18DwGHSgsm6LyDH2sK8zF5LzeAJu96iun3yF0wzWBzgpUWyE5RWvWC
bSevJWgXmoVAhuEb0NlPkC1Wd0842PP78QCgXvuoFOtfzrUalUxrkeV57tlvM5cM
4IbkGkwEHvtYDTllfjbAgWgFOQesGAjEAes8jLDqdFicBYPpigib792wLE5+/gfu
e1wrxWvfNT0hPAc+oxug3bPyL5oxK6ayj6m74aL0wDjVRJe+EZBfq9XhxO2yESVC
19UDqUxETejLCAoaM++1/UKQmoBQ+gyIN86lRhd1yWy0kjOYEd81sAZJM2PNFKYN
vzxpcv1s9SDu1wTkkZfq3/vOccPly2bA51mtedMECy9pTqYwlUM4cUgbdZKbU5GA
JgQjmvicQ7Tj5PwxObVVREPxzxADilMus6iJb1WwrnhvPxWJSqWz9DqCbLJJkCZC
Xb5sKOO3fW9wZvw5AMTo27YZh7UcU3zFrQnfgriwBppvEm4Rt0r2wn6RHsHODOWJ
jrzzZO1lcOnxvB7xrmzqd5M/SOWP4yuoOndUBUT6YgvnhwqPZtVPEM0r10ZI09cm
yidvCxvNF72CeKy7NZACy1yWs/vSmMzF0vHJ7YcH2RbwYQih/WBpl2iVa7usQFyK
1SLwE2lx+xUU7GND9pnyghpv2spdKeEIgEXgzl/T2n69eBQOLutdmG1Fl+9IFcLs
bO2H2t4+FxhaD+g+Qxpx/Ukv5YDmSWSJoy5JdK0nZ7Wt01YSZzvCUnC90G4xg5mQ
kpPaEtA7TnZF8keCm7e43zZCYptLSyfTDiIHZXPMx+p8pcGGOJcuUttes72bKRko
01q496ARzjf2vtMrZnH6Fjx6Rw7jWoVafohv2bLWai/WBKLT86ZKZHXjV3xANAzj
jeZMel1kan/pB/tH6gQY/PuaI48WTxN+uvKQmZuzIbfSPjnPiplhkyWVC21LRdCB
DGA8ZNUuybWJNWKOzYkGju9fdOAVvK4KIpgRPY187uBvzYSCJSWHiEgesIiv22iF
maGxEY5m7lh7z6/MaE4X/TheQuyuS1vEGScauknKhSjMU/4FoAl1QjKamc/oiZJO
bHPSZ6d29fhMEe4Ddrh4Og8av+jm4jLcqGb59SFkET5G+iXIPtTgFq0/VlMmJ8Qg
Q35ka3JucfZ6PtvigS1K6txgoybTQ8hp1MaGJ8+Xsb3Cjs2Lgy0jUxdRWLGUb2Ta
dTtgKXbZk6C56cz2M1MCe6oJ4frVB4x3mjNg3UVws6052ZjCpQbrURCORtKTGvd1
9RXMPmHuczax+zlbllxX96iXxRFCxJlRs1waWgfkFfntopElFdzeBnd8s0UA8+OG
P9/4AlY7XoeQqMWfPZZXY/W9RuDiHFvSmumDMs9MjOHAtDIlAZAo0nS0juytGa7E
1BbQ7kYmh165qE3jeYdpGjT/VMmPEx37d/O1cK+XkY5dWOCakHhsSbgBM5UdoNzU
nBThB2gmSwz76I9XNox2PonshuHuNupnVSVmeV1moUqNsRJt9nTCtq90MIfqRnBc
CjARMdA6ZjQ7NTCznYAsQwRBo6PUnlJES5zsFSOWPwB5qRY3zgcQFaRXJG63O0dW
tqutd6eH4A+hSLwaUbmRPZ4xfxaxfHTux33DUYzwHGOKyGEoLWQREbBeDMQD4rru
hk6SlLu5LkpkaK9v0wYA23HVMyr6M4WKjvjvEZPfqZdvUhvWX7Crbn6iTjrBAl0Q
RRC875k1pddXQ5z8gNYNNHYHcwmiwF5wfpKVFDCB66xu6n2UcDdw19DQK9uk+uDY
tvvRQ4qsnSTx0ZNuJ+G9Sy+8MkOpPhofxAWk0kzBITlvyWIc1XujY+VxSfvrb65e
vv8OYHeafMUursA/O2PMTLbCQc3WCvQi8lZtNzn/Et+KZmnFand4gRY20v22kmRl
TYTeaMPxUY1qvNX+/He1/j4LZwvzGObL90C7xxKaOu/3xCnX5G54p/kMD9NYKI2d
FmMIGLgpvZBfETRL/tlxNP5ZT+aEpR8PnsvEriLnH6mNuQV3h3pNsjvFAkyo6Frk
Sjcid2vN3K7khsgWQJOalQXJfE9ArzZuQeinxK0r2dWUdeLcJk8sJlfG+MQJvpMA
4rRmn+VsZ53YzLXdllqtZHUEteQtNj0HrUdnq9fKKTL+1mT8YfFj9MN6gNqI5GJ2
cUxuC7a+6UjGOWKkbcN3y0wmEn2BduwupDIy978zHjPbzQeA1JjuRkYiS0sPgtFG
kNrllTQM9wM8qKUxFoq7j02oWrlyKCMsVrEI8FrCMre76SlStLecuVbE5smSWoe1
H7D/wz8hOoyEKkqYnlYA1ilusAUke5NxBdu9C0ma67Nep781TN77RYpYbF0fDYyQ
LG7+Ci9Zied1/eF8Gy3W8bJ0TzQAyexI7D6IUxP//OvLDT0IbF93J/d2PtEsIreV
NEKDkQ48oBtmzqA6zEUT58UwVO5KLNHbVc7gvN8C2TFPBFFyVz+ECRpZ5RfhnBRC
CYiDyEeDWvffwrz5aUhi4Apg1lj9t1PGtLUbLW5trELXbvluzqJGTYwclAChctRQ
eyBEkAyMzcaeL0e3vjJequWlY2pSTBUcrA8sk/0TQN/VLTP42X/AxzwYkKL5EVQL
hj66UJzESjpv1I7RE82nnBMcosY1tJINbB9nraZlQG3PGngv/N0kblER9ZcfCEUQ
Bbz/oDXcpBKBYxMc2fRAGADJBkDrgL6q1/W9ka/wDq1oG/uT9sdN376bwrotQmnO
K7pRtVZag4Gux7JKUKIggkI2bhQjpB+hEDhs49MZZDsHIinTl49opZ/JOSE1QIga
gk5HJubvaAwGnvV9IcPUrSSR60S/hzzjdbCT0JGgmt3gNCpHHT2DiMqYSaFMiKGP
FykSUsRghQ2HXYs5QVaLk7UhkRRIb9W2HuVn72/6PAPYUk0jCbwnQ5xStrkx+hWj
kiWtaWRTm3nuusEfOSWBU9FSJYFXafceBpVBTz85SmEJxH0cpkJ6x19hyUyJuMbO
Qu5zsv2vsmO0OULXCam8ikLfzVGnfBWHESbcJLfpEeOhENv0wBJ8/ntbRdADWXId
4JnIlFkOhDjCHHcNjnDLFr9GM9ahpbo14SuQtI0nM90bgms4tIxq01KxVD7OQ6eN
sKFk5GvMif96xzzsOO9rNS2F5RlJS2mxaQvvvba295T6VM4Ud0rVFULhzAhl3VHQ
EZL7ZSyo4fySFYGAvJsWK44T9Fz/136NvpccOrtSygpmp+86x8Wlo/oc7XmYGYPO
I5BN60laK+WN1ufdlh0J9VCkjqwnDl6npss5uFNh5o6O90hHHnHmpe5CJTfUGwa1
O2QJw45EkJG8XYY/tcNwuu2EjNsNq6cbbpEeHQXl5nrJpRtcurOEr9zhXp4M+7kQ
mlKWJMnzYu47OiyU0LxjXJGS1l8DDQKVlQ5sR1Ez0PZz4vRWJjBdBWesjCClQDoZ
qa2Kz+OjFYgF7kXHsUtmhVVEaXQakJzY6XKeAfuQ63IZ61TTzRzkdzwf+ld+FR24
XAKT3jJFE6qfrj5/NPGMoIsojgH9ZaqbLRRDRekWpU8xiyTZ9RVkjQo0ew7LrZt3
hHqrVEtfBcv0r5J5rqUn8sGSrokNXBMIhLIHSRZsIjfzvKgTWOUB25uMMTSwehe2
gniyKzIyx+d6lnEED647IKga2523bJ4EXJaUSCGtyJUBSgBxbfNRn6r2ozcDYZY+
q2BZf5kclhV7dNrOPAocWHQnz6AVwIIHF3LLK9e0CBBD/e4VnRQn9Af+vUG8DTzL
UfAbGHPLgavG5vTfSqpMpgD/vbJ/ZJMUB5hczR2+5SUj5MeSecFaiJbzp5/DjBv+
zVUP31y8pSHpzXqhsGLkfMBNA+8eIaeDWbF2QzNl1c4OyVSwEmWh7w6HsOtO2fEA
9RgcnSvS4Zqq7TjdMdbUilFqCjCe0QMh2nE8x0wp4k1KgfwjkJtyziywDHTyEduS
5GhW0OF7WwfVm3L4Vd8D3vVubQTJXQvnd8QKKR+q/adUCEJ+NtxLz2ehb57DjWWM
uCAaQ9rqe1wKRGkPOClh2U4T1PFwtcX7IDrlaSD/aXLUuxsWim7rKqkkIxGCxwcX
LsTkRw3VzHG9hAq4TQQJDi1HzIDywTWj7r27Alci6SNXqH608sM+festSxgGekfg
U5BDQ6rKz4r92/dX4KpQDPTKgVx5Q0vMtF3MiTX6dMGsxHns2aPOS7h96MJOudxE
tFj8MOM9cSNHwFpUh20z1XyRZWsw5nQo06jMpXdcFPvkiCCXQhXrlWjOWiZvClDm
6ZRRNwx81kZbrSlfnRaHXo167MHSu5AgAhoqwsYWZV1DbSDS9exx3m0vWtMUABiS
eAj+IsX2+HutQhNGGajmnJhi4qneE3aO2mTDKbkPeycbrneM0z9bwUAEg6DvkkPy
y3WLNcIsBorBC4U56VC7TVVdV3s7JO2EoBDKo/H+IfjAH8MbfcYL8NuQn2F2+UL+
UA48+Mdd1NECVo49U1nNSNL4rQ5yUQEuO5rhBAysy89EzmPm4lEHEXImbqLlMba+
A8Wy4XS9Tse+pkYezhFNJMShZOZpn+JZlk/htVwJNjUBj2V/TG7CYwV/If1kVPFl
EsxhvOZ3h4HKAoBsvFfNnAaWliNU1wNIfgSVSHSGAYtjNofpf5JSScTtcEX6FvKw
GTK3YiBQV/OUOYfqiHQ5vDDDuUsfABkSZS/F/XP+eBrDlZE0XDLzAbz7AzvbrWbY
dbee2E7jbkMBvap/mMs6QvTqINlgXUg2eASl2NY2Lj0jmUD9cjl9V60H2NfLMG8y
4M/i/nJiyAvCky5Q8A7buRo9CGlwIFMOochPN/ZnhB+moNNIn/a2q4KwcB6ZCX1S
3FNIgoN7/CvfvtOoJ0Onb+vJPNSfCr/5Iks+6tAvd47VeMBOEiYnHK2X0JcokImK
Ba0J2qItKwbVoL/TTzJEME+YzhYwsQglhMH0QkDwkbg1iK5jHC/M1x22liPh1F91
c/iAukh48YZ/9kHOOZ++iE1mv8cbKMhKPfMKWtlJSmvKcm0IPz5HX1ZBwdw4vc0D
AJzz53fEzeV4cUUNSggjWtG1Z1qAWXmC70bJY3OKNDjuheyn12RFXYgVboCNkj9F
ecmuA4hquicD0T9es2QT6B6qnhRO+EgzxXE3JLKvUfmdGgPAJI/R1Fns9Rd1qm4W
sM2x5/06RH7tcaa9JdxjXswPaGtZ1C9SHAq8YFjEXJc1S3b8NGDrcHkMrvx599W/
fV266ToiaHxlUvEWtZbRUd01f2IEDCUa838n7sDLwWJFifw1eebJaXu8/AuUZv6k
JRJm125bK5OUsNTECb484QnBeHs3v3/UzO6BTuH+2C22HKaNe3e82gVRJLgQf/Mb
PyKw5WAcK7RfD2L679Mkcigh74+sNGZm0dvbdLYQ+zxkrzgCMhgK0ACbFNKnf8Df
CUPutLJbOw8pYzL/vzYoceQyEMWQXVK1KvDwmgoKnU6KOBoQqAfKRY+neB+RrxYT
76UgveeMATOo26Ev430UYnihvx3LMzrg+8ErSyAjLJmBDwC6HYphME5ePDoMuCmm
ThE1/FAgiZJkq2zKlqQ54xruCXpDqezis3OmGLVaejeNxIe1TzbqHHFYgXu+NWp3
LEV8QTvqiFT0OlsgcBcHKTnUAOKWLwCBYNpYUN7oJM/mTdF6PcCfmLjJICPSmnrn
qLoTuwXOuZiHMEZdJhJgw9gh/xwG//aEOfTWTWfOaEqSsSTuGgX8CO4Go5ZVLqwM
/aGO/ODQLrdMw7G17nmfm8gM06f7yqZxt/P35IDLkdvnczsxB55uTdoJl/B0WaZV
UC76RLQa2jEueXQ/InxE8RnXyQtVopZx+ArD178W3ayZmvfPGDpUedNci9Lhycxw
3/9hrN8y2FVacsvKtjvja4uMXP5d3nzsEt7ukibiOTCiQhsjohTf3np0VQ64RVRi
hBMzewl1gYnbYGl+usOooeVBgn0j/oS94zMgFqwlK9nFEhP1cMaEdIBLPUMg6YPo
ha+0KRiie0f+5aR+zRu0BSRImJIlFiLZng+sRZ31d2kiFJ7+zAxXQbQGXllLF+gc
qVYDFJQq/F1iMNL9O1tGAxvc3xnfvdoToEj6YLcH+1o9SJMFZ9xqwjjD3n5gGsrA
WZ9l1iGgunujOvMWlF/3jIm+93p2tiumC/JonslX0ah4bIYjHzAmGoq5il32gPl/
cj+LsNERWi9OFH/MA4gul9WYtS+ayT2esfNyQxHCxgKAHzjktsxIo/X6koGnI+Cn
Evm/bPg7SYA4pDdLcr3SGv8AuShxcyBz0MCqiClHqZpjz9xr1o8yf9LVio6X5bA4
Nk6OB0lj7gNsZajvNvSuHmp8771GH9TlTVaBqnQ/ZhWlWBy7gt8S1pegtfmvgnu/
xUCy5FnrTCU1BMe+erEdm1QYhkggvEAr0Lbzlo/MOIzeiVGwsjfy5D4JilvS7ckL
OHitH35+NaSywrtIzrfJC42xWbfKau2aPp+O4th/O14Ad2TYFTOhWib/i8eYSIQH
xY8LpobpJ1ue9KFnHhYjQIn6S2fykcOWLq+B4/Lrj+yNbCZLGMhjgev4Sbrk3bs7
+gFcTn13zwaBy/xUZpH0++f2h4DajHdPQFKURanzcws7ZzP4eiDqdfh5GG9kMEdq
7d8ravAcEpbv4ie8FXlXup925SmtLFGLM/4OFbLQ67Mytq53zyU+P/vdTL6/F1PS
+3Qof7T2U5Z/NbrOmnKlPgiQ5Z6NAQBsdGNlRtfM3PC6X94zUNODuJBBGr74F8ox
8WnPtWNm2+IfuImRzDogM3kW9kUF8SlADn30egb3Q5Qm5tKFwsY1gi1KXFd5TSHH
/MXuNkNhq7qbKPJ+BywAmOggDN4dZCTBBLUxKiqE3NKzGhDJYfp3IZC/grau8g03
mjmOxMSVk0NPc8Y/MsVNTGfOmxDKgkhH1nK8fz56GWfRR/6IHHWgmdgwchUMVPQf
YRCT0RobV09bMa2kQbZP7Ez9JlJQWHDI/rHX13gozyNqiThf81M9maWGvuaZopy3
D7IbCoFaiwfPTcoHfNyRU+i2v8mQ1ug/q1Vkj8HH5nrkfVylixMz0iEzXXFLBlhK
4W6t189JPs68+RA1hfq+XQT615vgfJ50EN6ZEfN381+bV+ByJkujMyTfkqSaq8r2
HG1y/Lb+0Id1p3UMDiWWnRYHC6ME3V1IbnMwmYtoUjxgusePT9QIXTkJvpVJb5yw
Whx8JqiuQyBcQLoFBkwTuA3Q3aW0olJv76mdCNzZBtz0eEkIGv+Z+l8ly3HnKYg5
/AZ8Pm23niFffxh5130B1Pi44irA5H7EzjW+SYNaUM/4H0YEe1bWiGHpUsvzmh1D
yUB1t7qqtMnv9ae8+00DgjLCWECbvYjx32GnNT2fP9jG0eXaU8TgxO8VN4oaY2pw
C7Uduc+AMS4NwjArCkuhnM1pgxVJzbRfJXRT+UpDgvzunFDjZzn4IYJ0f0pFjrZS
PE/UubfxUKH4bTZoF8PWUxddOiSylhayN670vHR8m4ciIuzrB2Z0R0eEC67anuPR
hGlgog0AhxOhJi4WyimX5kb+b3iitKOxn2RzbaCmhv7bmyMj3vVe0Xod9cqO63In
9+RWAGrsQka04qnsGgzryQgo7PMhYuD89w8/L2K9p23hNaFSutjelI/y2ekLBf52
wFZtrVvEgIFlcmP9mnWAWUZNyVo4iWDnXgPR6FH9jrQ1ehg/FtEkGwBAme9bHs9l
DwseIsKe62FKngnDV1oflsntvohO14sapWA8uW5TUh/RydE4arNILWDVUOkMYvse
QsIxIpZuKI8zLAUrfRQqNJ8YUczjdoQgMFJ3FnwVmwlgKRf4E0csMc3UXl0Ifyqf
f9/hNlTbSnjSK0XuHSljWoribsxBiFifdKRfTmmGPEVMTRrOePtX/jvrV+rjcYpa
IYE/iNKVRlLzEqY3GNypq1hLb5qImlpWkp+NKDJWud3zBa9FxKZf5thLOzT7i2vI
4mxx6sX4yDcq3Wo1G3UqwPe5BNqRTs++/SztBTxd/nTir/6IMYl+apYEhY2eqlFZ
QwHFhwmhhJKOMbWaYr0ZnpGkqUkgI24zYFpWMHMbeJsBZ2z15Hbvm01ppJHi4SGZ
KCQQd8db2aF59QqrgQOuhTfIk+espCggICxB5A5N+kI0fOdXJtrrGCExzm/9PQy2
PB4CLbqdoOajyi41PyNrfeGsazeHPAlqHPuThC6Kv+nlVY0ejrMCXljL5cbLzzK1
pzpGBmmDI+b4tZBrdlFDmrBSS7xAvwhsWfOXm6nUD4zGMi5dKWXsgzeA0+kBL1fG
RJs5iJz77E6r/p+JoE01mIimo7S2zidAMPVGwcY7hXJEQBGVoV/B72U33UTTPEYi
mEGSuO0JTVRS7TmCY6y3Mr2OY54fMpSeb+C6j4C93fn5bQ7uXk0o1ZDB7c/kZnpF
PNp9Ps+68U6y6nW8rz0BfyWoqX8fP6zoehDVyF0OuA8fj99Ry9FQCgoAVNSJkX+e
nqcrLXR2Qqy/o5v/1p8oCaHynEwKyJmHDXAX4LdDn3Mjj+mweok7l5I18cZbHGxM
81h5J1G2D3OfY3TyQV1zRK1UyRBZQiqQJ3YQwTeStdvpNrx0pdoyampLwyDP32qP
bUyEJLSnefC7GaEpzA8/Ej5jAXAtRGCac/VBFZqUy8tzm9Zw3rYPza/qlkBsdigj
WKPKlCt7zbdgVSscmzBXI5dxHqQ9ZV2fY1HptJRSlmVYq3ya0eujCSrWmO5KTXfA
Rfq/PqiUBvU8G7YXdN6jmcBP5C8QsXRiP00RMRJNuQm/aTP05TJH5t2eXqfmJbEN
zcZux+MNMXzMV0tiNkGrGuhrZ9hdCSOdusmkT86FaUirgdDJVuXsztvwISUdD6KR
S8ccJFwynJBoXH1EMWOub0OXVY4sW6wQwhxyA+8MdO/wRvAq2Yb84NWdfyY2RZDP
n/xZbZPXj3vzwfPDIAzgooI+4oSp0qALWK7BZB4Hzl4V6poUO7egqLYhhxMSmOTA
2ySFBVABJX4JgAhf0AfyaK58YPct4zvE3z4c5thGLh2v9WEX6cS3xANc/1hI2oQi
XUdrkcVx8QGwRE06Z72geXGiKNAh+tWutNwtiRPDrDVf7dYLPR8I+PfRkd1QePfZ
SqpsK4ThhSjmpQoSLc5uM2C/2Iu2nCnQJ3a/E2gF1JNx07n9Dh0Zx0k4CRkMHUBO
rxkL5/AP5hc11PSGNV1Ak4UxF/MrPj6b82XHw1yxxEdIJj8D0W5ffqlVhTM0XrsV
oh5NNDJY3grk6lrqpDoS00kt4vSPqW87avN1YiL74nyOah2SI1i08v17FfA19icA
No9jI4Hy3ROQRU7+Gw0zUSMplNIgocIJd1npzy+PZETXi/DafNPF0G64Gr0vjSLG
ojkc697YYesi3K+SafZbzayGzMXoEmY+IhN4J5qCJOct/uxFsU1MJ4sZUwGPg40l
4ZOXTcvNNtGkbOQtfcXtC8/5S02o8gJTQr9mNdbURxn77bSYjli5LOMJ3pRuYMTH
yaXO/BbGctjJbxFurW/fY1gufxzxQBqbuMwt+Kq6hV+yqRyNoNkRYWAYnhK0CjSM
4Goe6pZF1p7pmEJZz7SPY3Jri9lzyZ1YsyCkZ+/h/UwTa7R9JPmNgxgSFVvp3gCh
lR1E3j5sszxD7SAvaVKC3pirR3AwSRM8v1lP+cqkmXL7Iv88wI/AgwF3qVumgHBH
61ubUSbwDXO2DUlIkyQ0LO2ADa84vrYD+eK+0ejhgpZJMXuKD9M02Sm8t7ISUiKl
CUA2BqAy+LmC4EAgZjPkqasbrJgCFWY4njcoxg7enBnIgmdJrFPN6YYh+T1hfir/
uQ4Vzfht4jPhrEFEA+FtssAqPwKULNSXFFGBzhCP7LsL7H3obKCmIoiswBOMRQGl
1RRwf/z1D4eKvcKaF4zIcOOJIh7uoEKj16E2mVfdBKbg7Xry5v8fdV4rZyIaTih7
Ius8s42Ht8m78Vo54AmlyNvvkRYbMYPjt2PsCNOVICoX8YE8FWlTdvcsuV/nwSEF
7+n7jSUGzhzyCo4mZd7zL+MSSW1IBhAFjtfHiQ5O5STokeywVF5/aw7XI4Vn2wYC
bh2dtAWSE7dSw7qfzSJnLhLXfiMhgSR6rGAA6/O/qlOGrUiv799N3yIKfcwfVLBe
+2RZlDXsKy0CeG9xttO9xYzMkQQWXsV1gDZX+LNcYn4yJBO4SQT+Rl+/cT0SiYs8
tcCSJsiT7ADshXspWdSSswPIxBCVRHsI46PjuPtcFH7+v45p43DI1k/SDQunF5tJ
kTJpnoeukiSpmXJro3LCzmW9Tjkggu8t+X6CVss4PrDUiOp59n1xBVLsdxKRiCo1
NjYwTXZ3KUee1PxW3EGuRYjJdfCej+T71rokopB2dM9ariLrHdzuKdaOBAlpN9dz
vgutca2CV20zoP7k5ojVBUs3SUU0igiHJINmcEuvHFHydJix3C8daSIhLwgq0X6c
m1hvGelQ+YS6WSBVwsstTaT+Jz34OcePcOrkDueXS7N9R0OMS5sm/vfcIdOC/Ave
I1hNY66Epzvseo/oZZEFW9bjHpb1ACp9GrXZzN46KI7cApvNfaSl3F1seB7pbVOS
XkMMMWGu2E6fn4P3fB3MCh5r4Q9I/iJrywe/IZEl/Mz3+mLPdBrkeabqKOmcEcyr
tBOwfGzd0ZVUWWA9IEOfmcXT5ZRTgiI1DM+hnS35jAExLRGvkUVYEDJwev36M54Z
up/ZdOtCPSgnL15xesYMJFVWyLHyI/NrT+i/g//OLv95yTEehwec0u2QBvYciO//
bmHetaEB0FuSL2yZ7xaADF8GGweLlXos/iuuYpMZOLYHbyHYCh9ZWAhb/XEnQb4b
V0xm0C9+Xol9sfxuYtcLQ5QBXZTVv+Z4ZoF4cekHlBc+T7qu/kZ+tPKn3ILuej48
9REg1DhiT+b9KV//FrQ7gJmx4pJAD1YOtAXbr39H9BinhRlOQbS+em6BZGtkUdTB
96t5Gs5p+2WQoyfFZMIE7kZ2EVOIWHVnHrXxP4W4rOiO9EGQKuxrcy2TNZioO/RM
Cqly8WUc+5/z/tcASXuMFMr/Zk5xjgJQoFYWkULiBlIuiZ20JEHzW5y5mDf3LXYh
xBFoVjmrN2UtSU7PanPhcHOFGYd8gkOcI4EWI0+ND67b8XEvPntKh/YL5JXorXSv
sAL3KmJG8qdxVWQriBy00jcMM0itXkALvhxIuKqCvjIiePZdov0ozl4epYAMjJkN
uzjLUgYLtL99NThOkH7FdmMAvKKhdhQ6dIiWUhxZS5eNuwbsDRWFcueOhBI7R+WD
kWQC96R/whVYFJcazuCM6hPmL+JXAsqsxnaQuNU9Jwoy/wIgpM6GKQP5fTr8cUjp
QF2gyTH5mT1djkBD08zz00TCRFiGy8ocwFwcr/kxkYhBQran87LbRndg4T8iZsP+
6iOdSnQImqw0U8NQatUN6/3FnomeXz0Gvt1wRFjBIV4KN4fDOIm6oBsQ0VGzsay/
5qcj9PLw3EjebtsE/l3H4lSgqlz7QoVfXI8pdfIQTz4ZTdKzxqh0YjlVL1aOtQKL
`protect end_protected