`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sJVlH+palpt42Vz8KbH9lXglwnvVIZm+k56kVhW5D7ljlb4zmnrHkYEcR03NrAbN
/3Mo8ip7mdOA5lVIczGAy2VQJCsS0I1tkOIu3/i0v6eFINnjQMsTtIBrebf3vEwe
qyNO9tSdEgFPZuXeeukdSDSYlBWN2HRPtEY3jZwhT5MFnDqocnrpwLtCWGHfhVUN
geF75buApGxyvm8+vCJmXSDIbhYsqzrYVDR+NaQ9/m4M4dIEyq3yyPfygXe094AC
jm31GmUAQ4ynp32nFNEFU+0JaPvUF3JeTvQuuk4SECbG2K94DF9E30aH8lRAig9+
9A34C6ax1YI1T0/ZSgvVHkxpx9ExmeGNuQy4lWbJdKWph4FaDiT4fyKhp5U9Lp25
/cL7MM2A7Kp13iJLYOjB4W0msE6nMn5IkNSqdRyQVEbedsjBmPoNx8DnCPcTrkjY
u9XaI/z+dE2SrrBc7uEgVDTvvFaKG7cq7aCnXgaVPHCd4+P6RGaRnnaHNbP/lGYn
RaIcrJqJ4aBBi5z6q6mb03m13ugYMZUyD+6D+N51k1TxlDvMUlZ3KUOQjl+GYCh9
VN5gMhckTFT4aDCikJ10vLMjBHIlfYFbKIj6H38KsdVo91WWG6MKHITnVSVTSRK5
GClsHFhu3SRsiiKn1TAYG01ZnHonQe4T4LXe2fFZhuaNauTVyzHva90GfStzLwNW
x8ZnMoV1WN76Kb8MbGtYyxRpHeuH5SIEqntGqbmeHhN0AmeOH+tov1qWjvKXdWeb
P+ARV529+H75AKeJel+n/6KoHJ05z8WqA0N4ND5uvlB5Jha6PSK4tkSEeXKqSwFJ
I2XWBMLDX3CsFTncUpQUW+hN7MjyR+XJFWU/NBIrYhat+2vpH5qX4YueRhcRmUTV
Dv5m8/Ne2F5fUFpZhYQstdXag9LUuVAWZaL8RPPcEZFacn6F3m8hYNlmtwP15Q31
nYKAqNGQVxysfrwOnasiVoCQEkXEuE73uwG0QsIyEw5JD7XrwSMYlBC/EyvuxVFM
0YrsDzvf7RJAi1JmO23h7rpalhWaVBXWrokVr1CQ/3ASLjTXdW6ns/Xq5x7PrxBf
HqdMp9meZvubZa8Egnky20lROmdVnbSg3uniUQtNK2zn0QyvZqHbtAQXnF1C0QO7
76VIQ3EndmLVusqCv4hhx6ymLM7d/FNin1XTjU5fnuYLIu1MOnAro3iNq32h6nBg
nmn5nzWgmjTe5R4WFCmrIoCq19VUIznvBVw+DqkDRtxXlHB/0msBFjLmxgbQGjg9
1fiLKcQT6Jl4Gd7Sh/PIyXF9fKGBskZv7nL7CCdbI90cE04Vcgfs+l0Gi7VO79dc
3CEYWcEsYdbFSdpnu6q4Ajd6DAlBjhOKHW5Llq2vpwIQyaGmj6hCSYhk0uXlP2ou
gmpyHSdvl44VMPbYT3I1S49Gdd1tX1atekVdeL5kHa0eTUb0hRfIHH7eOqZZWh63
SLtGAMAh87liYrvPMp9NibxXby6XZPwpFQzPVIF7EvIhcEUuNN6ktEzbcDQgICHX
bSuJ1hKV027m6hUR+y1VGivwPn4Or/bo/qrZHnHKlg6mo7+laQIYDNZTwmJ7bQCx
vJHrnDKpRcrbwnT4HJ1G0HrpWoG9Vd/hdPXICjCiigWQgsf/JwNDswLPDNjyNdrz
kSXsjGBk3slTNP0ORwp2Y+RtB7C59ZOuv1f7TDxlRokcK/W6QiSdw/7ZYREwvdA5
5LTcIoyDiCjYefNp8D5dsb+0/pMOLwzWDttmEOwMx6GT8ZfZDx5vDisAcHyiSHBc
Y0pAVqKtT6QGvuOruxHBGlFcy2ghofhCgXXvKNiVNqfrM4VDOPiZwz0pkvoFErrn
N0DivUmyW7in114tHFan6cfu8mRBSx+pmz9RsQdCSwHXxwG9vIxkvVbHR33lclpn
zfk0XzSXulSfn4khCylKePrpbBF+fM+Kcs/1THWkDmKoScDKohpr88bNr7iliBtU
4PZWKXDn/ilIcVLLmUVfwDedgPByFFAuTrZ3HozD27k/9WLAI4UEs4GgRjjhEcJi
FOdcCVwu6JJiMBvtNP7/NLvDMuhiaIbKNFpFzRgPUN7B7ng/KRsqu4+RNIx3EQo9
/Ft8OnGAaS4+HHTaNAwf8StAcZbHrdXgp8gsMSak+bB2L9CcrmTYQDyq/PeJ6bLW
q8rCQFYoko7QRHOWQehY1nVZEjKmD8c7QJI+Zqi3fszmt5CYWrVH0Blc/BleNKRM
EESK29RFhgKJUzAJEknXgMGiHsKAmzWbSUOMHCANaV4KCC6XM2QxSkSmao8fIC94
dmSrUTtqfmFry0WeO1AmAlwe9g3pFGJ0Pav4pGxNkm+bmMeBBnyZ3+0vNq90TxaW
fut1pRPii15Rmg8zNTHhhzcFgdbo+vV4b0K9KVLf/CtIRLXF0TmvfIb+H2UGShx2
zAQpnv5BEys6LlQgWNDhW4gY14pHmZIj2eGJdGl8oIugF0324BqIziDG7CXqDyVb
TlmezcjswEfe3yveRFL89NjIAIB4HdF7hcy/CAcnfOJiQUdVMe2X+pOmoTDHcV/8
wpcBbkyr4VpJ7Bm7fajHKRtuILBS2JhhkKgXd1xRhTMIQmScpAP6YvZazFHbSFJn
/D3kZXO7/WULAH1wTLSIB0uqu8xyz9v6rU9/Y7l4y+YeZLKgIpFX1WMeeq5hZxhI
e0iqLUPoZjFBLK6lX5Q9VVpAbD6Db9rPUi3UL4e6DhfImKp/sk8C/78+ov6W+893
wSdaFniiDseyyu/M0vIoDQFEQT5Iox+mYsqBO9wEM+kO9M+p4fupmcYbjZJJlUFE
WaCYra79Ptc32P3thnqdxDNCX7LR48uie4O04qg8JcBSIqqIT9e5yB6pLzoxsZT2
836Dgvvi/dKlJBAJCebhRNp7Ob5WKXwgluMucmauKmPNLmyXc5BnwmFyYvIZ4bnD
HWlYqfgedjugjJD7WSEFvprEY/XNPl0jlNTFN5kM4aY5Rjx5nendIc880yIROgfp
HoAhuQvrZZLzuHdHLC1UyBW3+aoKDAKDHHo8fFWZzcrThy2jWv7+e8YtPvblBQUF
GvMcjWrLXG5Fyu9CJrr64dtjVCseBGnFaE3/gM6pgsX2mgtdmNodST2tDfKj+Zmi
FjlOgAkH75lv9ck+jcY6p/rZWA1+SC8630/qSe5TSmEDivwIncJJUbrz4uWBBCdg
h3jOI9lfZA+B6lohnyAqeawe8/nbH73b2s3M1PA5+ZiSGv0YxbXVU2UM1CSjD7pr
VbGRqNe8M0sJc/36ymvB1h4/SN+whHKCr8maNyogr1/psgM5PLGscpmfydwtYL7/
w4WnRXr2Dg3lLLaOZV8t+VIIb/TuljFaXb365ynXLkPUTYvwo47Ylr7PTCQbHht/
2w99N+NDh3SXXcC//AGCD/l5N3WaLXCdiqcJf5AuwhqDD0ziFIWnJ9pFzN6Q87W6
L3/uYEvS3hZaCyaHxDt4h1B0Xbu+lLT9hydjHFI3TS9Urf+RbVuJ17w8lg2vuJjR
HEL+ve5e6gi+WpsKB3beJl2dcDuVPLbv/rEZWHP9LaLm3vhZ6d2dYH5pK+LOdxlN
nBW/0Kt7ZTnDyJ1XEPm8Kf5/+g74k4vkNfGwNpOX/rXN+2GVdNgnWo5AGC2jiEt6
9N1rWN6dHK5v80aG3STB64Cr1KKBAlBz4HaLkjLi/tNDIuNMyjXWHVwOEQQR5MeQ
fVjPUZ++yas3lcO36MGIVqp1LcioKSsCPhO4grrSaFhOs9iudgcCk+s6RpQ/4x6N
B4Ak1g1CBC4zd82nbBONB4rekYzlq7myWPgnHO5kQkxtIATtwHfKq8OKqDqRSvPB
Ywc/zhf4t984cIWdjan+iWs1xZ85/YAw3KaYaqME9RUZFM3q90q++bNZaBUhbPaa
aCg5upvJjRjrOqH5vOCc+ZZl5GQJorVQP3UEOgw9BUawE52bKH4Os2qPtcQ5t5s6
cnYBRMBBqdDWbYvsqJ9UPsffGy9KRJrr6exi/4H7dMfj551XTkA1a5GLxAbL7c/q
xV+tyNWJbN8oxecM0PxqaeJ6MvGABSon17qAp/u4kfGUCZpSLaME/JjIbEjy3RUx
XPKCi3K1GmZ0UvrVNisdx+8VFKkyb1GZ1jd7OfoD14nVVSCzUwY5q/EB1r7G3zfD
HLz9Np8XKrwsZbajD0by0R+4gFXwCw3fAQStyeq2nS+GM5BamNooJaPsavvciurH
Qo/A3fpgh/mpxwlnPIFnKd+/0gV9zZjJM5Fentlf6N8gOdSZ16fViWivfTJ3UUGY
aIdYQl+xLBEv1mzqc/d1j+LKiwJhDb1KF/kLkFo2th01y01+ZVm3v2tD4GkZgZfC
P5Wg5uzzo/AdkD7RcOKnrbIrmc05RKyQUfTVMMeBNRi7v9ER3bRqjbreQ+gnl9B8
qjj0VGDIa1ZLHp377TgUXu5jnZa39gpZgV8/0NKu5/4X9MMOC7JmYfXWZfkq/evY
vkeEZYerAm+gnGCX3QiTi5Ck0igCRfeXBQg103qeeMGqdGQly8UhGVCSKIqS6ClI
qU8Of06XSdHBGWcuNZgOk65HXCm5vNNlZ/xJ4XgJ4QUrn3cEopu8t0Xt2vmOOx0P
13DxKg/ye6lGE0gbFQE2pVn4pJWqnu/hpGFLitINFJdWnIYftgzm5jJdlMGBk7Dj
RCdD3d19tidKuN0IyRrZc3oqfRbBPLo61sjvtlSA8k5D6DjEfWmU1Mdvt5Fv1hdt
aLsoqZn1MJyLHvFKsyCtmE1rOOBOq5HCJySh1DuASY/v7B0onO9TlcSjAeCD4xHr
VzPKuSDAHS1zZOn1vzt8q50WFq73p7QAnkD5tF1dC6oAufmICyWSDJZnno5A5cuF
TBod1p+IQfK1kDZp882hWzOj8N9FTuQ1xQLUW9NcAPZqQUpQlkvOg2XFbnNfuu7J
xXK3vz103jL42DtM9IsQIBcqxX1Q1rCXoD26eCAGg7ktwrZV+2m96L/1lkkTNFjV
JYTuoWBLvHqi9au8dsKh0xW4u8MN3sOKWQPBd7KE6hCslRoCI6uwXlcudqfayndH
gt44+JaTCGU5gOp+WxkFad1uUJ96ty2B11yxFkhvFe6pAiIrE83L5ST1AY9afOFK
LigGI70YZRkUPUZTCRUplE94BPOMzptXZL3V08FfY1DRNpepGGi4ldQqrTLDCtSv
C16GltfzUy/q7073jJt8XNO9ijmWWs7SNCLiHMBbPJr1rkdSgSn9Lkf+l54LnHhW
j4NAfnjnvTL2HQNwFHKg95znD95QBpe3NSEhjNG7R5beQzI6on0SeCsXxpHWvJao
+S37ZvjU8iH3LCkDTyNjSmo3sBO3zxDMUksTiWoj1xxMIjDGR29GSWx7TFRLuLse
sGgjf0VWVvgkE7Gc2DRWtt4pH/sq4KIRxkNY+/LSScajrDf3aOPbWpxuROceBHZc
jR+VGcv6Xh1K+SttleAznY8WwQoHRvNXaF+/YAgpYmsSnJGLNb9gwm1MfW5YJBZ7
JI0KmgGnxUND9gzQx1sqqMnuVrLdgj6SdFtoJ2GBfZbQi8RbZ3WP2qJy8WuYJJZC
5dIJQE0v7cZSumiKcLSMo3GPYArCyVASYrSwSRoUNVqRyz0j06rtJWHBj3gjknE8
h77eJXGr3gBL1T/8iC331qgP7d3En4GSayaEQ0v57jBDsWwj+K2ducreaPp2/d4R
wOxWsvRcjctDfNaHwhACgWL1DUjeQ6J1VX8kiRFggf+95ldwnqTXWpjuWYdhi6k0
34fZ9X3bf4W7vYONzH5gj7wcQmYGFmwCp/b8XYeI2v9c3obpqLHHVIpxwKnRx5FX
jqV6N6CH9c+Xx5qonnuWYROGrDLjNVbEqzA4FtZtaqb7YnptByUSnpFZuP9PLWa8
lBilb7r588x1Hu262fuDWdfIbliXAvho2XnXsj3rlvqiWoi6RWKQsEHH/XYPqwvI
lU9PID5ia4c6Xy8pVCuIB2L7xwQuXsMU+G8wL9ECjGpDDsyTfaZ+OmtXkZiK+7EX
ieuJZSPBhIh9WxAEavbr8NAOKnKGwpsgKyRuGRY+kjYco3UPcU2nuzc8MHRbWyvr
Rp/l/uKvXsEbIawyD0ywFvdI9KDF6OneLRnTeFsdYHZnOby3XOzBzayEyCvY6/si
PszK5asWSdRhv3DwFoqRvrF4G31Fo33z6Gn90t6PuWoawSarkwlCBY06x5PjHait
UQ4ivfQ5Wabqmg1Q++pnV6TJed7GVMYorhf/rJ8gf1LAelVVlp1qtUKhku34pQ5R
bTfzNBnyqWrDKNA9utzHDnjw41YV5B2cTTtBtMy5B2qP4Lrh6CXo1VcDvKkTdHCr
GNrG1ouIm+oFj0Xrp62+V9s2a6MSmLiJH0rydauJeTFR1O6UDUIsRAMUM1PRG27o
ZeZZYbpMaVErNpAMUEAdOZwa/cn6jOwj+AYbjvv/JVjgFhV47l9ktyGja6kR5jsT
OAra/PauRKauCEGRy06pO8QAoBMcx565QrfbEwLHGR70Lgk8wFTbfV7qcxXT9hRX
hOHRSalU9ctB2s5eCm07Eg9nJAEMbvjeRmKA6Me9gURQu1vt5EcjifbSA0qNlNT/
/eFHxeFs+fjTYTxDwgaIfej54jG3xj8RpC/wQ1GUK3+ktVubVSntx9YZHE1IxXnX
atX+C0cBxBcHDwFeY2F0gs+CdFAhdlOPNobv/8mM9wC8nbEGhZRErWi2u9dyXK0S
cyTLiEs0jlb9IvYNHyloRgDvLZErgkj05J6C7d1Gx9oRd0UOEQWD48szhCdp3m2D
IOF6CRt+i57NnYlcfwYHXUwAtZ2qxFNXbyYbmvoLHR+KKDZlNJM18KmjZs/HIZr0
n4iIn5poqULZJBVrovzdyLQePLjkGLUs41U+fIO5NQzk9qaOvutDmXrp0aoxCnDB
l+LdPdEbZK/hszXY58UnmtD840N0l1q4md185obK/ScKb2PAst/rc/JX1CsQzQPl
eH83+a1trP+xShFicUx8VirGk6pSdeHCu7QCM23Lt+aamFbZYxV/SZhzUVytpXMX
tJy9c8y5Yzvm2uzvOl4frrLe5CT3bRGtIpjzWU/gVw1jOSnAP7QltvdMbVzfyu8S
B+JvvMdT42nltZDkRPeylDftQKVZbnntB8mwDZMQD8wQ+jRx6UmgzuNiadkVWpt6
HDnqG67XjLtlPqleFvrQ5FfcQVQD33WoUl2wfjBSw3yKxGqo4qPwc9IXnAu2fMZD
aBKMubprkAzU+WJ0TAxjHS+jgTcVzxfxJDOVUg5XdL/42ZjW5jFTfefJT4d4SRAh
8Krjiq9hbxGsxQzy6diRnJMCZxCebSrryFghiitZxRc3rZKDkO8kBgK9x7TGQTPc
H6sJJnnBeH4A7pYC1b69TiaIgyPm3iAWIEzBSfjcYuICPdkS5xgVZE6boOsiGosi
6p71YTjQwUPI+rQSS0Wdjz5PX6NBR2L04oXlFqn28StZcu6w6SP1Z5TcFV+PUHLz
LNsruvSaL24du+azTvyIfcqJUcUfMnVbo5BR8H9ZDPK8EYLQ44xeaRLnFq6e41zb
deQl1YDSuftq9v3JBuN5kGm64nMG//lqiPhRX7Nguq8hUPNIYQqCPzg+XsFf99hW
dHN+Oeiee52oECkGqyH3rWlQBVl3m9KGyaH3E5iME07wATc3+Jk4iDCwuYowuCyj
zu3IAeLXLwRol+rbISR3VezAAPuVRmPLapwlcNF1W3zXb1vfqWY3i40L0Q8Qsnt0
/YLnq2r/BTChr5/Z4NZ1bCW0+LMlu0CcBvNeYVaDX0q2JoqxG0mGlLoxbduT5oGk
B7FWmnVOfaP+QuEvGu4jcANI+pblcOa66tz/gSEWybOXaqFBMtyt7vYdwftMa94T
ppz9iOeH6gDImh3UFRTOFfYeHxjNfUfX48XylQ4JyvHrtIxF9cCcIhl97kpN2glv
xZJmCDQv/qRJAopDShg+mI2eQEtgWFczipfX40ZTjFLv0biUFfQ4pzNxncUUhyeB
XVlpJmAF5RxBpcMHtv1l8vr7zuwer8XoLGlWx40/qPVBgxrQSaxTNE5QsJ9Kg/IX
qHriN180NHSDEpMq4zSYyzqiPtaFVDTvU0yiaFMkWoeDtyBMdSezEycW0CSrbiNC
pkrk7dpUS5Jrb5rqYcc0Yjjj/sxualDRl3VeNVim3pjkwcF3hoscsvsnnhhMkRyb
uVz38MWFSmktXJ9LXdqOkFDrrlX0WJOeQEXVP2KAhMC1jnkbtI1mbHrnZUvglnQL
DQ0a+wfj7m76n2q6VFOTp/ar5EMq7rrZHcpFZ23j/CCYekUx3kcd4LcssUMet0il
V+YGJfxXX0ltKI8bSbpxLuo4o8h77SsP0tQr6YtX4MbwdwQuEKq17BC9MDcQuFQB
1lZuntXNcIDuvCMTMjxtyck6vxtaIUPDRR8fpudxL4SPenDm+i1L2wh9/fY6Pp9K
SQ22IDhj2E9v1MxZBsm9zPW/QBck42jPaw0sCw8K3k7iMXVb1+MD7Urx7kAXuJoW
DZm6BVofHbY7jeXf31vWTkoqqopk5PHKrv8loCBWoQcAXJDu39PS+MWOQtqz59/q
wGa4MVxUUJtAJlS/dCfLEQFEoP4RqnOlKCgzb7ve04C3Z1s8zee1HXb07EOwMGPD
/dhNTfKhp0lEVjFOuew4bKRnICqTx74CYQPgzaTrU0xhFtQBbk/Q5nhPpGLiL6k6
+ncYXpZ2SAz4Kf4wJr9vBLynL2ZRrsV/AwlSykyCjRxmJBoPqd0On3i7parGcE3P
VgCLqkduMPc3n6ADeX4kRt0Q+4hBWGp2jF/nEF4nfexXuruo6Ma5ghpMoU+Tq+oS
PwIwhQCBonuw6ZJfGtJE2iR7b82TCXMp+ekJppSTMeWhe4AlzIWfT0ABR56aL4+F
pKpnqStM0wnYWe3A3zRhuwDrc8cbafc8q3WjYmHbts8r+gObrQ4ZzjbrX1rlAX5E
ogd9XXeU0DSJ/c8n8sE9kxujM3ChggDJNvIZGAhrkquE/z6XIlG5rOTW00lFYCeS
zEgECOloILVYA7m/S1OyxcvfAO8J7HMLYp7odmlbxoJgzm0+YMk/LAXzaOcnQbuD
`protect end_protected