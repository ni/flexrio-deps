`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1HmsKLichBLC+2/sfbmxY8U3jfdyMosn2gBQ6C0ju6S8
tlNJwlOL9wJUkzptYblkdZktOe7/84dAc6v8XuhbsHuoq75aj+j0qASE2QLW4f3E
Foyds3OC1cIFGN59E33gytnDnLN68KiQ4NGW2AZCiNB9mD2SpZO+Wcpz0YXD+OM0
tPYFZzGqzyiebi0Abknlq0Ompf0GJP0LTwUU9Obva7lbZMD9OTwP5C8/8ZIbNeqi
KgdAFFC/jCLdDJBDAVsgUYhjSQTCvqrggsTjfvi3qCBhv6DTDIldeI005ZwnPc6W
uoOCvVlfjpiatsc8orBPR8Q4zztOqpz48KFMFfFODkaDGQH9NZe0pOwED804Runy
JkZdDrVhOi7kFMXH9vXRAYSSMu0kS3q7aWtDBaQWCpjL3k0Yka2zH5tpBGF5Dh+D
ZJ1upkaA87p9AC3TYuuXL30AdlvmNRH1zX0w/p2dmj+pOS4+rqczVo2oYOS2RFLN
99AqT6qRNRLVMiq1k10U7xc8BxU9+KkSgJxZ17/yKT/ryR/I4ilsAdl6HijKSbaP
MhuC1drmKd0nZLiQYxwDQ1feTNDn6l6jIcX+lY/QUKMjlEQeL0jF0clN/NfmxXkE
h38kTdZOiPtwdOw205ppqrkueK+qEtXaR3fq1FP3fEHx5NP94XR4eTnP7y5Wb/0l
WWEo08XeWQjjEPDs6VBs8AI4Jm/fNKHcTOrCbSQdihjZVBJhYhlxf8Ch+raax/XY
vL38W/Vtyti0Fyp1RqPCIfgLQDnb/g2Klubz54HCXK1kenU0S4BPksmznoba6MOl
ZsI06KTimV9bKVSkCI5RUCBUL8DFeiYxjfoxLsmNSLgvG3vr2urtrWuGpCo3PhDW
0ykIK9yY7/47LPT+OJRPHATDru4UcL8L57wCH7qBZ4mXsexcEuYI07haTTEeVFVo
lax+2kMfi7qtOnLI5Ta7naLf6QrlveoThzlxjOUT73I8b9xu7KPEmND88G5fSI0E
tFQeMzUgyQwqW34GQa0o1KHR0zlfXSnxZDjO+sJ8tZ8xF7A7q796sFbcVVyYJrut
6J1URxf/C/D0OX7HUa8Itqmb6G/rH0RS4VjInI9DwQI24AP0aZRAa8SSxScJ4zEU
5AwmcBdtYcApSlM4Y9p3goJOGZZ22UJ6OZaGl6ONIiCbbHrhZskjzi+etdsS+oi6
3cJr7Y4B4boUfVsqGChP44DWNiM2FFmShrTOLEyie3K/KVy13xatUvcIzM0OCQqp
pWz32l0clyORfoPNWpbfsxpeyy78p/aF0P8KGV0PRete4ywIkk47daG0y1iUNMFU
y1YVr3ScM8sdgtE+2oOjd6+yoZvBxpu09UkqFjkLZxV/EbYkNtbo24dusGmtaS/t
rLYTUwMqPwLgdKvndvtQwgrObCHcUtjzGHNeva0oGdPMVMQdGt1n02LV88kdzCZS
VuhHnjLIXYqNWhWjBnHtkoX3OCwn6edv2yG/W6ElWYeix2+DQn0ophkHJtzg3/kr
1R58geGCx1TaSo2otoaO/gB1BU6fuUr567nrB8MQK43+yICHk1fqfTQeZJDM13YG
VjT9Kbp3YFQ21bdRRqQQYH7Om8lsXCUSSj7lBfkREnYRJTOl91vdIcOOjjiFpcj7
N5Hm5JfBIwRZ4mRrGsjfTKWQOtYQYA6irEdu84zONXu17RWV/1O+uaA8UoarZqXb
JJta0asalxIskdOFivOZ+f98IHKSJeoeTRFfr8eJrVTh17B7v8WbTWLAY4jqDjSF
uRCXs7XbyMfo0B9By8azfEuxOYztdmExyH2LtQvhH3KlBcjLjR0isXlapIuq8P7U
EO3EPgeu0OjjNaluUJtnPmveywrOmrjJeM6hgIxxkTQHJJmiAjL4yasYA2TNXLPc
bz3kIEwJdvDSlTE5Fn0ZVlGl+E26Oyfh7hy7Yf/LrdWJMehnB5qjNdYlQmw+vFGt
NGjKjo8AkVr28eMpYDEogCDQmbOIWg2qbYyVSdhmZSq1rQCZbtJHvOip8+STO0Tt
ENPmAwtpMWhbzeahjtfbUIrhonLWY1JJvomYTdhY9QnmfG5EBVXWdjAXINhYfVpm
v+BgNq1Q0YQn9vCbxUGM8Bo3mGInKKhcfhB5OpeUtF/VD15hTj2u2DJ4yZq2QwEM
Lica5KgW2ykeNDTEJmrypaxTNxTM1NtoEKDZcWcD/+z2FnXGhsIWo9G6Awb+AXAh
URcrAJmY7nwF2LEulZKBcleNMO9GeriP6PuYStqPVfAYPOAKT2756H75J31bQAwe
ctaMrFVwGE9NrFpVFy/rlij7565Ef/lgJZ4rBBe3EynSxpDRw5oDF2z5rXKz3/gn
EwbI4h1Je7ZewV5hhaoaKGpxZiCrATQ4U4Rs6CDM7fT4FKE2rbEI3Cd9IYNmAKPY
v/Tte+ETCJ1p7IVYnSS+WbMd5Kcw4XunU0Q3P2FtC2qbyFK0dFxhJiGAy4yRW0ni
3o2yXqQk3J3I2KpUIil7Qp2XyTWqo/vAQed4siUF1FMurMcmsqAZ95yAt35yM44Z
KDVx7vAVZlVgYLW70CUw8REIVH0zlYUnbM0pjNKYHmZ+HzxUr20vz2BHZwz0yvTt
ufGaOjj1zg3pjiKSchP823RHuDwavG4meCIUbulykl2YJ2QAIxpDgQyT1+4aZJRH
YNNy8ErcuyY42veWP6KJEcEWQbtbfEoXW9U+s7QJ3PNBviWAW7Av0X0/x7yjcKgT
IRpvAqBDH7t26ZeVTtWaXVUrGIqvVcb+ug2VI+WDQ6stQVCsOBkjF/U3FNq2Pjwp
Ph+ouG+Ki/FqD13YNYSPbMdZxDdoSbDA4rOKN85LYlonRIh0rdnq4ayF8f5RWfBD
PAJ42/OMKairWuviNsu3+EaJj6gxtM/biZF5ccCw0BPw2VMCTVNcgWkABzF6rgz3
TsGvKsa+r/ApUSMUGYPmDa0VHC+vvzQ1lHLbrUwoyJ3GIelCVktY7SmfHVvWHrBn
GBN6YJ+3WQnN5O3jzljvc7lorCVdRshNIrLHXLFOZsgL3AnfiuHflbOqLWfiqVvL
xws8sWpkctqF4vFc49odEiAaKeBuBqwOD3O+ILh8Cki+DUkF1odVc/ZpdRfpP6R0
nPozB59Wb7YJa6W7N4SALbw3F12cq3yr9MxR5Ile2658oxqJUlmaJVglfSmYZLxt
HqGe3enUQSPpuzTXab/4s29SSO6eozqA0idBjeTvN8itGTQENyIRibYFMS9Axvt7
noZg29uc0DdvoThyT0tcAkHvZpn4RKXE9B+wOVXAQOWJHj3Oi/D0T6fLHQh3Hcrv
Jvy3/7RDmin2Jn9R2XtjdSNPb1O8iIEF57iPXaMmKQeCu43mHbaM0QvEP8XWREEt
NPSCLO6RBxvx13GblhNhHTIAZ0mYqsaoc2ZXeDvi92k66pUbVr+bCtDBt6w6kM0a
uoa8cUcioFjHYwHjq/eoTzu+oxjQCYqoc7jLR3pTkk7r8cPRkDasfyBHkBdMKVzV
Xtd3IFwc9T8fPjxCOKpbvaVqak6oofFzuiMT7RywX2Hdu4Yc69PMMlGv4OF2FSWv
gsNeCf61jUYCNIn5LuQxxUw8p218S+s8dHl795T8ENyroJRvP0eYEope8sCJvy7J
J1jmbTG96Rc7jd0y++CljHpey7pDtzEPusOvGCtiTrdt33iNjbcM6+CgE55AWhEq
2B4G7O9Qn/LmrO5F3e2WII9w7ucM9vlD+g0SIKPYJWJ1lIeLmtVKM3nNPfCmXGZs
5Cxm9jBYPEdZvugH/EJmk3sJH3e02Z7D4EkcW+S4SdgXnUNJbyrB9j6Ky3foqlAc
YS/bh72NOfN7/Is1D152O8PEkAeKhyO+HaouwKHBj7d5ypJMCtugzJq7FI2Zj/iO
Xr/1hcptzY2/xR/OPzz64WMvOFctsFQvkqMyLz9ljxQT0cM+WFweyuSOmxwlXYE/
qNWJEG2XXBQFvrCcJJmY8buEufsk3Adl/RfVyulFTUnqz22Rt/pqrG+bRsMyUgBk
KMiePYvLDZ3HnWmUBxIefw82T0ODyCUkvnhlGPGFj9Di5y3sWDremdI4uG2+gYIV
32FTE+LV7rOrFwaLrdQ7ReTDRrrQ7U8EjaZagx0np7WP3zAZlAKDBFf9VMsP12Mn
2P/k0sTzrZzFk5mcC8Uf+hEh/WmfIAgsvbYlfDbCv5nyN0Oyk9w6esUXOVnqqZZM
DSgStvWc9Tsqbnr2R+4gen0HN968UoAliCJ8pfG/R15QHM4nK6F7NdcrDmWMiAjd
sd+XEGucHMODpxYKHcd8SgE4R7Z82TCCUtp/gHox7zERxU6yaiLM3fuqUt6MPFV1
sug4Bpdu09dAFiU/MYQig7iG9xUf2VlCLg6hzOwgN5Ax00YQdi+f04mUmYXI+0RW
t4kRXUR47RFAVud1wMZi8V82iQYcm+i5nt2Ai9TtYtO4y09LMLwFhu7mwjPuFOmE
aJT9RVcEbxdCI9QXifneSJxJ2wG6MTkAUQ7ntxwirH3R1hUsN0dbgWWwpeDp2U3L
pwEM7tkvMLnfmSwcGIDds4R0u9EQa1/dHRbXvrNkegIlK86cMRaK1HkhN7CC3+Wk
cf1QT1wWKyln99Cuyg113vhA+1naAYhXAeFmK4g0ZXq9UeFPgO6x88DmDIBHw4m+
Yeqp4mH+Im4f4MO/0kQSSvqcup3rYBMk0Z4R4Vlq58IwXNF+EogtN/6r3FlwUQF6
4bbN5jh+iCTImLM6HHUF6Tna/ZPvdy3sfasEc6HJ1C7m/3Jl8/2uUlwqntt8g8Kp
agO6x6z4dDytydRoIDbmQpb7JwccNomlF9DA7vMy+md6GoE0ieLlhmeytpdNdnsJ
Bu4mcy72oyq08mJmW/JFjgx7X29XnNie3IalOkOHK/gHeIJL5tDwUgeqB0C/6ncO
mkLR7bBifTG98vXzwCD/aUlBDuNJGrcBo15ZXBYzOvGakunyzWJV4jCYgffKvUV6
URGfWIZGEiBgo92CKLRW87yESW9Q6B8FP++l2OftpEDQcZ21ArhAIvLxessM1H/U
2rUPjJ1EVFhyuAq7mMl4tXvijWIYL9dHjLEGFztYGW7D+C9fctf0FHWsbcdqekHq
eAj/RAFbKc5QibDiTgJIJJ/l9B+1VQZXxQeWTGyQarASEbMaUIP0ls7TMNFRZSoF
L/irkhwv0V0t1VDoJvIYfltuvpwbntgtrnYEjk5cmFapzewxsETHeypJnuOQ5LJI
BpahMg9jV2blFC4+iMNAPL+hcGTdMqfrvVSj1dzrMPNRfVaOVtJ9AeCA2SuvinM7
fOV/NLlRSLxAGFBG2yqib2IlrH3RLH778QOQ3UMhBBZwNdUDz49ikLpy3+zP03eE
PHGHe4c+hNAERjCwx6E9tRBvdni1gkdeiKneh9nBngF1xeBDbrglJaTbQbBFrd4Y
qqIdz0Vi8MV5RMwgmMiQVU89beUjpJJC1CBc0mHD5VNlZg1XJrIvr0jozhFt/O0D
ms8BLYbKr2YJ+iDaBhNxQtgYtmJmPZt4nQBFNd9W3HqW/QMdl5hop3Et23y7m3S7
hdpdI+Ri+x+91cgScvaMHmMOix/LW1OW3GbPSsWHAfGVS3JZwMlmEZ/ZR+0YaX8U
GsIvN5Mf9Dya8IVyFdDHk6TSWjpOUmkgJkwQRUusBr6Xdcb86s+7IOTxeMfRJv87
YhH7goDm/iN/89r18pyTT8nX5JwNCW09T84G1mbeW34ufne10YoozvIgQCv1X2vz
fAZ6dx4IjlVde8Lvs7Du8GAZKrDYe0npb07UYQ2kK473p6ZAjQoGw+4hZgOxvVoa
wNFzxC6uD2pRSkA2ALrA0GrXm4MWWq6y9WeTtbFYw+VpOeAnDgW3ACrwnSznNYYd
qhJgi4x8m9A64zfb5RYUA7xJBqHAB2iXCbVAEabiVS2wFjdh2XLOfsfPIlRlou2+
9E9bjMzGC+bo9dMbc79c4N5bHrk73OjW0uA/TSLfaNSzMkkMIBnrSQtC9fokKigh
LY3x6+yr90P69Ei4SAchHc7rG6wmMjKRTzDYeqJXVDfwkRpEAL3zFCPBLEVdiXfl
C8r0UpP5q7igqOh//puuyd+8pWU64GvH2PLxL+6xyUsw9X7wWpVe4+LE2xW1sAPM
MKOBMeUrRUjDARsRa8x70CQCGG6n1V874Jkt8kuQHfN4A+QxJwAbWB73cn2HkMQK
lUAPUSCjhrcSeCUKgG2xuN+ymbcLfMAoiQcU7z2nvIwZ++8CqPGkzGITW7EvLMes
Olzr/XKvkITidIv1FAa18zx9Mv1uxRyGNYDXtQaIIXFJbb4CCE5orDwKPa0pCAAV
uJgFqice2XCGpOHivg4C7E1VlqmCPpdPCuozJzPAJvZJlo41I1QO0tNncbA+lsEd
cfPlwGXY0FzmNwIZaqLKmwbWgFGW6ExXptIvelvpCswYwIDGaL3GcXLZBUMvErA4
h9wVCGbG5h4aM8wK3sWVG7OD/slW5VuLxaXikGhoE6dH0HQbpNalczULlzBn74al
0VnAGbxLXSZk3DT57oq648rDj8SffWsGxi0q3uCMaiUGxYGgCMcKIKDCjgfWIHOm
nOytiD7OBogvn8S26fcPI/j9u4JHzNNpNNoCOVJbT0vZpsqW101RWgopQi87Q7rP
4FAJfc/EhHBC9XF09Fkw6UXq/UZHBiFiq/OcJUlrt+eglR21UIyfSPqUrFhh1oJo
UB2U+88NthDT0QtWeYUV4mMHgUVtmri8HvTQxPiL0nTYSNYlPTOvbQQ+AtV1x5dy
PyFtNZLwfumW5eOqpnEfLaaFEVW4UVFH9aZSWlNAx/KsBlYWewTHNZ1bDheLCESG
0KM3qOZvC2nX543Cbp+jLDOGzsxSWl78eVlDZSPqMFsnbsUrKZXsPFOTEhoHRhGR
YRzVSUTOd11skNOwnOXmcKkkp+XRxBOvx/4O5SewFnHX469elupotxAiohrMxPzV
cF2mjfpU6zxqV56RV1AZBWdnUjPAPD70hDTnSiX9+CS024X1mF51eNovJ/CdYZ+J
8OJZv2TWVWurFnHVEu2ueUDMIAslR6NH1nryk+tjG2vlG21fSOmOpdiTZsKMRKVL
YyLnMe/FjNGXHslW5xyxYxxSmcageTOL6/MvwTKEfkiQ8n77uCKoX3e+2l7x5Zin
WsVl02g3RCwl5Sn7d9OATOce12SzhtRMW+WiY86qM1VF5x63mQE8q8eql5IyFv9T
LV5mqJr6PQQZXWFloFm+Go6/rp2jPLTPyu/9CcpdKYclr2GVndQAk4O6k/wf/rl+
SqhaqUmQ5TFtqo4WntJyPEXYdizVFa2MuBI95ArpcFvsuiejeZDaPKo5QNgnrNvg
8EmINYiC10PDtkkZnKeIPrUc9xyQi9Cny4NlhDihN6eUilYIX1b8GR0CWll6BLtF
5pJ3PHtiuAenih4Xzw3ZWpmMiwFeCu8nCoIJ+TZkx0QcZ9bhJ5NjD3g6vJdiR0jT
4AEtQcYLZBT/ftNdrXS36HS6K6F+W3ENPUsdP2E0tz53bvhDJlPSLl8mjvYWBtOR
s30X/PZYYUPI47OOWqdA+KZeR82xkUyIXg/LL+6oOK5yCyGHwGDl5g6UDJGAxruM
71jViiLd8Ty93bVJeN3K946KaLxXImWE/tPTJQThE8jHzbQQFcpwR5aHRumDeP4K
1YYh4Qb092Opatu1Y/Vi6VidJuozhj/kEFT9k0xuV3J6nlTCWGo7R1n9LPutK/gH
XiS11FdY2nwcy+xize1eIFlnMvVrUmw3kw+Ha2Phj2AWEWPnLi/9G/mWLyO3PB5j
CgEPC+uzo2aU1cLx1h5tj0fNpPrWf81dPx7Y1d+dhj6gWduOO6E0mKu7rJaXNLF0
t4kV0164N9yb5S9ndDprH/YyvNDfkt3W8LobE803b77S4K/KW7JX0fZwXAkJLzIT
7uvG+lTF7TRHxYY4ACubXnqPNsp02MV4BB+D4IdrqF6d1KoE7mbA6BdzHYHGOK4i
0AAfCxLKEAFf/3SpONJw9gb38VSx8hWSExkUqQB+MLC3620ADbvlrHxJlOTichia
GIrwyEV125yAkiFuT177+Wo7cOJXdatt21J3410Oq/rdGIHoAyetY+SRo0NFEyhO
ADQKiqoprrT/vNMrA3+Tmktfg1zE8G3F2o+b2HjFzyBX0oP4efdGX9viDVVONNBx
6oHz3Woq7wCbkkjOEiAhNeBRtIOs4cllNoiNkCNJhdqo3uiHPMalwVzSFLC83E8p
xRBaRy133kMKAeQDBa99SvrwMpoBrg2xTEtyvc2HTtQ1H/Q9+U1pUcsu6HAtKEMC
3IXTX46ypMugFXzPA6H1H8/M/zar7fP11ZZjxS2VMNgX5P7+jnTGLBIIyKj02UZn
MAyiI+a+6R1aGr8woKXZ61IsykHqDTztAdyOxErqTW0UprWtXVoYtPkReaa8g4g9
Dt6dw9+BK6+crbwo1vzf6TJ9853G1REUdVBA4QzbeAxfG6zciGPMvtjcFr96sIN0
Hd+cKuETI9t+Bm2jydiQlPcMYe5AAppxBQdzdP9XFijP7vQCfB5uMYXGjmNHSyAL
jgdEl001vqxqMrI8BApUf0kUHwHuilGG+SsC1HPfsiLEmGX8czJx9BGYE4ARXLIR
StGT4E6Olcddr0XokZXWGkuActYyzRik/XRLzaMug9TW2q6sr5CMLSpbnWkZvir9
ymaCYxlUkl190ujGGESWi6zCLiOC1sMeJ2bg4ySNWFvvnuZvRMP3hQoYJfRPnQ8n
/X2nSnM+wvsTWnfrfmH13CcqdHLotjiUKYbXdyYPER5WXiUylPUE6bCtGqIkG+FZ
clrTmFeUb6CNjZG+VVagHhUsodl6MXdLMIHuPIkFcjzIHBuXg6l5anIcLEIfQCat
PfYUUr8Uyi3KH+HVukRhNn6da4O7XC/nIbWs8yPwMDd/tkhtAOD1z/Lz7rw5rPtD
GctcQtx8eLbd4brdFOHB6Y0Ezx7g2h8fqAw45Gqoyj/OH1L7hCYov09Du+tFeOXV
cNJeNWdlzfwlDSW1O0rMTte9Ih8ywYPc8CHCZgKKwBHALkP/svL85llhe0GxsFzf
mVFF3pOMGRCRKh6GXJAgGoRZZZV2aJRhR9XMnNlQjU/7TAWhWnq3xj8kNU7FDULo
samw+dtCZziyms381TuYqN7qV5FnnO445IaZO8dXrtbbVrGNokwyBog0/UTEkQO2
3hghulpMoqTK/PNzc0ugInSjcJ4VZa27GcTTR5hAwZBcak//bfTCuhjtEqeu/NDl
NKUeDisny3hpJCGSy0A8OrWYiP1ohJUM7xwSM9Z/WY0SFd3hmLAQqDbAJwnIU9b4
eMWNIrf9k4TKlMRHcHbCKFRhrCbYWm24rdxuTRBMPoDCbfYyyf6D6715f4iMaMDK
YnBytseyjrmm1Cw9ZiFTNkDayM9Y3dqFcJNgaADSDM7pQy5p9E3oPbdrp0faKUgS
BrVNmu2G/04MCtacfnla2YNnI0ZX/425Nz+tDYnJXGOmvDh+nxCUEc2b0G0eG9ms
xjKcUbEgIqUjKJSm3d72qdJOaFWz5AkmcV4YEiz31nj31S7W+rc6AwiCdhG4CwTd
FriF/nv2O1fHAXz1o59yMpEO3IiL2nT9CLcynp89cNaM0dgwYe9tsmOzSiIB0zpx
/sUu2GpDdaJddSTHiPWhlH1Kc1gHMi8jorivQ3acdwyQ2Xk0z8vodQ7uFYZpma9o
spPDVgRFlLBD0D8YKI3AY5X/O4MAF03f1dkQx5raQBZJvGFMblPa3c1MtR7hzIZl
EL2D2yshVDRncsmAEpyAz1F6uTfKqgMbhRyuAZTbguJrW+iRVGhIMXOHn8tAicE/
FK8QP1NNB8f+zHWv/lqL8mphd0y/DpWTM9Ynu7Ovisd2KQ6TnO4YxTpp/q6XSvrN
5G3hAyDsBVUyBKXdvvP0+bXNvE67XsSy1yTmE2gEwdc2K/bhT6Ey6n/ZVQoEeHv2
TILa0saWdu+/dHYutLwOC562KMGvqWEufKffziG1Cb2rLMniBeVyAzlfSAR89qj9
yu5Qv7YMpybHdiHaG9TcyU3eow7al0LtlTM73clBMtxUX4B26zhgnLxzfJvfzdTc
TcR48j4kBlrxKTl4l2Xnzg7n/IhpCnPSbZ5RKgyoskCQDg0hORgCBonAalvAOH+Y
rugUMmER2Hf+XanYiML5HK1ADN8GEG7XnytOjHFAV+whLcnpZnQSwdn3tST/xlGw
mNI1VQ75e42Mx0s1ymDIT4lD8Akb9Hx5s3XVpa0+0X/Is+PnIs3N/6qNNN8L602M
nww13RUB5WBZvWnx6z1IndMK/f8m7gcP0VtW26LL93qdO9J2Hl0FVU762xf5i0QB
K0Zr8CTMKMKRAm6MSYpnZYbnrG1gplbDiAz5ck4hUzGtTsdcehnekklFcHRCIaz6
6Y/waj09rgyAMA8pDVaEAUqN858BPGy4UZYpzOkgisTxuxrhNAGm+PFau04Or2od
3T9ZQ4BviqfG1FDmj4u+kl0XIEZhm2H6DGvMdGdrmpfDwyETXlCPMuJ8RhFo34UU
z/wZWCbTfqnjlBnLcnN+t6QSjWS0Lju76wVoNj7KbNe4EPdmB8AgfasdorShYBv3
jhwtNn/Zlj2ZaMjejIhWktRHabLmgEPu7wpMR9hBBMLQwvcY/fIEpriUvD6l1/i8
VHZyi2LIWrVwLIXPybPYF6sx9hL+A6n6G5r523d6fs9XGiGOPcsotZGzdMFLn0sc
dD5zB4rUECdgv574gEhOJlEzdFVTTJdU5yLhdPAa4YyJXhzlxwL0IkzCN0oFboDA
aOayjKfFlMhR52UiLH3GPNJQcDLldbxdHuRoX1BTQKm0AzgQjz9/ffxi4TtuW5iE
EFSfVmqSoHOGGQx7/ZXk9ZbvUQ/+HLWHBFBduGu3YrbgMj8vRyeXvdHsWbTUoQTj
T2+5FJ9A8UOD3ZzWSGMeJR82quaR0EP4gfD9zEta7FcezHRBidTxcb2vBxSaRtj0
LYsDXXhnjMVAnCr7P1gNBT6SmIaip639p9DOfDMTOJfe8+2RcSeP1NuOVbXsSHQd
9Kp2jbJ2fFxD6VVt87waxJC5ioAwl8vCYFjAxkKNAYjQr94vwspp5eyNHDXfzn29
h7BQRFEtBFv8WN396b76y1GQ4pRLRtV0hHKwe/j5Z7FqFuUXJugPPw+7c8JVM0r6
yKtoTuiwdaOXEidcKUZAzk74sxpyko9KQPeGGBwak8EAJ/HlwqOEUJGoojQpCzBA
WS38WUXTIhcJI6cM1yL/xIVsypmALY9rD4RJ+uB4rRIdPS60RZw0hy+eAD4HJZVF
FVs3cprot5Lasea4gR/3tjphirW1arfDoxysDQyrYqlAZDK/oFuGtmCYY1Fggj21
BzMT/lHHE8CaXuxWiSVTR66Sg9h/mGjAYTcq4YtIpizqMV67Bap66Cb3HmTuWYeB
4xDLtIqsI6P3x3L5c91B+4G8QaxSzsQHnEVOLatcUKTx1zuV8dR8wdJFjv1su80t
gOXsAdkeklmV/HdybVIzg6Nvt4sD4V9f3mI6iVgvytQcbdMcpNvdAiHZocbrvrWu
wOOebehkB3IKOLOqUKdqoUiBukHDdD3c2CCzQgfve0SbhmKIEkn+rkNCjU6JwwYF
6CD2ACcVsBOubamiJL6Cz7IVaqQl0JkEQJwyxLVdym+BJaIztuPlMnhaCQpBOn8S
fRhwAoq13r5tOf0D1iJFlL6poF2nLCd+m9VznGTpHQUE2D1hk+rtKKM0M36fFY/V
v8XVIwrb53SRV3knNLM6/B1ldPYrZBPs37JI4XzN3FJ0x2q0RDYHV6BBcWsJiomW
VQkCNsIA/mHKUDkqRoYrSzPqip8bLAwn6QFtpmnHrSIoO+FdTftqFvbZ0aJdsKuy
ajeVfGnB4uDyvU31jzMe+iuYtYQchw9NWF1GLNVq8jMM9G4ZqwT59W+4qo+lpWB+
CYZfpE/mknnNjOU+eAdV8Glocy/67COUhlfCOm5o81eWkvUZyUxKhmzP3guvb+Ec
9PJQdoi1RdrVh0qLvtm1ipwUI5+eWKXT0m809QWkHxi0Qfy70i3VJezr9Qse/6Ae
WVAlzaWPoygEhsB0Q95aJv2/rFt/cnYcW48wo60vCuzVdFSCBAeXVYwUDtsGXEsQ
UXx4jdg2Z9PMV0KB/YJDZB8CEyEmLVFWnGp/NKofGDCCdCQ8hAxNRFotW3aUMbtk
znfLSI5L/xfY9LYznLtUSSBoMlQSKej42tgivp/1teUljgIu0xaxkAk+Z/Wf6JIK
dpNuACrQhk0CtQDAEo8LLHGeP3eX97S0dVIJkSsA8ScBZh+bSs1lR3KWL2gjFsqG
dUJ29PXzzLlAiJhrtJKMlBsaxb6VQ6J7tMN3zLwIN4ACOJStX0jO+87SB1kWEyWy
Y1K3Mel9sKYMABBTEB3S1rFcxNOqWY/s3vBI1VnNagIETkmaL3hNcGUPyoi6C7t8
yk5rAV+mwlTVG4H6j3RCPdQBC+R97NC98pZY+egRjgTy3bF3pc442fQFyTOFGgDL
LQvlfdDiQABaHDgy+Jmx/z+6WJQIhGoQkHOPPePowsS1RHlwpRo+0IZn0BeyrM7v
eWgP6jCJm+/hRuvGZuGcT1iKoiCOvLrQCwxV1HLGwHqFkj68EAs0K/Hz1IbrVJm1
G7ac9Tc/dO395YNzwBcdCqpMZsk6AXtd1B+Np4LGVzI10usLnBkOhXyT0Vf1zFBw
5rEECzAhplTh5Kj5Zdi/+YMY+KgizzXPqTm8LASZ9FwSOSTk5Kt+QdjF6ZtFzw/G
qVS4/xaS3t69S5TuzNaBEiBdnarfoR0V+Rsa0nf63W4UxiwJfpF8In2aUa8SQ8Au
gW0XLsg+IIW+fEEe/Xb5jT5vwFh4EDhELIpmjC//05X+9m+XzkiiwG50jzhhxDhk
qiuIJK6X+RedRdfZYk/KY+SeA7KeCspZfalrwWrJgV4acQhqWDlfQk2wdQ3lxyin
C0eAGXLpPOiGD2dvQCtCuKVakJ0QO0LELHQgD4Y3PRv7EqDmqQ9JTJNGSBMqkzir
F+D4B/RKdhMwuc9HoPoECCLWMMc9mKrT5+JTQFBFc60s5mIP/jLusUJyLzBs8F4Y
VdAEQgqxRplNQgyQwqihs4it4qxZU2XIwVgE9h1WfElG+ic5rhWKD17V4p17cvhX
ZMHqXEPS/vX588N6O42Wmh/TrM2yrr1rWYfO7GatTF/b2xxpppD2Sqtpz7pGbYlW
DYeUJm/lSkP80or3TN4BrHmoWoDIVUI7y0cGuxn0YB9VYJ7Vdym4Lv4m9LHPuBzh
i+D7ByMFRVKpdRmrEpjYv4G999LD8UT8v0RKOkRuh+EIzQdpHRs+ucpToPoLIrMK
A4s17+G2EcPIkBmQUZC7uLONx+46AMpM3KaY2YuF4Nu3Yh9ge0xq+ggavNoNAuqW
3qfoAy7rI2yXERDd54NNKxNWuZ+y3btjhED92kRe8Ti947dus6J+Ijh+Ltly6mJn
3n+PQLAVRsGOTsc6IXa1mNCIWdPNw2gWdKbkaVAJfM8rqe9wxhUsF1lYibQ/qV2+
hxrHwdSAtGAjI0Ypmlir3WqkNX7vGOrUadgNQy1GVGxkWNVj4dGQrRa3roVQOOmU
2Cxh1x4v271H4wcT3ryXe3XzBkIDxID6U32uMpVEbehDF2IL6bCfCBb6C9AMme9A
yp7FCboFLe2BiNEhsSnpcZ2Yu28Bkrs234dQFx1h2x56uDphAAlzUYbUAgdewxTU
zTC7QDsUH6bir6Ic4YqP0xSyN/TsueGRJiQehf9hNCGkNg0E9ypKeadJQw2mr3aA
XD5h2uQOt7U+Vwv1CaYjBw2ySWdPZvJXdzJQZm1MFvubXQ2eXc5UEVMo7bbnZV+f
hmt0jREL8OH/S0QfE7pWa7FoN7ImH+9kZJBvwSek5hQPRSIk2HJKhrUt4VIeOB9F
FxNwJehhe4VTYMv7ZYZZay3cCn6A8r0/y6QWXgaYNZiBxlDmZ8G3+Ul53c+ilxtf
91MQ1gU/U305H5mCAA8rrW2N8pmQJgtKbkDg6T2tVTmezTnpFBHso/5zmjtJOcEj
AlU7UnpVKE68Kr+5NZsS7e1scIP1WFdPlXDIv7fQOlnhdogTUAuXJQzdfakeXnij
t5SoxHbbYoOcenQgR9Xe/8QxvNHg64gk5kn2Zo4kuYwR+I87MhFbclH+Zk3gfBkG
chWw7zSaK9Aw3cyeid9dZx7gm7b6EXEOoBW3fi8aAngdQoMRySGnfLnGa7k3e+gT
TQ+ZkaKOz1C3yNngEwI6oUiSLZQkmQ77Mka+WOuPS2G+DEQgWoZPNHsjcJ99btoo
Tgms5aQHurMc/RqSODLB2CkbAVNk2VlAYngn4G91eLpVzuKdxBhZ4D8PyTxltaqS
1fEXLR3olfO1LFdmhqPGX1YHVDUm6eB8+nOgJl7VSYeSa6d1JaLZ3pBmcpsjgXvY
sv9ac+Alkx0p65oEiKSuFJGoYHDlA57uN5yrJMBJo3ZUkuuvGbW390Ic53lXTTa+
0nr8RrVWyCW04I7ZD0PPUDRGiPA3dKxcgdWp0d2LdCA69Bs7Q2RuVAEJm6ehqssS
XtGBv13/MQxr689q+0hidn6hRRXcybHzqpZbMi8CE5MYjvzDqqGAJnKOqOSzvQ6+
cDOQnEJtOkbJDn8In4dCeQi38VucYmkFkxwl4mjb4tuWjmBA/ZM+SIYT++zjC03O
+3iLnOH2E5EGagLIFWrE3qommJ0zEAlR0+tJVF87Q8wHKFcx1jxxrfpeB3Y1zsCS
W+JbNFJGVcIrEZAag2X17X77GQqoK3Ye+q2xCnOcWnVil/1cX+h9THmEvlsL1zrc
/aIyqqfSVfhAowpAhkBciL1rVbtPLx2hdG7ZHMrGs9icwhEYiBVPFp7XJfuyQjrL
XCpIcOWOmk+9TIrtV8gqvNXFaxr7LFuev5Zkouu6vhdpvabTVFYXawuS0bfzOu1i
PBN4whceA5/dd2qjhb45Lvn8FKBuW8oWnvo9Tbq5Sq56J32llI1Vo82UlfwT+M0+
p0sTXFcDx4vZid+SJJ6zc8Ls2JNIABCCIkAh5e5lq6VXY7TW9Te9noDPySmhLh5f
NyoK6V7D7/3/mwOLWJZjDEL6Gy2DXMhmx268RMClkHvVcAgw3ZkTWeOva13m8dPM
X6d+aw4/ZXehRxU4ZhPkVrYPlYdnGmLp+oLQjSHbgVaS9Y4NU2uMB4eYCNt8VU0u
o3eOhGcUkStE3qbdatulx1Unmo4nLekXwl0/mEW831JbhdznHisq7ahThlw7UwoT
RaoQBe6qaeyYPpQt1Z6MAWsXx0NlTjT2D5gPK/Ip8Kp0XDryPLsGQ6Fu9DTkjDzq
ZaMYMKC3cRkjxYAdZTBki3MdOZx57bPyLPHgkeDjTxdAYQ9sTmm4zrKganZFQf1o
EikBFBFtsPkDuSjKRVj3gxMc046CEAVw2Qiq2L1dUBNY1PYsZNGF79c+EBVRdut7
/NU58RzvfwC6zCG3ZvlBJAz2OMsvXatT/ma9Xe1twPU3zAHuxloVRxcFbAYkxJ0A
gBM8dPLz/rt8DPGP348DNaAxQykIvLmoSuUBmChCkpmmmuwtVnjf0AKpNazzZKQI
vAaTN1tA572PY9TobaSb+r5y/lP+xVeDnAt5yvprYiPQ7vYiicozjutLInbN0Yal
TpHd+QKB9EML8lM3q/UJexqXqNpj4+xh25YM8737oP4RwlcZVUIN/4cB1qFdRpp0
JrZlhn2GUdaC75oIzpmeKL1zxk9+q7hQ6ywANMdiC1Mx0WtrK1uY2Pf36+mgJqqR
CiXbR2hKGq4Sq++H2jkBIfubvi58bZ2Eu/NKpCpTnYRmxeFzJJaBKKw7hFP8PVdB
hBUYAWrINc1uCAp16/Wh1e2N77h1BDs7M+ENu2TH4BREAgmhnm9fkm03siPJaFg4
sEUIJzHgqAvS/MYd7ZgWwvuWpDGdIo+t44NBZ/diL7uoPyZuGFwwtyYumvDv+Byu
XoxnKkv7RSJaRWszWBiBoB+i/W3JY2WixP4mvw6YELUa4pFMECNNnV3gRz61bob4
f7XUknBfqiDqmCuWB6uFA3pJ9VuShJ8nU1ocRboRoK3/c3K1BgfXsQpL844qUMby
4GwxalRXOknAMArxlaj8VYipzzBwXnzOqxSoslhNPAEQYsvHzbiJaqGoAE3ghu3k
9ooT1jLy9PdrN9LkfY5P6tAZ2ajSAvarS0g8clNi3QRNQqB5T21hrbtLnUUVt+ez
KaCcHYZng+RhCq+TIuLvnYrKP5l4MxHVuuOpEDGFZr0NZGtiWFhqMsHlxDI63uBh
kChm6v8htvxzU//Q40Gm8eONg2sTJP9SOaswmLlgBji4jWA+uwwPskrs1s0mSmxO
Ab3OxVPu9v/nu8eBBg/j11NPAPUKB35XBngm1CEF+L6U9KBrTYROsalZnyKUBTH+
1hoK18mc8PncYQFSIIiYCo99qaqZix8ZqPA/pTLzv3Rdmaz0c4JcSjsX2LY6+GmE
7VE50IhqoOk2ZOdIOu0Irk+mN2P1ianiMV+SdaH/rMB2N32korvymuC8XZdMPmXY
6YeZ49pt49Z4gzc69GF58PUGwfP/D11rkoLiDeFCxXmbO+oj5fLGG443hIPPmsDJ
96hZj3FoG2QNjLIN/drlXcgUZVjFS+GwkErx7pEm1Krm+AFGA6Qt9Xq+2CITcUxR
v7sEAgQ45XW4rqZhZEQ6CZeldwnh8mpB9km8DAivreIq8A2hzYWoHNJOliZMfG56
Lqvucs89R+dCNPrp17U49Eh+4FjpFRy6nNVgjtBfQNdZrTdzb7itm+aoNo+GKXlQ
arx638RWpFkzeLA0BzOZ+OBbaBQ27KHhQIl3xKB0p64B8vH6N8w7+vkUHkOZ7NgU
5AQVoKbKLlVilqbsrZq+RHQqZQhI3DItswlKdBu0emFdoXOtqFtwufbus/7tAiRK
JwMi4Q50MM9vayL7e4jXYS10iybxucciQie/L/Cjhm/MApWgE4lQkcFZLpZ6/M4F
ovYNjGWj/TJCq/xnBmuxRHM1NhcsfU5+71sadxo17qvuh7aVFoLfJ1d8KnyiyAFC
k2u5hy4xnABYBqifOmBTgsW8V+QNUmpJzWZm2QZQF0pPrn7qsaY3I/Etc4NLiRMu
OVuMG9hZ6UXS6BacguH2nh0amclmGyFeixLEH7MK/pdtzy0nEBaiRP3Y+hhi8e4Z
OgSYBW5OTkZm+KOX7vlIIPMb26aDedWCCkyGgOYk+SQXFzXP34+5F39NgxNI25X7
yjmFHThvFvnwnpIpgIU4GO8oqCTzElAi869swaOCzAACXhKe5aZuwZon/jYHlLvS
i5kloaNTdRoW0Yih3iAuUfznH/7rsp9XkuDeQOZQ+elIsvs8vNRVS0IQNoZaW3AR
v6qssLfb2VoJYWfrgXA4wiKCDFwASKSKIkFWhZcK1PqGZ/h8i5PHMy0eN4AW1uYA
Ed7QAmV1PdQPW4ZpHqHb3gevR8bTRlxE6oW0CFKYqC+SGyc2w7cSw3eFF/EzcwD+
dUt0QoVJlmU6lH0fEx+FqAV92cqhGQus9+1dVUUY6vwnqbaY9K9ZBVhPRDyHxgMX
8mSbTGyluvzxy/+M5rWL1XQ9f+Y7UYF5wGch2kNScBXqdjJJXETHX6jxMcVw96J/
Zf7ickt6lY+FlPE3c9WGEWp9gR2PtuwI7/rC2iQI4fwKB4DMVgGNlJLQCvkN8YVo
6VKXeA7vRB7zkkmzpxl26LlnK4VptmJcODCL8D6zROupx29Wm+F2TA9aaqqorYkV
beXmcr1MvZEWb2K6bXwm6UukolYakE1tnL36PTD1vZw0snmBQF8kbkX9a5j+yv/3
K8FnBaVmLGESU9aXBhHjgSvcfJiqOuJ2m8RYQdqcsU+TFnsHpi9I34r1WCKHzXTH
gyOUTgSbBrAVg9pfox6AETbcDU2zqjUbZZpieKK7HjFgKQvoEFRJtp8VjlPcKRpD
WBqYXoYlEgroxQfKiNGe7C8ByFVBA2lCd+cskcnf4y1TRBKrNkDg+49ojfIFUJxl
vvGLrB2T/mpKSO4GZYeS5+Dk7Ze0WSkzjvoRy1Fdvt39RthS8JLdvE58Rg1FOniO
+tjEf+s9UPaE9wQOVvDejEU/nEoCHc5FL/OSFbI/3OIfDXq2cYZThlQxkt02fqi5
9V/7BCnjit68D0J7d2Px6AU+iOGpsn/gAzrxndluKEODfrz/gaBQ9N+MRzqNFFRu
ICJ/+qSDTTd88QondMmJPbwt4yNUcP0sbCJo+IrzLcMhbXOqZU0hBjAP9/DY8Emk
GTadBgUXsL+uEcJcVI6xt9SctYEckg/23OiDyHyK1G+G+biloVdqnaeLUw9rfArG
SZI49j7Np0uCirRPcUQhDqWeUdODxK87CpTMlM2zmG7eYbr5jQ1T+lXpeeWrJRsT
7I5hEJhVTFnquT360t1gQ+ftTYJqnqjXvdaCkfFYXCJNMxS9+nLLBUtW/lkXqsfx
oSoGMWuieBrYCQuu8Cu8bzJs8HznqhW0fOWBPSBcmfYpL99VV7kOVE6LWe4uVCvh
rOtcifTp2HSQ2W6yxrKuIuvEI8I2E4FTFnIfqlreJi3NsfR9HleY7+pDP4gyAuEL
jOnFHLmMPIxqztvKbRvShJ2wIEecYsigzNCj8u1OE6LkdH/nUiSatm5v/3tfs2Ip
nBdU7XoAZ86MsgCv0PIejFnXvfs28kvZKNLpLhB3aFe5LZW1RddmffeByBVT/Gqr
jMSeAgd5G0gMBvaOE0q8tqksXAI8aSOPrqdXMQwx7JiuEo8pRB0eK6NZPWmaDtxl
HkC4DXtOe0SMapVH+1VYxoQVbkL+REjarbVy3gY1UnJtVAd2WMIs7hWIdc0HXlmM
Fv8OdDM4SJqdYcI6cnUGnKpjhTTaBJVJ9xE+bDn6LOBACbpgUSVrPQV6/yrJ9s0+
REEu6iiO5Ge8lD/rPKZiJh4y4vOe8ky2FQ4Z0KXRyP19jguYSeS9iHkPM2tTUw/5
WyTdT4v0sDDZXx8L7FBYK5XAeKMs8AxY7XnIhPT8p8gj8hEoiXs3YBAnmjfyy4cb
takpGsTLI+Qj9a++v7OqrG7fjQ+f61w7YDQaXhZfJgsxfv3QNxRoeGcUY6BzogHS
Z4potASZUbIF5M2VtsSCJYySMu8oq/auASVquTVNJmwsm6HM/7z3Rpa5XS+VkYJg
jsOwzJ8qA8cRb2qHitYpTsBeuhcPkagHormlJ4vhl3zjRg6ZeMl8GWtK3rrDtLUO
rIakVRQ24De68c18h8r9snRqZzXDMRYpVUHi9AkFpI3Kq5TTtlg9i9JkqORU+l2L
0NR1bSJmlWlCTyoBPaJ89kqYoVMXTEAbwbjnquzVshT5pdjqh4UMxw1pRwwOJ3hg
htJAMYV/WVEpxWvFGHNSahrLGM5IT7RKcNyVx4RNK5bxMtgGeQkJgDmSmzmvudCS
HJB3CL4c76hNNKTveIZUaRTJ61AxSR+k5Sk9iN4E4uUjYTRotAcfXNJ+v9VV/Wr+
AN/1H7R4ULePn3LygmzTuxl31UQQd4t+2wCb5G0Wf/XVD1e0X0hKnsiKIfqtT0hM
qCXKfZmeZ4jlk6fhw3K4vMewNdSHar5p75bFUcM0B3FlDL/RJwa2zpd/9yUwYaH1
sLF6KP4Hbjbao9Ugi5uztQujir8rIjVwclxkT/5kxZz9CnT81xExd0MPMmy2FerO
BHD0ywu8w9K+XBotTIsWV+3+I9o+ZN5Mfcw8NEN1ooBtoojh0pCaXw1Sko17WkDV
sCGk7XEyM6Mo0W2B6w/HBk1TyZcYw6nnZ/B0/1EB+DX0hQZOacUPlm2KSgwGtTCi
Res4JY5VQjIZGyW6fO8ZcvuFPpM3KpT2RWNPYcDO+Yhugt6X/BX7EgcDao4OJS0h
QGfPtxjSp+Z+oOJMES9QS/6Mhq5YM3Jj1IWi2B2k230uZ8TIK6zQ7uVVdDqV5mbQ
9iMXIxsyp1Ir1mpKHZFXd9LivFGFFQ+J+rchWsKhj6aj5+pQRHUhk1DBPQ6IdCv3
okD/sBEylymmG/haGqXC9U73wW50YVzqW4nGYlIjiqIdxhfXPJTPzXHvDjLVvbKb
rt5vD1gzQLakXLdtXBq7jIuCi5ZB4awor9tf3WuJ/0BVxMTbeuuh6OBtJ6msAT6N
Qr1bVqDIlgtWv6M4NB61asmiHp9hPGd5FY7wSh6wEO4wIoexvRFbVjGD68XNgsDf
+ol87CTvAvlVI8bCPLL6vVhFUJMYy2E+NPi5wrWL6XLXdE6U+H1RTRVIBYtr0Mr9
LJVeaow8mDAd8eOSnzFudClnqxPyU+SPvAlKUBmlEqKj+5/n97FSPcYfzDYc4hY+
ivs3B4lLg/PI29APG7rlGsGaS/eD6dUZXVYkUS7dDLruW/lMLqOTHxrkZvVcTWzw
TB7lPIpfyv182t/dbfbtWqR5uCPlosdszLDoYztk3WZ3uFNpzO/K9CTlsiFCchU6
Q6KbRg8oRpGZ3Fd837y8IP3tYXroJeLtlLYJ5UIzoL1SBddsF6xgNxLoAwX1PYKV
to/rSJ4MYtCk9FQIZr/ZPop5B3cSyHOrMDCE69W43ObHvspsWXV8w3jNKgzbna5E
PiRLNTz4fnecqQSSxSdBLKcoSZI5y4fffD6QDnC764GufRbgPD9/t/9e5AbNwPLY
5W4T4YaSKHLJgeHFyroWm1VLIYnZcTkfPzXWmJNSOV4HpgzFe7/2AuzpkMzrQi3n
lQpJSnYvMjEMChReCnMg5Z6keapSnDXLiNv1zg4SnQ7JrD57z4k/qj1VQhHff+4Q
P0x/6bqT0TC2C2DUZhQfTIz4ElophHaNoX7jcqaMdZuDm01voO4aG53BHSwzVRf3
lv//eyH5WGYElyV4naaTvK36n+0cyjBgaCk4htxdqrM/5JA68NhpFZfcJNL052pd
ZrSazjPLU+8ZTaf7iBrULh/yA7fzIO8uXV4HDD3N/ivYt0P5oS6wad7Uv26jCExU
KtrTGV9oXUdChztyDkLRReAVf5yimkf59+RyUGa8mS1+ENB8ioOZAM+5Bund48OL
GiOtQ/YhqkrZX1R3P7J1tH7zpU9S+GCvafJlgMf8blpSHPDnFAHkbX83d3Yh4RlB
nrLqGKKzTW4zyWSIYsyWktXH24at7AqUVgh2vpqpkhy+dVWytlefUAvlWaGORiad
hR9RxHE9CFl9jCwJUyzJMbeyQl8pyg2PRj/crNksPDzwO8c2bTS/9HpPKgHQDiIt
1BDI7GaHBFngGC7Ozwh4fohg6b8MohDbJIaavrB8UsopPZLyaxOpmcLTxiFU+bis
zFUd0IijCNBj4QQMSSj/xw50Twg1/Dmo7wQtCZhWAEcvUn+6kxyBdie/ifLAyDAW
uZRk3ee8ikPDJ9eaQVgimY1/t8C8SkFLQDfIubWtHG42iePnMGlnDFLi694Y0cA9
0/nwbqHu8UESbjMOdgwuYz1hodsFre77gpBjkeTBid8RjSP/2oiuSV4p3fHIWrj5
5wRg0eAe0mK520QZGlu5OJqLswuQr8jv19GioJ2ihUe3lWQpWva5p/SFzuMeWImp
1SnjD0NdYtFB1t7BnOh+O07RKXRUhhFXhV/V7rcWmvsvuiqEmtnPXUQ2SG2d4jnp
xCcIUtL347FJTQlHtAyHzgH2gKyiuf9iirOAzCNr5kXK+tMJPpDb93fFt/1quPW1
v8EWEu5kwnhn2EqbQNlzx70MKexshhIVK7wyGcOqAyUK7JpXbgg1uT8ukHCrZYM2
54pT5hzTt9+4y0Uajskm/Bf9v0J0UabwnF2k+TvV0CgF739yhcNPhdfK9UYHkax6
TvBKtPNTlQomoONyr8xPRuaA/towypxpIN8LZBemfDq36OMUHPSVf7lk8agQUkie
L4K/ZeClKlL1dt3f5fgsN5GBSnRQCAMig6GnA1CH1DVIa7VDAFGF+cdmraEauOBf
ynsdoW00CvsY5h3SM44HugkZ4605oCJyFu6aX40eymP8M+bgBEx7v34WzjatyiE1
lyrzuR1nWujxhnc/8unJvzhzIaEBjQYk7U5YZOgh9YC+sG320fMO0sp5lBamDSQK
zAnC6gHQ8FQpOCKZuBEShvtRloi4SZRat0bKb8DE7Pmeebp2QRN9QEqr+90G3GhC
J7byhuTA1oGw3Rlz20MxLxxokgA1sn7aWKWd3pzy4NRLUQBYhfXiTI+LYnztyQfi
7hVGEHJ5Y5rORo/3QKV+gHL8PLcnU1banRbwM9Jg48bWFqBkgkrTiCNgyLef4seo
chMQ/e50/DSZZFwe8/qGKG4ZMs7cPh14q0Zaxzh3yC9TGlUwVDL3R377Rdtv3Rxu
9g+KMb1+233a4vWEdXUc/l5Pu/bVhGbdlpvQKXQKtRSCGqyAAO0QgsKCeBgcoE2T
iL1aCW3vOCTbJMatn86kwHgRncF9ohsKmcetyVI6irlJEiWFw6ULjOc3Ks0/+z5A
miIsuODiz/xAnChRDyN58IY1blGwqp0NznKj1p5bU3KYc0XI1cbMgDN6T+9PmhxK
QuUcoNoAH01uiZKjbCaQnH2LDoT+GzCgrot/Sge6crW7HfgaNwGrRWi8Kqzyrgby
4KdNa+1k6wHuV+CoQ9sjhnuT+DXOiKM2GckV6dbXMe9/Lpxse9N91Tes5OALRgFG
b8ZasfYD3TSk5utNWE7KyldFwT5UWF+cIZhwSHXc5D5dklu/yRCAZJpHatD9iPTg
SleUS53hf4ZZ2w1vZC+3RTEBXsARpa4Z1GcahouACvNiPfHjB8DtuYkLELDTfLGl
lOCk40/EfMC7ereVo9K/IjZcPxwtTtRjQh4C6GjLHn5w13eJPFj8W2f0iwM9TGTQ
Xt6wOqg5rjReQEs9wEcyX/37HQWG/Z2w2YkfetFIsgEYTkIoJOze7UP3jwwk5q5c
c1YKQpbVfzifbe0EWhFU3kaltNnlqxA+BQDn0Wpcopn1SLd0cJw+ZGAIyMcl1nlj
X8FsJmGmlPKy5Bs0QoUfeIDqeUZRBv2xqpgouYAkdiNmrIcx7bkSgfxdeqUDb2mf
9x5wcqPf/4j/SIJl3jxaEi9L6pf5NUOn7af2jbf6dbD1b+egXNsIDK41opY4SWT9
AOVg7798NYmJq7gD/gu5H5N/GBwfpsgxhz0M4TH2K8y27OezVQ8vfZCx/7i45AvL
iQ+HS4jfomv5sOsy5OREiJTdHVOLlJBUWWOYpFeW5IQ/rCMKkT67VRGffBvxm7z8
Ja5Fxox1awPl9AIzMb5OSbDJpexNBk9iZAr1izUZWDg/j2OQfd9IFV63m1OU8dHj
grWb1KYhlj4fwyDIVkuzD4MV+UCCXl53hF3dgdnv80u7pB+ptuRrqQrNQICiRYCb
a/ec12JwAriJftJHS1m1kBroZoESFicvOzEmcHzPDtaOHMHp5E36w0QgT24LNgF7
f/RQEqpcumABRzcOGhs7rj+JK3zzzqLwq/NhEHdzuOaOC2Gdw+FrjJBcc5HPCiXf
o63KubwW+r3F1PsuEhZneCgc0ceKZja6FlAyo9NX7PkQ5kQwh0YdfieXmAq5BqKA
eUOlzkobEx+2e1mDFQ4B+Dqq7uqGcyeE7BnmvxYutRUah503M2haBiNa1kdkCsNi
Vi8Dwoi4/iwYeOjG2lWwDIcp83ZewU+Hy7Juxlnci5iWeVV0NDktRry91pMcCyFA
n8eHQ4FpyCZsxEG45Yh0d4Xa92Z02cobasQThzA1S/MxWN5vK7D/AaYE+07okZZX
YTbqltpWHkivutuPv9MRQhnDX68IbSD6dhaBpq6IHWC0enI4fvMZFMX9s3Yr6BXP
VseU4nOQUbJ03Q854jOBVCYwUZQp6BIHpnazBxxOe0CwBiu8UyTTIIohRNJCwAhZ
RtITmeXC/5FdVaKdh/HAfcesMj8GLRDRip3TwCVyPN6YXMZgArCiZSUYeOybjixr
oYyDjMrd+p+mabcP4lxtb7PoztiPl3u74nod8N6i4dMkeT66SL88HYfClCBeDTUm
EHxwOygMhw3Kz+pGk48Zk9lUlE7ZgfViRrKnsj8CKccDfj/6XXMqfEmhcB2IQzMh
VPl6VBxmjLVXCFxQwTG4rYGN/E0wgL1I6qLh4IDt1K2V1EUiIyhZgwX0P+wWF8Oj
V5TXuFfUmqlDKdiCjIOqQ5tPKPFSDXKjeOBZqdniw60QCH+GL5vCGefcwa//IOFH
vZ2lROh/4sYyXaJy9l3QHli2RtzGI2xg4D0BTwZ8Nk3yCxUphK1N0h5Ki/Uxa2XS
1miwmgAahkXJ4zom/ciIepiU6jxs1qGc1RoEAbNmwjzFSQHNy1RSpiLxb8IJ0PnV
pJuDREnIZIPC7rRNyflLCwXJ1l1vFq3a39B5rY3g3jvNTw/UHmF/XGwTJx3P3uGn
eQCGPFewHUMqqT1Ci4/Zp1GH+bo7o19RQygqL4wfbhEupL4urY4KRrNlf7f0hakW
BQA0oDL7CHknOVS07OQbmWN8eKdfJwdCuXNvjFG/UdOB+MfkHz7LewTRjy+bpP7L
036mQwLGxIvMp/lILUt2DTIZkcLej9ULhSpJ5vM3t4WiklvVZjekiY6ElYqzB908
ZTabOnB0N9Jpr+9sgitwvpKAJG3xQpnKhR1HWv6imqBnPSDO0wh6KBnSz+r6ctdo
hskwgt5drUR99nmeMsLcJWKjl3qm5Zj0hrv+iqV378cuBa84mLSbCk9E/5xFh0uU
KU8vqPoveQCtk54WIlWcn7C+8WIwsMK8RzaAfaj464cyURsEDFDuVEOXBcSDkSp7
JNS5gyWE1NVhQNR7L7ZoCnmZVElXabEZ5J5//kke2ZGRA1RWv+RSTbarix8Wlnms
swXNleQ76DhvAqQxDFs8Ch4rLplSh6RlEpxGFUCLQgSMucsNbyaJawKimLlpUmZK
uQWp2IypvXhR/DynDKg/nYywOK6beGYteMvyGehC4dFHmJrVk99WPPK5DNc9XWE+
tyFjzPa88FvlCLHpZ1hJsTVuPzFt1SaEgOre8WVZwRY+myrr2rusrpjo1qsYkhvy
JxooeIEzWb+eNW2zmquszd3yHMZyGYDLFtmMLfj0CckTjwHZElhC06+jGpaYwBry
08y+vO+ozadLCquT9+W3U5Ajpoj71wbbzeRApFkKSPyCx3TpcnqXFWbvwBATaU64
etOIc1RqD9JRuxBNBPaORH9UxSBRU/37b/r0GsLkehgqeQgKGTGWDwaQ1q0QnCr/
3e89gq9xSJcfTCwJkM7ifxQsv8ga/WXYFLZxWBH2Tx9m/9CE1L8uwWq8FeY6c+Ng
4yLV3VHT4/0K2anH8qfS0CheeNOxnBBEdbuAIQt9IKcvV1xJJT5cmln72lXQeb7w
pVreDi5XCyV/7oPVr8Hib+Jq2YLhgPu2qPK5nAfPsITkKV+0wqkEXNbjnp31NwVM
XNNP58xxgfcnrH+C/ZDr07KR4aaXhAQTdBX+Dsm0dwKTvLE6nvWMelitB5940AA9
7PqhyQnrPa34UPOSmGVhozukL8uVVn4bNiE6txUenCTAsY37p1vrZCmwftpMaFn7
X7+T4fVxkI9ydvlZBm3GtO8VgZsjUfivS1Ez8xbALeivKsi2ALtO2JvKO+vivgPj
fcLAY1ws/EkOYeWUt6WZ2QJDHLonTkgPjUFCsJP7sZ/Dze94vOBba39eYx0iAp93
KI+PY0R83EM9ElCK9T4HoDg/q9k6yBbirc1DPrRKLio8ExXjF2IMyFmEavHEUk4f
IX3NxyLp0qo36mwRZxGVLZkVN0nCYDg2BhMCEcKNBorMRJGiulvtIRAiXP2fkTFc
bYzzYMvM+CuQXcehE5WzxJ/DqZHKwo6dbvaaOIHXiQYutkOtAfnhI983frFvmjIF
z55g6n0i1XIszHTzsDEEUXapIAAHqnb7BjR5CyuhmxFUr6E947CH2vhgclzQFzVs
5impyXlKKCjW/u1m/tqsP82XJ3f3THVoZ0FhsdZbXqEKWzTWrlC7ABrarTkGD8DP
Pa3jPusQSvH6+RX1qqKrehXdgraPWkqyS/jS6lYZrd4LLPO0dop2t/9PxViC9MDO
V/MYUuOorXLSVw0Z5CgwiOlYPHLNy7WFthDw7gjMTAG4YgTbmjaHtxe0eDumnELn
SS3mZJuaLf+i2flh3ghxgQitxumVElYl/CIELiTI6fGoR+9XLV49Ry2aktYaqVPp
3YkzACN2pW0OFZ25ldI8haKhTSs9MZMqavahA3HbMRflcMIZzctBG3iIWw2Q1R3u
djENjdBaR1pJ3HUtwgxpQKEe4QOjqPJTBooyclxA/Vuqkv0Cijouj5lo/y2FbXHN
6vpA5Pa+ltQNlrbacOxuCvM1Wqvfy5KJCUSjiKi63iEoaR5Yqs5XfOVLrBEofN+Q
xR+5pCXU2rlaqic10rrkTbiyWSMeGN/iZa3Vut9PuAEqy41CIAVXxUeQSNnVAe/Z
9pI0Ml5DV3B473kq7OkJBUpXVGuwx4w7uSFNaB3WksWy350Jiyu/Va8o4GbF3Ki4
iPizNg0VtQx8c/MX6z4y2x5d3ogIgWK2i+WAHIT/LifXSAJDU9J7JTW/eZsoZoHR
fCsT1e/OpMJtV0y0u1Zd/cR5ScjKQgu3hjKd7GQH07FQr8N5Q6HDfc54v7MfcY4O
HuttfP262zEP5onUIKXt9Vib0MdlKynsC0yIMkw/PjR/YQnfhmm3POkq5nsjDa9r
6dOGAI1Gom6OVxkGd+jYCwkNr7bgfXhQs95GhPYjdr6x9wp3d0F0M8HrAJ+Ix739
v9mq808vPwTnaJyhiLepRuZW4jycDF8pDPjSVEyPP0IYcoVB9hbsiwQfdRks4ABa
eyT0QkTO4AXkecN0EwzMAs8+JI/SxyN+v3jDZvMRzCv5eI5szqeao46rwUkPIgiq
Inx/nC9hTDlqDSh5vpuEVciCbE0WTgW7pX1o8XaqxdxgmUI3MWj+30xfp4ocz9+c
sLN3EUHeh40eOpDbGlZfutYCYsSDEoDklrBOrQkFNu/PLjWI62pmceoVDHcrGwx1
uThmKurYjg9Nhkq5VXGk0TlSe2THFdIg1XSfRZ9c0ogsq/1KjN2LzYZS+SFRufI+
RnviNgnJpvjqGV31ExSh6akZw8iiOEBgOCmm29240bDxo4GjnSC5bQIeZLlcNPDU
3ovExikivKBYrL35n/qwFoYIko26lbmIRbK1Dbpk1dNzaxsKPqs5gu0Ba0xQleY7
GrHouJJIdMvPl+rmKmXj57fhpIZeN1q3VdbBykIw0ppckrIxq/AeU5sL6KTjQUvc
WmY+7gj40/Y9mMpIYmx4b/uVXF/wpMSjiWUVe/V32eDxFup5gCqvV+xYmqHFbgDE
EVY3Rm+xO5Xu1GJyhCyCAti/8/+8KtwzmacxDcGTSKQFwEUMFdcGqszN0adNSp9U
aGDC4nBLcYggrt99GZHzHOelG38w8yMfxze/czioWUvxt3gzQ2w9Nlt+dngj9GAi
eAM60E77rpVJrHn1fKpzHhBIIfPoShk2a3MpK8viElVPClEOyK+nvGz48gBAbksF
Ny2k+Htkj2blkVblNcskKqAwRank6Ks4gAM4FgXrxpjT8m7Hj8aGtdVadc3NLuMn
LguA2nrdCzhVePASBZsEzwPTQxMZd4YjPSCjLR1YXzN/Oj89KKT0DGZnv5r5mQxW
Yggddb2CTdNmRp2Fk0H8Ke+VFTnTl7T1xk7qzeuB0kyK5hzszaNHWvNjDxsc4uyz
6hXGI2H+n7kCTuFa0DapOkT880teyKWOYrxwT3eQTuxv+XrOYCLxN205EwrCJiDy
4d9jJeNpi1j7lBlq1YpqdtqXTK9wfVzgnWkMfUf3qOwDoxP6wV1O+NVO59vKHAd+
TtiQjt+yMsgt0zs/eWsTXoRPZ9H0HfDOhe88BvdLT7IuJNGBBflKQH3QekmBkxTB
0nr75jGwYM7ycKGAMb4hH9C6wwz32vHxBcVd0InWomBtXEWj2eUxec+o+lq14TLj
9HtDzZDFEIDqLeB1lVssv1og+x6oixhBj9y6mrjhWzgMjm4GUNPaXH51Wnkw6pUJ
NdkmtgjukJlNLSaC39h70q+EVi0OTE9594ah8EI8rcu4q3iElfIZdpNl1u5fP5DN
xOcYTZzclSPN3CEE8HEX77O15BVdcgqP0wtqb7MOnMuVQ/5jexOVIlyFOnTuiwmz
hpUrlrJTDljaHBK3gzQ2haFxJaLnIqY/9uKsS9fNzE/lpr4hNlZhnpgOJyidfI3p
wHhwzJT7VJ9GuYw4ypiUFUnFE+urtPjl6OOODL7aOjRACeBBg8h1GsXie1i0Yprs
4cjnONceQBUtHErv7pYv4rgcEe6bM36jCSmMTezo9YnZQAYnxwy7jkVIuZ2gxmQE
qBA8ChCjtcwEtCt1TFxMXnCjxizXbjLnIBPRsUX9u6nyXt0JdDFNu3iBWFfa4R/q
9aeQ67gQkl4qMzekLSUPbtrpXUK3sVDx/EVAziXGHqhKbc5r38SmPUIjIuDea40T
Go8voDVMPtAYFoOAGHwLAQWkovJiJcvBEApooz8iwnsTI85T/cQnHTHj9NpLr1fz
NXRFdYA0pznQxSAIUmiiJBD/3EDjxL/9VfPfSARIqnMalxIjcEo1boa70/TDtA/n
UwezANShmvYFa6CP3DVMfYxF0RAY+P26cTKTEzcEYzIzbd1hz+KVrDJ3NQUWfelE
nWmNz+OQxZCH9ZVXpCVmN91C2LGT0gbFr1K15I60ApNu5QwDPlnsXuewieRyIyxe
Bkjs2HyZ9tl4vjfTJ2Q0XxK7c2EkxG6xIycnFLGK0nbo8SodzWhd/iNTWZESe0nO
LPhxxfIlB3yjwxdIXjRLnJfT6+CSIGplpXXLVFNn/3h4stfqGkrv+/v6ufTEGEgN
mVSvCm6Wn2jlpEbXG0Ydx1jARXfUv8iy3K7r2MeKJbiJGipd/xjIyrwVRZYrB5lv
LAXX858U9nFpL7X60ty8dFIG98xfiZxBqZDlzUBV89LDJLebCG6sHkyufAlajAT0
tq7WMV5fkba02OQ+6wJNqeiJpDns46XTDv8Zh5UAxHIgfaHGjrwNDTgBGTQqi+Y9
TAQ58t2GrmR0xjdO+p+OtVB/j/Jul1ynyPOUxyHZBLz9MG/ddxmf6IKIJ6rcYCdD
DlIfuaqvQLOg0mleN9lZAh7Y3uvXNkx0Yz4+hcv1c4xw6bn2j1UBSZZsSjELXPLr
UZ8uC9q2+SgI/CrzzjKD4ARfvMMnvhjwwgP35kYOznPCqUfR12fWkt31INOPoF4I
cMExQAb4+KruQYX8P14xgRAQpVk9KM1KZgTMosLrAFCGDbvnVBYIiyJSU0xGeUj2
C2uE/26xQw0owLNFL3Y6x2A4Gp3UOKPYCuQ64JoDnzwfzzTAjnRVfweVN9dZuLlf
tToQuRgzB3fCnOWF9MUikz0/9/p7U1XClp5xRFbJnlPrfTXWOdP3K10dq1wyjI4c
3wq+V23uT0Q79kcgb695IBIN3CGyggIDsGLSA6NujxFT/xr0rm1DrfUp/Xaj3BIe
MOKli9PSq3V2D/JLBrk9XBl8XUlJLwpPSen9BcSS395126AXrnRghQrGZiXUkml4
iscB4gYn0XV9gomlOKiQy8ujLyLg084eM+QDk2c16c5DnWuFyQMcZptt4YK7mwor
qJ305pxzYFiS9TiJza3i6EHp/xq5GTtA3QB5Vb5h7egOWiB7mG5KudZVTKOaljFw
bh+tz6K7sbx4SzHbuhiY8FoWlUIW2S6UqlmSvyySWP89YhL2WbHoCPbIJRFyY4ZY
Zubpo717T5R2+7+LnEBS/RnCGUoYZIoi2wuif7cEkDZEA1oLMDJcyfsYK7dLwZbH
9w55hG2yOVdlbqVO76HI9bZi6ulF1K5WGcIlr4PvYe0lAmUNQN/1V8Mqs1wX8Yqy
zYFJ8LBY6dMzV5OZZxdewbn7+cY2nkaKgcjmFAhXYA3XJQrmU92yfdS2mtO7qNtU
2TXaRV3gCDv/vQfpcA+XUOJljBJLZfxlAU6hHiJgR7uRpJb+bzm5bAmEIHc5GRdN
YBwNceUxVNMeXQ4NuLNEwurTYcoFWhj9BMdsRpQapgqBllRceJzpd+BGSIf7yBGO
sDQ7Lp2i0dstR2fBwEyZ2vOcdOcHOxHSOAlerAtRJeKmvc9934HCPFHgSG/oVTU9
2fdrK8wmrGQN/blUBgK9VpPAg/VLb5UzefVEku7KVSj95k3IYrZm3GEiwUkXtqrd
9rrzB61AV2xjCwLXqbPLA5cnqlX0dK3p6zcKNBQOHSJKF9zlPT7YTA1dJzNQ9Jfc
z/F2mQiZ0Y3qwnXGOmsCn84PYKvcy922n9kzSy9mhjQFNtCGfmWYzWQwrmkLa9mS
+3rMMOvD7aL3QbKYOYX6iNRE+D/N5Xsz3irtf9rhOYEqWB/Zf0XrzgOMURWNrnYM
73zf/pT1elBRr5V3xkbzaWOqEhg0Mt7bUpxJlBntlCJP/Du03QFpy4lzeyIaoPNP
q315X7Ja9p6Y8m279LrDW7LhHdhKgCtCKvmPxdQzSGfBcY9A3dh63rYDCYMaNf1C
tnBRPxQh5sF9pf5ACMbvOWP1eV0uTlDFQ3Xscy/1mnrGyyHHHo8GJCc6X/Plb5jB
zSkC6wwwV2Iuazi0YJXeXO7S9aFeOaP+ZW7NTIprASfJqwbVODp7b0y7uC0O3rej
C/2zDQRZBmrXzYZVLn5R+pDRBKYpobZiDXuBd+TzzU3YjaupuygNOW/pEaV38gV3
cSQebT06bOvAF+Ghau4TTSDWlKiEbi3xYEvjwrIGxVecu8ooufIlty+0Oy71ngKF
0M0Gj53iGav3xnVroz0bqOX7WjK32E3bZ67lB5qlCI+he9SbGZu9y1fQ0tGpZsHn
ct/3UINcohpP4s4a4Qt9syGZ57GgEvd11lUVZ6+VxDzcO4nhEKp2G60SN2Zg+Yl0
rNmSZ+Unn3Fjhw1SdtEB/pC0OJ21JPEkUUPRpYt+rShmNczsAMrAQlrSfa0RSKEY
fm15KOqP1FlmXWyB/d5CV0shshJa8/nqr0O4QTCyW0o4fNPqRsG5aKWDs4zFBBPp
uyKRhSz+Y01fPBo1b0X8K/YgCegopn+iXdFcg2X5E+Cj1iwRGaBPoBaD4NoQurCP
Es3+NjiEYQXa5O9yt7bFQk9TgxefdvbAJgR9n3ya/z+GBdE9SzF4InZ94NSg+bvl
gxPt2cDXNUIxeibEy1Af8cFSc87Ym70pgDhi6MCppW9O0BnBHUl8mIUgm1zqcL/9
EBbZTOD0LfQB5wTEUyswGp8E4rUIiu+Lmf4t0CzlXR4YAOgr8QnWCs5pc2t2v8DO
VtCsofRI/lji0F0XWEAIEoouZ8C1Woz8TIShRnugvtyrc8SSqUOE8xr/4c+0cA2P
cFvCkk367appBjhcBDGG8mhehpZigX1hBq8yFDmE7XQkKQMl1O+GGoVpba5h72by
8saFa0LcIBfch/wqh3PxRo4BOiXipsfze0GB9EQzD6+E7686Qi7Gf08h3AgqvlT/
s5F04kYKe+bL8gzemkK79GTJx0PFlsSvhQRKI3/sBwxaj55sGRo4j4+5nnRHm9Ke
7iZFw1l+0ZJdqgwEuBSDAhjYkbpEy7O5qwGEnWXEjSmrdFUx+tjNPkAMT4145oAG
OuvZVzOLRL8CkV1dKT1WIZGuD7kfcGjVMTfaEO6kCR81i6E65ChfHT+gidvIKv6U
+GuPLHIt1vgjItFynE6f7RO7gGve0i9k1RCUYbfl0QqbICRQYibPl451VhAvHAub
7ik6gFI2ekrflkB7RE+TXg1ofWVUiuTZ5ZtjFm9U+YU1Pb+2zPxX3pZEzYgiUD3J
8vdWBEE+zrDceHBeTTiOATiMn8pezzvB7b4vF68kkHeuANt/BJPDZfR67OWa+XCK
5csLP595CMO3FYIEixYFhDlxPYNDQcriY/PJdBkzYLisE3CFMyXtiQTkyT4cBYcl
X0b2YPBDQFiqG3zd5L9tMprVqnmWnN5l5G+b5LdYDhr5uOVFs1RMwe86M3WsnfCq
IKP7FjPMqfahgPz0sE1nf/GS6wlvUbgFy8MznnaVRKTvCfXANlmI3XnFG9TCnoIB
HR2UKOaqIDzVRDXxmMRPmK+lMrXuAQiN2jRJ5oxj9kXYZjvaVsssO6zTbIrmE3Cj
ozK6ESWsDWz5xcV0gUyrgIlBJUciGXdohEcgylilcaF6xJ8J61cKZlq5FKEoxoRg
DqsG4WXeDvU++v8JdNCJCN+YYFoHy8tE7klANYl9ewjOtUR6+4xrEduL5St9MQGz
r8VZiyQbef1f0i5DaRcZx8td53CH9brW7tqDGgAdt10ZoS5Iyt6cFT7Lbe9KdCCU
DFls7MmLj9jUExwmX++Bhk0z0i1aLB64wBJkWdcxl6xh4tgiKG0m0CAqjWi1JO6d
FenqJ0u1IQRp0WZW0VRuOPSa5+BKzYLH31bVF7g3TcdYc2reVnHTr3cs6YkYEtB9
JN87ZgfK+CVQJEXs80OU0quRUV1gk+5UCDd3Ng+lFKq9/l7+Z+kzrKcRdc9MXaff
PrsZY95XQt5NkCslRJwhGBoQeepDrHvDrgXT2FDcwJTMor74N0qnaeQQrRfcmcX1
rHeZ5H0Q42s59GEaJwDYcdBPGQgxYBlQjiEH203AfFKseRQvB1bH3VFxr7GdCVeR
NK1r/JOzfE3TfrS9PnvNonYidq3pUVqQxAkq/QyUzG/mKYRQSgaYZJww7oOfLJIF
4tLl9v3E30X/y8JwFIXe/JXpMNAILPUcov79o04t96E38NGBRQVuHdbDN4FDQaCW
AfmPCZ4frVZaveBLWLilFecO/oj0ZFuX9IMqhBPj2pBXiU0aJPaWu9kaXc538Wl6
mahv/If0/7E8plceahJsI+28hoA7lpc9PHmxp3zGFPF/wE5xuZYmzsbzP9FQvXhj
Ap5tVyAlD67dHyrOn02jS5DAR9U1KtBIO5TwoWAQWBcWN1JF8Ku4h2TQ1OL+QUVj
tSI0uAfQQXcMXT45HH6JPZHgasgQv5sfuXLuu2LGEKBS8b7Ve47Si2WsAbQ2FYtv
ngK/W4+ADHt6K+EtSwxbW4+Rz/eOccHOJdFmr+StNvBhIN08XIZKZcMpgW+U79Bv
4nNMMAYLdm9a/68kL2Z2YYMuLhKWyfYlbj+5t9jBFgGPRc8Tilsr974c95LelKh+
R64WlR6dlEvfL1UEH94WIV/JGYVna8YDK4Hc2PgFy3C10h/HhejK+LWKMuFV3X2J
X3Gtwd4pSfVBzomTuDkoUMGtAWjNRpo+z/g8cycphc/z5wJ/Kt6jaTpCw2LTm5h9
fmNrAQZ+nQRIu0kuaIKmCKnhzn1aPq77qDj6LbDHg5Q/YmeBX92gxfl5TlA6NWFT
5+DL4JfIxGPYzB1cltzr4VyJHe2TxRHcDVSLFUlQamBF63+jWrB5/PBjtF7OA3L8
F6sLmjxmUuMsLU1gZ7JE7sMqkDUSOzHirNDEGdWxgdd8N4quarOjHp2pxcTBG7t1
SQrdm+f1GFGmy3g8ogqRjPgWn3f8p+jTMcYGgUN3phjJ+2ggUWAJKlbQbIBW9pN5
yCNnezE/8hnqjxf1X66TDVXI2gF2KzXWvUotloQL567S67EDMSzivWfftlmbJ5WW
5C7orgYshYcoGXT9rq+OIFScjDhPOFBgaiLJZ8+g/Bz9+GhzNRIjV5wBKL1hFRbi
hZ7mORSy+n+lwEwjCZXrfOxUyaz2TTrq+38yRRB98nFjnszTwWXii2QetH+jqvZ/
vQHgjH1RIG4u8HcT3upjPxeX3RQb3HXb2dOcwOka2RvNB6p0OEUdPuWX9amwsUKu
CJU07gWCj88WCNDUPnO39Tg7aYcX/trpFUFIl2ZgAvLkXI+ddu5gZDLqrgplTdWk
ESdx/rOjIH6/u2dl6Wc2IFLbnzhS4ii4EC8lewV9tuYWFoX17Tu6rl44799FD2Hw
Ueh88yO0Y6nlN41NCVjC+Iy5JCnBgvbSrYW7TSoS6gVIPlVb2Eyfyo0b+AfDWFJs
MSjI6HWRKwlSQ7AX6t34bMl6tKgDHaTxCwuaIvH/6cUdDyzhiM75HvBtzRbObxMA
CGK2RlR3VMOs0Mkz4JvN6Zly2KFlETYfKciyOM/1/qm5mZZBOfoH47LosGavKI87
rlNYnQ7m/WAjAUFmO9/jzG6h1XQ2TVCA17pJZIgmmhEax6iL+2O6juwW2zf5Srp1
rD+D47NDyyH4xopB+l4NCrvW5/9PBfQJFAHLFdNJkthlYxw5AjLDmHMUsrUnXs7Z
i8uDrLxZuQCnSCuoLVrO8ZJ5CszKK1FCZI7gDFWiMYQOa3dNGGJHfN+SFJ5H8uW0
Mzd8G54AZdH4SDgmcsmKrFYdan7ZIRCZ9zcTOuRzu9XF/YedjVfGFzsQ8bKoLX2e
B1Q++jGJIAfbkbQmE10quR874QMOxjrrEMofXfD1VwR04H+qCCDMu3jNAlTOsnvW
JOJkRanuaqsmOGUgeYKTUu1QlKu7cz6nSZN59/EYc+UrZUL20/udybrJ9ykhDLcp
yAyny/j9uhFDxHC4G0jb8OakqgzsDjkq+bVoRIkHNOhhHNGKFKsQpCrG2qTjMt9T
qloyhj2v5BH55or7O9WT+hhTrkz1+BOr92JzxmTLsuG1sUxmMETwi/4uMgpSPAD2
lDPqdlOUewLPOHwTCCza3qLtzhL0FPSICKucC1SHW2ZVqqnBMsGQg18NTYMJoH+D
TR8ty4qk7rqzzQ89fOn0LiJR8+zsKzj9Mz5hQFhlShguL43ru25E8zigrKSvii66
V03ypdtuPofK4FDHwZsM6492HolOqh7z57R9FmrWlbiJYE92Vz1IrzNJByebYDwG
+W53kAbWKzk4UvTXbUu1AwPImBNrtmE0oxISCNT+L0l5/o31mlLVZZS4KnxBYWwv
kTGgsRz+ydGsEAffUbEWNtxlNS2r3EntVsuhDf5G0GOAcj/em94vUEa4BULJ1PyU
Mx2YDilmLfu4HQpLmPWLG02tgTPuZ4Lz1hLRWJXKsde1i8l1QCpvVaTz6OXHXHB2
p3Xhj5opXQvdv8icttFWmeBQpTyDxmP2YglMEOuWdVnHQQONumXN6Znq+eX7mFVI
NP2NR8M8lvvE487nIcPvEsLVoxh7GenzCm+Le3/whdOLeNzm79Xada5E71Vf+c76
XkuvxKAcn+rtDXrKqnQsXJ6c2yo9UAuF9keIkNyGQ0OijvwGis6a3a2zls/Wuo98
oAi7SmqSGdjtY9EGavHj+kqs2syA3kAnGb8Tu1fKhRrXfqu68GHgg7f2A9y4XseL
2qOhZv/qPL4A3ZymPTQvCeP639XeD2R4GueDLnZHiPhMYCiBTgGN9S9gI+DcsJhx
yWLABVHqTO/Z4tXECCFQnkpmpMe3aXX+ZDhMWoVH2cjHC5VZEVkQPNikhgd6x9/9
/PYVTUNE1wPe7OATLOqmyovHc3cfISh3SMBkc9tbveVIJv95f2AvD8CSmjmek+0/
A/26rDhB2Plrb85zLuyVsvT5fF7p8QRAjgnXs4PvItfnkxd3/uYjzshkw95cwNRN
v+OkBQI9C0empehWBXcK46ugdVcov3JmRFGqLGAIo6sFIIhZWq88VcVwDe+VErmV
bt7dbbJYn8tGEyWf/1wIrcISWyXURjhQGCtLinqSzRccwA6BvAkmptpgQFvmSPGr
rvUTYSDyqzwqyX6mtNY76MaZoGlI8puqIiEtZoSowBna6cBqyzPgyk/u0HHqroF/
G/s7OTFQ6xoS1nUgUNDwP7jLs3iQl0WSBlo/YTa9/II7Tozw+2NyC8uy9MAUVKtW
D78xjM1ic+cEgJfP1rB/UJT1m+REh9P1dIVENV6Oa//uWrVKQL/zGO1OiYGS8IqN
1jKsUio6/hNM6kgnjKxKv5ptotluZD0Xnvgz7c6FvYzcsQnrmQnaS8mpejnNvw6T
XT8ZCDh9Jrr4j97At8US3vJR38n2UoraMFmIoLq2ndFaLndytwR40I0LJkJJ0ON6
+Cy52dtuG87hLHwhZT4II5CowKcQtodYLZh03V9UO3YdO4XlnY/+2MeVM90lC5rB
g7p6jT9pFlgTioC4sxIA1EcfzJ0Fll4bfNyCvdLiq4McCxqPNp3oeerBXQyBI158
QkxDvSdRfihfXw/7Qd+c9Tdr09tqrNMGL/dWRPPYEkUxeiUKh+v7nWjtHVP8x0xT
BZeiOUl0EtobPAOOJqinKjbxslH+N71pFIZuGlSG/RdBqEP/lF/SAr+sWYo7AFWu
qu552OFgbwfxWIQeXFey3lRT5DtbCMKfTZeNw3rOac02cfUhyLGURSAjuAO8oLmD
ifKrT06jZBlGKQESLor5C1pk5a+bjTM+OgIPZGraLTkQdnLCYpwX8cPE35LClqKY
Olj5e6O8SzMbI1bo6sI82h7qfuH6yxVQY35UwVM8cL1a7qlVavubNR0R0lSkJ4/s
LPoRxq+OK5N/PsXVBs/So7NPHGRgAc6Vp73N4n8y2x4alm17JjUfm30/mQDHFBYm
mQdK/4ThTm1i/3rfWTWpa9f876z+v5fFq+6w0sZ6Eky4V1xZsRUVb402hubbxF2P
PerHS1+/vgqJHxTNV4ujI4NPbyiJIApZyhIdGj8rqocE4Fb3wSAbK8d5lhM4G2Ok
2fU3uVrYCFYpBt6NBKNqU0t2BNq9JA8K4EavuQIITmSbOBxTkAyCFBEW7eaJwmiV
Mk4ax09bHCHs1vjkyGni4ezKQG5DTMH6Ojd/6yw1hgpZFRyluEu2ZSIjIM0siY/+
k8/6InBLWkQNGrumvapnFfOq6AKbqo8/1HpEhDcYuaFabVqS3NH+JM5GkkMwDNVQ
5v9PXyj1k6cU+Drinl4UG0WrWoDMds8M+bfL3nVCTUDe8fYw0UIekXl/ZAbkpaA/
d9cl4aguABlJSR1rYvmcNFW7RiS9lfFF57EKCuOS96uy5ASCl+nPZdaL3IhNCY0H
DqYI9at6FB/MaV8p3p6n9o8k7DYddHDlIzYnnxUfZg424mR70QL/5+12XtwAYa3u
NNvUkuNnUgD37zIZKTkhwsmwnzaaGXDnjk1Bj90l+LnziIjh0RCGYS2fWwF8BxUj
UHwq7BtD2ZBl7Ea7hmhGwLkqZzKctXLLreNhKSUgcJmM1hyl4Fw4iiW43FCu+Y14
rdzRSIl56Gzla0QghsImjkDcwdhRnEIYjfW+fhqoKGMLeUrSN2rPfQrMgLyog3wP
Z1PBrC+6tR3EuyjC451q7ji/DyK8mk8wszXIDbrom2iVxThYNG1m1AcjR2jP23m8
nhH2IsHzdNIRzdNEDi2C2iJZuXQMy6/SSb/J42B5VRn78BtJAtDGCgpRLtTKPkcO
VJpEBQhkqqvTix7QOGStH6IAk25U9+xowRBe3aPrJy5FOTjXh/GZ1U21Bwm4LBFL
pJ2UsEJFT3bJh5XrZXizVRJRoWAwxPvkbkga8+ubTwvF4d8zBu0K4SbuH3gxn7WP
W/GBhUBqV29KpNJxEJ00Z0bfywzfK84a2EkCDFmZJsBkNxGSAxitG5cdOeTWrCdf
wUPMUTdh+7CNKXFy4QttZQZsIadzdfFUnDDODKzzSzjsT8eFOBKIDt+jNGYXs58o
iGONJz7JGQgG7PNNH8vGrwEMc1g+oCB+SbK/WlEdUZdltZVa4OUtPvxw3NoFIWTv
lcMapHXnGg0OoX8D1spa4KEFqwgegbQfejvU18d5mIGVXU5rHdj4VfYAFlSzpD4h
E36R3oATy+UhOkht2sVUGEecPFp82oyyMeYmTymSptiRNPFXnDwKRVzxB264gI/J
lM4bCFoJJB0eIE4wH57oMg9ISJmW2m8yoYtjeeSKJvc9yjrGKDHHlvuLIzy+EgHo
XU0Xu3TbBFLUaFfhF9EP2TensHEYIGYFJ5o9T56Rw0fVuFiyNA+HvsfPSu7M+nrU
WOyTY9MRo/fMH8yV+ky8nGZVVErVU3l2SPO6jWYNUxYeZCO5tYpqGnhsMADlHumX
1baiKau3D9KCDNEnPLY6AXIiulc6iw3+N44Ui8aijMIuXYHp0CrKfF+QzxHxG3CP
gAfpSXLnePJOMt10aDSDAcu3oX6vfve7wT/GdJ3V75FPYCtqJBA89/hEKW1m1j5O
nb+T07QQGyCeBZ0ptq2NBqIlMVhBA0K50X2Zxb8FhQTRVkYo+DyHTosm6NovHX3G
OWvWn6sR4/hXSadYjwiPlSvaks2GRplcjYsjrXlh+5cuNXFBAucxzPjqrg0u+SNR
1oDRaZ3BLO4ciKN0LS5SM4qEalZRxyJpTgV/JfUE/R6vqP4x/orojOkyh+Joy6ZD
R8Wp3dT0nAfDgojBxun22C2sD5DTBWPxEL8JQtpKvGmUdtkRYMkTVGXyFBYW1GqE
qw2bFYWxZXTyidis9PkcdmjJyneOXo1qtPVQuu8tqV1d+3lA2Yjk6tLGMhN7CmNR
4MU86Q6L14oQhfHTU3FWTUAaXJbsoWQtJnBGlvDQ+kSPF8+bv1b2VMQ2nXAWTm65
oiAlxCQk1ZIwQwJBz9tuFA7JHvcaNTUq5HAvjGp8q5dlVsFkqiv11HCra00gUIne
u0xTMa3nw2HUUUT1e0D4NFo99cde35V5MbC5pub3tv8Smh650KBJpIT9JSh3lzNx
jSFesyWGgekRDXolKyeO10dXx1Pt1Jgf4hMDtjRTJ9/nJet/jqS7azLI1y4zWTb7
KzZowDMTTHo5WGq80pIcruvyF77AD+SlfxkIz7xVK17uKJh9TYxOanWsGhP/b7Qw
OlEczJwiKyKujIvSYPI973J2WMROwyprmZJio3nWvNWVIODfklBb0ncfF+cCtExd
4Vh/KrEQS5ssaJem7aUIhsfTmbyQPHj3TkJQFg/MuCfQKSO74tChNnyJZiSbkDr0
cjMYIdW2xeQdOQp1UhuTZub3CK1oqMf2p8CtgNWQoBWIRvBOCUtG8MNVa7djICMf
Jxd3XoVtIJawIU8rxKi7qsvAToA6SwwUDnjaon+0aqPTAmCCA03Ihoa3zI6r3sRG
EmRUaK/DbUVJ9DW4GKKs9tjQm44VS1bnkBy2Ol4oKYEkfQQBKGSDgfrsfB5Iqfl5
Min48WIRFBwhFYlA0e3BQ/0bAuHhK/GVPK/Gt5qzdMGci5+cleNqu0advsBV0alK
PGrIE5pw9pA/2pQzVgoA3/OHEoA92P/cDzXNgV/7B7iJPrP9sFv8YmPK4SRDsrm8
vgjquhKCJLvGCPuzjNyJ0HErSLRy3EF11s0jyg6LllYXdEC4NKZwiOvmfr9ou0B1
wv+bO9BZZniTSq0w37TLAEA+H5EoPKlFxpsxcVypmafag6+Xmv33tAcKczmHkwf9
I9RMkQZFxeutZyQ7DiWip1TG0IaV0MfzqnsJhOmClEs3H923nyEBTaJ6mFFJBIst
HBQ11/h8MXcgOyfUPdO0uQkzjqiG+UZTWFkOM9O3WPkfXMSOT1cWXJsrmVWihtP8
GzmMCKu3btj5aHd16TDDDUzfngkgXFoEpB2KL6WNS386fftrGtSiiaO0oRIzncpn
4LMASOppSVmdQR06SjI1Ibiq6+mYJeVUxjTNfgUzCJvrrFhMRiHS0jb1jbGgKNgZ
GtQVkwJKIR4+THJXPVOAm1klyXWkdsV4P+RSWJIpJA5PoJwxT7mhAkAIPNog/tVC
N8fy0Id6pWjBh6P0dUX2lkEhxGGth2Zy6MNpXVHkJXqjm4gexXrDB04z5b37lgQg
OqXvVqbqN9nwFAIgTUKBPVfJqJjabzJ5HRUmFGxosKuxWSQEFiSIMgtDK/r1nYNk
lCScK+lBLkm2WPp0n8hvGzTGkbRVMarn/Dt5Tzz2GIGwkuCXBWea6PGJ26Idm5A7
oHuetCc2Y+lqstmAmBURxLPebt9fqpUPoqbBByR3g0yFW41E+PtKXIRnTIjJ+gS5
kc8/TNvIJl3+PS+8qYt610+ykZM79U1pmp7TGTTbw3OkB87ouLAyaO7CJMt+K428
Oovig118guean752BB4b3PZ4uNgRMrviN32cIbUG4kDwDv0NU23N+hFc1a+7Aj+h
HcTvntUmFUpezOBGKM36zuu2Hglw6L+2t2xSUoTH77N4gSMjP8FMNOnu/4AgaiDi
rtJf33HZmqvZRQOJyhancTleAK+lU5e8vK3NIYD6hafjVLrDwJ/Sx/idIUtFkizE
irFtsIuegBDTsRHM04LwphSEM85f0CzJBnufKoNI6P2CfE6EX1PCbN6fukEMZ7d4
ThtoVmcGaHJ1+Ccsvrz6Dk2YezMczvTyIVp0l3h1hG5Y2LlHkCV4YcQ0HWbB6AlC
5UkX1w7l7ylAUjbT9ugjVy9Uct7FGHpOvxqok51jsS5us8r4gxDMp38STvGa3Qus
NajTjajDpPz+Xs9YEVt6py91txpaDCOrgN76ZieyK/S/bVU+Z3c+y/lPhLfUIryK
wMpDWkwhZnDnsx1L/igfNXOoifffRZnC7hE5qshqtCcq4z2MAOumuHyM/EwexBaT
xh9u0gwwrCJmCkzLZY+ncSnBzL1iWQhrprtb+fUAUnZiLfU6GVpXOaYMiTuhFSQD
emMl+2BS5V0qfNuSPfvXqIcl8FRbyFy5WL7nV4QoJ8VRqF0RNjQQM0JO7rQlPyh0
hamdn6D2IJQxA8V5ROKAVV3qufKVnM5I3xcoT6thX+nR0kHtTmIbMvL0wNApbxzi
1G86CLDu0rFEMjHB/hn9E865EttOWRTQPRJ4HTqJ+JmkoMJaoo0a3EBaj0hguY5T
U/1S0nYQk36vn0hIo/EabxrZUKgDBl9aRWt+eCvLlQnMKKTxRrBgDGYQKim3SQcm
HQOD1hsJ/KXYwDSibsPS4LqCucP6vCwP/X5RgccWVLCGGaFVSzq3lkEk6IC/nEqU
FuvGbXfxVy+aZTuCOLB95qjQUVti1lb9kcLnNWB357I8L3V/yTPVf/waW6+C+zTI
oz0+sib8Hu90kbKjgj6sRWytI6iLN6VYd2SBMVVjeqiuBgi3NDkjotKL3PHxqAOs
9XtHdeinc6FrRwDa9ZmVv4JZCEigtnMwwrsAjB2xvL7wicfeFIFWvt0cq3RGSUnZ
EjckiT1B93Mk/eU9rp9Jlcq+Gpnc1KLsWQx5Nr3+W5SVymw8w/t1KKDfX21zAeCF
WfUiOmffxpmZYFpmDwxezOQHSyO151V4LABAFuS4nsCoOm14fSoElGJuM1aPSJFM
QU3eefsZKBFJcfy5vkMdSBhtVeFDr5Pl287edxKwpZaV+u2ogzBdk758igcJ2ZKc
tRANGsL90AuGmmkcli0Kk7DY/AY+AUNlr/uIDaixZoHBKa7E4nkVS+IBflawLmi+
UZMfyW2JuOfJ3TS6QyePKWrJdDX2FJZWAXGc7Z+PZGLS1WWkzL6SvB2zjH0w2Tsy
Hp0SbTicoqFAkm/whrUQIudpreFmCcVZk/ZsVdaIXqIke453YHNh8k0I0QmLOxkk
KIeC52+mJyjqw1faVq2Uxgp115xDPlJUlqpmZzbf7iJnOjd7rN3HmqDtqjSIs7OH
Hc59R4nCDdCvcSKdMkQv/iqZAtQrPZIXrYFARzH0YzJqgV5Hst0x8WJ2dsauWpNV
//LXpbKt0hUXEa6CiNNqxdqRUyXhJz3WnJPj7GULeOk5Ypu8QvJiaE2BcbtXTgiB
26C3bxm5ApUsJjE8XwN6SmZDUPauzob9tLsETjbseUIaIaWwSnaVfqcTYPbeNoid
vO4oHZulw8L1/WDDqn2Od6taxLEf6Y008yHS2s1SuHwka8suiYRzuey/umbah4oX
UfF3rpUy+qNftzk3wlk6RjAVCWvvJRWTgsWX9wIzG8yNT68Wc3I5X3xY62/JyPFC
AU1ZpOSZhndnx7hw/CvIfZ8qIpNqxFALb5uECwwSoe3WV+8eGUIr3jbuR799SwdD
BbC889df09DnIs3biMuwnGaOuo4JIBBmUxgUy83KcXJbCo6L5uIQFO8vC/jrbEzF
Yw1Gh1Kq8O3W3fj4lFWpRfZbG8oVEH6ywI/OKuCmL/3ZsXcjRjF+QC3AgDcpYof9
mZC3rO54pqpy/TOXhNd0IiWxydAMePtvdSAKGJfivpILQo31FKq4HkZoXXZgOw4D
2Z57W5H/6/sBHYHuqcxt+nDpnTbjZIgC8tRFNG97iDsGfqQd1br90GMTWcD3qcU/
u3OukLH+Un7KSa6U6F2JE0n+T2E0akaFwqtJPwl7oOFYmFrO8w63b6XuMda8riY4
jtx95va/ZMl/u6s4dCUIspJ1EY6c9EWpDRO+mYS65qNqHT7MhyZzVVyoahQJ7RF3
ymo8MwuQfAxvVPPTYLHrRSpnPvQRCc3Aw8viem5HiS3A9nK2wUh9YOVrIzzmRxi6
+4UlmDCQixLE9H/XvLbRyiWEY9iYdV0fwG/I8aL+GU5rPnlMnpWSnqyOEPLFbMH2
d5PDvLZUPXOyjuSzQm2WfgtWKaW4QyXHGOnz03cfT3TQ3WrAj/ibRIaIge1zyJuC
b4gv2XrjshVchpns+TL/66A/djuQYMu4uTmCUE9bhONbKv39Ff3ycIWWC9QhVMgQ
jxCz82OCn58rlLzOJASYdqamqHSf7JKVp5N2a6WqDR4IuV6NdutHasL37kxWXOvY
m0zm1QvF1Udf/1m/DF3tnAcnhSZPqQMFVnfgnTi2H6SJ3jO/gZ2fYhiSK+2WV6xn
HtEVQNVafUFOx/HraoPfJ52paz43r/r2vx7Rjb+yfDuUvoatwU4F595EdpEGeoSS
vALmAo7a80mUaRvTJHOfNCiARY6T3ansQxGoJCo/oObTr0ypaiNKJftsVQ93RUii
wdgHKnPKOssORK2+fhEG2CpposqF33XjuRtYK/ez2IvhNDHMQBJN0QzJn06q3twC
jCVqiRcJxA2fANpEGijrAQEqH/3fZy14SUiVgmVnR63hvEe08zAVT4oGZq0nIbZr
ZaEL97EYqrmlREwR+I9HLSosBD04NT02k2dcRholY8O12+jfSxW2KzSXF0ql8HEj
Kl0rQG7636/7Ii+O8nMfzN58O7lTBAEnh946tku6GlVX+JVxg+HMy0Ru7eo2uRd2
7I7QrcwDj7cXHp+N15FwNS9Cmy+blrQg4yjdePmHl6Z2DlRrmg8h8psLjbjqVhDH
nR8B2zc9l851Vzt5hx/28L5AELg17gE2YmR6FaMY2hzxzR9lbvceoKm8/nAAKJ5i
oDFcpQjPAq+kzJswyOR3qbq1Oi4qtllXs0IGMUcU1H8Snruie+QUR3iILbpN57c7
yCtIE8Y47qgANTB/oQvM7hD8wOQQAVeUASaOhTJ8rADxrgnV76JDuAwmfbGVvH/i
KDRjP2HJgUzY9R8lJWcZzvEBLo/a0aGkkdQAfHUozbh/YqWrqyKLstP/q2GdKZD0
mdHJdD9SmcRJBCUPc6X/gl8VAG7+pWM9BeQa/b0vz3I8S703QAqW2ZINVIyAmYrq
xgKSidxP28mxrW6E6u3D/YP65THi4RiurEUCQGajMiSKhgfbJABM7AcXdX5mDJg1
4fuONPnSJyNsqXFUt0DXdxjGOqwdGP6VeFEq3qinZJZgnNrKp/sIR3PO2UKw7dTU
UgpPjATYjejx7GWbVZCLWBNTJHo0hPt2hikEA3wEHV9ZyvEEmmB05kswR2mD+f96
5wifUV1xsLjQon4jqncmhwLoCVZfwyqVvSbhvcHvAn7aQMReD7XQ887eRn1UXnRJ
d3ezZnJ/85Y4KmX1YeDw7her7rhiZQ4kjgVE7tmtgXGdmqILjH1+OBe4nI2vSL2Q
SPrJPh6qPOyl7DpIr/CyD78o/A7+Pst2AWZO0fozeUNFloV1abtbgdmj6LPdW5kZ
IR4X1flnY1n0SMOIL2xz4qO81E0L7FbIyp+seeCgg90QZNwL52WjrGK3PNcpUTyh
Ot2+5jUyMmp1hFn6adAHuWSMcyHPCD0NzARNMAeK93oShFdK/Rno8vT0+HjU+Vfd
4JilwoGoegWHqpNFwEO4J9lW0t2pAbeBCI93d4hDbkWoofkWAMrPdThmwzxvzDXA
Fb5DhmlsN07XSJyMGvt5UpLhKHywEjrNbXiWj/fX0XHMkwNNgbWK5h8MgYy9T5eI
qLBvwvBgV+12/sRm24qNcsZUWm6UnN10u3Z23wmnQz4pnM0fxUcTydQCjeDseCaO
GBVccqIQ4VmxiT6kiR0bpmK+ESLki7IV7Ma5nFcAPsHnicUeH7tqSCJ9NU9YVfjV
8oWg1ljCNf7YY0gcdQDAIjbSOqBgOEk4hhPo1Iw6gt2U8oY8e9go1d9qPGuWuRWV
F2TU0byim4/wlRkZFxlM2X/2hfqUCd1dbPFc6LTJe1HzDizPXiCMtwNSqwWfNJyx
cS/jDfr5/08X4DnTRbtHMPx86yYCN9m8IFkUOr9/WebB1z/usmknDCKNsH2iLeMI
QNSmtw4UpQa9vJpSd31Ygfs1IPnu0yzRa/EFy4TOqctB1KSkiEp8SdnxYnIiyUmm
9m64IfQ0Oqc4XGyMQotk2OeHE0chV/xsb9y3kcePoyedxI3MNe7YEgfmCW2Qz31V
UhNAgB/PaEC3WwjUk7GOPZuZcmbIb+65fkyi0iGovfeAxNhjvn6Y7CYD/VZPDq6U
j1QcUes1Cxv9CFTRd8dY4Yhi7Ivl6GdA+JchQgEu5EESWxEBGXVHI1Os+sfPt5oY
ylHb2ICN71g5Z6tJSJHacTUD+G8rxlLWcuy0VnSvWOsGB9SSmXpm1XbsDieRAJwc
TYRu5FzOrvkfk/P6H3qbPAcNWIKJphJNlM+rv3UbVj5JklTSJF1bSxbd9w3CoI3g
7IO2u05rRIqGcosF7n94S5FiunL8xORtRaMfOStSodKUTyZTG3H49A3ebDFZSt17
0vmxpbUEcySfBLy4tWyXZZIXbXEvUiOTqpVmd1MIMe5coQCEfPsAqhmf8PFcWdXw
XXuFLFe/QJqgJCbjjSqQC8hfbCIzjWqaNfWKWk/s1aNd2RNKIzTvOr1nlBUXwvOt
g01Uwb+enw5TUXtmgYxLqVOrXdNNvEFF51A+B9slzlqidEdSVsH2WPr3HY9+zwll
EGB/KReeIBqUPR7tQAhty31u8gcb8woKS08Voc2ygLcFwyGDWT6AVzihcftwxunq
H9jaW5MZa4OeVrt1FsX9MFq9IGOntmcAQddhH9G7A8xDVa6U1Mgyp9GLJp/0X/lZ
5edObVIj1RO9GVQRbhij6R/guqOKzy3Gw+m69grhx6oerZ0TJNg6zzRUzz/VCp2r
NnqUvQOX9pxBhyy7Gz/6+x9V7sWPKSMN63JI40CV2TmiR2D0+sa9iINAk1SZ4Qvo
sx/59TgoTYLdslDYjgG3q3bsVGdBehckh9XXiqGHzquUaOozZEj1fU83Clebz/FP
i537jCYDHse/swxanFG2AtA21d6zPGrp8R2eyPQO8NajicqE+UCmUFU2R4Klb86k
62WXCZo2y2NvyWcQX1uY/fmEGHTlexBvTJjkGEV8CIxDUFQSPNIOZ4fcvbqHO9F6
OTlsJhuFvqyuZOKuhHaP/QzFEMaXBogjEFk40i+Tb53S/AkUvzLOcfO06fS2jbtY
JhfZMdvNJD3PnomqZtUQqOHrlp8LEjV3NMXd6tTgGBnIh7oHnXa4DbnzJYgMX0xp
mVv4ntBilCFR7ipzm5YmXjwQNfQDy+VjkVNeQg83567kB6T7yoGj4Aqrj7e1uMPE
qI6SgSC1Fe6N747Q1u6Dx3+Pib1qgfcApKvikjXPMMscK358r1np4Tja6NRFKvCK
V47/NQ3GuBGNKs7UGlc/MimkRwDmmJk8AsVsn9MYwhWDGyeiwJUGSNvsfYdR6+ve
9YVZjNV6QRpoHizHCaqxHANffvdCVbGiVxZZxheakq7r+OZq/DSNhu4e6exTd8jF
EcF0icKKYOJMcv1A+PL84oRTo5v8RvXWa4BJwb+DLQ2Y9mg4juidBT69g3rsPYQG
co1fIXMDRekUNQEpzbLoaR5wYSylO+4L6exrisNQOdDQHgM0qLJJ1ZyBXaPc+/K+
qaN8470Pg3L9GDLEM8lhh6IjHOy2q8yV42PBIucwXVr9mFQPvi/qXhgaCM63cM3j
lbVXfgzgIFJx3kvqoCTnkAZ9ZUlOxEsdFhCmQZs3h8ZIKECyBZsGLIZY9GXRCkoq
HeoMUVuqwf5jknqoIPYQb1vnhryAmUKOqX50E/H/P6s17IAUqGq/eAwywwPwD2bJ
D+gU1GfqurfbMiqIxYxIRhRzGr3g+EIjMgvKoSOTn523234/t5RP6NrCdc2Q4QE7
bU+mK3PAnouo9cA/Z3/jRFnPtbGfoaURmr+1OChDDfr/QBq+PHwemZAgeUhn3GyE
sGr22e/dpoloEutwjLI9ga4ssJyTXL9RgpE34UyJeJLPcBWJxaGp4PzclpmqHFVO
yT1oK7PF04XlVbD2TEJZZslNM3d6Ji9+A7pil1OrtPkTLVxKmNH37yqADe2rsUag
DNlHHsgzQvl+EGvXL7bf8a6RqHoFZLOMd2Vi5bGcf91AUAcsbylhxnMfmFg2iZlJ
wNsc5frael5OQj9ialVqgIRSqWI7mJTXgPrR76I4X+4uE18ClJgLRBxXRk7LoS1y
9hv2pWb11LR4Iseuyi5F90xPLlud1QrSv3YKzR1DDF/4txlrm5YUZFhxN7Obp88n
0f/94Axcg1R1PKo/r8MzR3kgy7tgy48RdzoxftB4KA57QofAbYeyGy8oPYQuTzuY
Nlb4Jo/6zpw6ADF8khEvIx8+DUwZ17oj9XtU7SPXZ1sleO+LsdqAl4A3d8ow3RMv
6uqxA3onvwRos8LCdJqm6/ACMo5KtxJo627sUC/WgJ6aqOlTanRv5zj9DiEBZZpn
MeRVzWd0uG+LBwLgPBHl6xlmTbD5Y38Ceg/NzeDUsctU+sRPayRj1zaHtviS3For
TFEXdgAGXUO22BzS4gDZ59rIQnxZHjzY7JkXR6NDnEZ+/JHrRYwcFbcsVgDH3Oi8
QTdH+91Yk+xvfkPDJL4DfTTm+i/VRRRkHsWAdaHL5R1KIVbrR27neloEvVEjriyw
2mQMxlLe/4zzD8JF+pzQjryKBIg7jXjPIJU1FcbuI26GG6W6zJA66kRZDhS5A7UD
++AQqdfGuLoJ7rmfHb6Ozet4Kus8uKgd0O9lL0jMhx2/0Dr+n5XCHF2N73m3Hv0f
45Z95tWuCe3wL4S+I/r6b0a4f3b5TRBt3EKCKAu+KbNy9GC21Kc2S6Wy7e2QP5vw
AWWfiU/Hk/885kTjonUPEcIQvGwQppbL5mY611tK//uTpCtvZRKeWvAon/1ntre2
cnfEpup43uzjaaKPxoqtNYIoDXVJ3l70O35qlpxc/HmuragEQSdEVm/RBzmv3CtD
d1vehMZbNImZ525VM0Wah0sg+bJ1MrSD3u2ObGmw/59znHgRwf4mciHtvGe5Q2Km
7kbpIcQu9oOw29p0zULjUAod7h3DZq3TJaESqEvrY29MeL2RzGFAk5H20aUJpAhc
0w3ThbcLGMXzgMiIRXa4ZKGEQWHjmlBT4wfPhNcbiCnbgcGcryJ0dnYjx+w9BcM4
z7EmkNljjLnSNGaaDm67LvoqAsKBENMH+uiR56JChYVMMyV7Qr0yvrZolhJO1o1W
GCIPKvB3WLLPc/o9GzZxKUs3HbsyD6flO/spMwyemFCQZZlteCHNLFdT/jchU9UI
oo4mngZSekLsE/hplQydXN4msXOvE7+fVJ/7ICsedmKjOlg5zzpqhOCLvMc8pMA4
OHC+MKCZ0JnBX//lKnfpZLv8xzhk7c4GEhWS7P+Pno80ahU+DghNZt9TUzaG4qD7
diqmjsxiAXZOHZFXLJl0YVjpP8R6vcUUwg+ZCdoTHcpqlHpdbzE2TrdcL5ik7MZE
DUXKbllHeptLGmrndhE0ywuxEMA+qOfnWp6rZ7mnGShuyXgh8PjNZhgrtTaNOXQL
4i+JREHYBU1jaKlTAAnqbt2l3fjRxlmtb0MxR10Cub4CnzGiHvcXsK5CSDefVbIA
b96RHu7FHD567R4CuarX+NPTCIkP+M6wyXuc/2uEJh6gjO41Lw2sHaevfgMJhN8N
AmXt0EVteuXsLWGxO3R1L4CNBSz37RjiOq7uJKM7ndg/K5sRSzvyqWSg7K0ZYGx6
cpLQ6BW53VY8l4OdEAiKyp/4mXMQU/IpWV06JSX/RQ3eUYoc6imtPNGcLf/NkSCZ
cXyecOGn6XnFbwx2F/r8lMmOY+D0g/fmsP3aV9oZc7oSX7wo/ssrGTpfQ95hkSU5
6kYLMNOTCJP4X2GBhn9dcva3amSX6QuxCBcR8lQvLuicdf3YguyaYUUBzEFKVUs1
TqWfHP8hESyRuO/A2lBzbl4syWqzjHMEm0p/sf0RlNvxh/p0oUOx+/x5gPJKCcZG
ElG7kPjJORW/OifujG0zMwhkmjewDVWZuq/yiM+lKj2ifTnTfzm3OLbscSQts7h5
ITteF8bGgiPJ6hk4HSBpIvHE+LO6aUNQnkMh3Tk+Tilfc2ZM0pc2NRddNQJzVflx
pRYAB+3vVG4wtTCBlPNmCPHctE8iqMhoYGU0Ielf9D0D8cSbYNhk9lFmQrHyZHMW
OuASvnazmzv8jbCffVNdWxPlvn2KN4KSy2F4y2i/nXkgn/awGDVH/lKqBpuLg3g4
Ai4CW5n679tLCGr/eWagMEbSuxWAv32yCZnrR6ROzYDmZI+GJsBAAA3c35VBohnX
1uLcA3qLgX7ArwWbX9M5IMqBnynee1x7UREb9nlkzikKUld+P3b4/MNnO+Yu7eWW
efOzX4F/7S2iZit7nqpXAq4oXZALtbN8ukXgn7t4jBEfxz7uedhVTO7M5KiLYTpP
73LcWJ3ai0+GxC+79ZTxKOehxmR9Q1N5s6ApdcWJJrI=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
vWaiee8LnCgatAmbQJm76HQ91KPok9U75lW9XkT4Zyht59IEvmW+9ocswzwHHUoA
+dvnB2vZ3UzRuKae/Xl6XwEyWqTsK97Y91lTDvN48S1bEBITV0qTgwl6P5pXZ+wf
HXawhpfc6BneMrHuJXWCBGqpErR4FElMLcxuqjxP2WYmbsOBlgl7hwl5F9ZwBLaR
kzPEEFKYAE+PbpdHKA3AZsuAyMsyhUjbyi0LXNKbwgvDMTq6SoQbsLYb8I+uZ1yS
jcJySo0AfhacOg4lpzYXIHcW0VFt50/N2KmZqXbQVG9/7g6EMtty+8LKcqi9D6za
hH0oAOVa2spn3R+N55wPKN9S69JZzcBtfIB/EmtvQExzn/sPHwr77N2HkbTOY74l
E+zgy8XfpBT9fQGvbBYImC3WoBg36qF3zFmiNnD7lYiD92tXF/F4+ODbUqdTpi+h
Rbhsjj5KoYd8LgSoliCd9/QZF/6koT0na5NTdB6NXWz8D5TUEZQQU/qRHkvVgG6K
1LbFnSAEV7HqahJcLfCJ93No8aYTIqcJEbJqLfZKO4j/kV1uKH9MKTaGPe/125Z6
aw2tKAPPB4A9kIQQdcBzpOrc22kjhANFNHP0P2kV6BC0zWrdU+/sKd3YqT3hU6GR
TGEl8YIMp3sNV4mut7SOE0YUkCHw8p9/dadSsvVLomiNi8mq0rzwcacY9ynoo8vK
gRf7GCK5EaMw01F3dYDaUP1cuX4OXs9Bxq45ZGVDPfEoD0Y71SL2FzFTKIcar7YP
Fh3n6L++kcuzD6UdEfriXk+R/PL8YpJeSms2L3fRaQqWD9uI5zyXT9uBQvQEHsbe
b8z4vlu9yb9XXReTNFgKWp6yDfhyNgpDMgMGw0kiFVaan1ErxSDDegWFNRzDDUMQ
53xSEjBTuv7yHY7uwZULo6TXfIXV6vmxGj4jluAstqnPeQcWDPSg2S/iabsjgYvo
t8mf1CU/FdG5MQDWGHD1OuTMzXJ2NP++vtcT/8E85yqfoAV5Sbw6LFIllChmup/X
NH3sW7PuXhwxC0bKWhJvffFERmwVpf+sw2saMkpO4TgfXD6RPmwrDtnGDul9BIGG
GHrHybVWbgU25FryczbM1+XpX9bsM+aj/X94hdlU667UD9yNRuBqXIxNxswRUXav
uVO/q9A61I1e72Dq9mezMbl/Cu8fH5Hom1Fvl0v14LNEhuTfk9uWIOLXSAtiEBQH
1xDMm6H6x1K4iMhZLtnTsy784bsfXOLhK9wlp3cvm3xM+DKC+Sal4vhvUvd7xioJ
W+89zsiAMxUYxDBpsWycW/QML7nXx2hK+WsW4+qu1N+ILNIS2HfCkUz3SCfvYYnO
jjBU0JcpTNhFf9bjx8uJgZSwPURjwEMrZRQLP2vEQsgAIjdCh0PxkgBrNROM7kUb
jcjcQPGvIwbFtzccfGr21aTmxxhVCf0ztsnycskwNlBXFseYAUZzIOFpl+Gtti5k
Yt8WosIMF2RHX02OedjkuwW7uTGEftDBBeqXmSJ2AS3iHgiVu8ejmpT3RQ1DWWDy
tmJu8BfzOvBZ0iprbXQthK5JuD3L5NzlYAfQonAICq9QKXW6y4r5V6uq3epencEg
sVAowoA5NwZZasFiRf3TH701Yzdz6fAzHg55Med0AHFIEuHQHVvwUhSo2rdYKOvT
sMFZrrfImNCDQZj82sWqcry/wkEo9jEl1HwzkSQSfwmtAaCNalq6cBgJQilbkV6k
uhoKfiB7N1kWYHcsbegatFvMTBzB46pQZmhNnUAf2hyhDmQMJaiCqF19y+U+Mmgu
PQTl5JZGWCsg3k3xhfTUz7G/4rnjsCwSTGswTK2WeuhbiE6AxkAuAo3gJosOxoru
61JOUPa7iPzvO8XIZ1ACrrUdQ7EwLXdwewYUaIFa2I8AsxZNMLY4ETsLowinMAe1
g5jVCMf9KZdE9ZdHzYAKGKYMuEcbHjAEJ+eqQIV1b4ynlPw9gZ1ehUoQupjOQnyZ
13TcKfZRNDBrWAESTsn++C1ZK1cx2crBPLLo8ZyAwKvilDwUeOc1Ux/91toBUI0P
s2swdFnuYy9SgkIvH4H355dkP0Vwf+AmsPyypXPJDrTdTL0F75bIkC+SLDvMz15X
1un+XwC+HfUYe9KEJtD+OWS0NwUr83hdRUhMrpwnTiUFMRhoeveRLXMM+PROw/VT
pTMtuGkkgzGnoIBFcuNG4b8jsDhz4CcWqEL9EiE+PrOCmDDyRvSj3p3jvjp+zCA0
m5+PjeI7cnD0j4xhE6sBC4QiyAlajkoEQ6CPhvOPRcDpKne3qF5mI3EoBQoyU5SB
Loy68eV1sg44J3gPxeRe+1ISd9phf+BRCU8v2oLzCw99YTRaXWRYZ6k2JSTMaxMq
2Fpd+ma9Ug+HtfcBDT3nBkpn+6ZWd6QBqqBZGF/dojU66joJF8bESDXWvSKK4PWE
OtlNl5SSabcSTajMv1HsOouQrEyZ8DUZrrfw3seu9JfViyEuNkUooiGC8RYhmmJM
w8lpPacTVRiCvSoSmAE7oid6sqHQ5EwBf2rRWEb38LBI6Hl/IIWgSIDFFKXIwMU+
YpDoMA0myoCHUQixAUEut8EOR4s5njb/Q9oi+ewrp7BUAODhbBFw/plmcn7BI/yi
3XIry9gfk6zY0S1Lcy9Z7mvfvMzPV024CD1OgD5dvFa2xD9PMXt/Z3SuBLps3/Ng
sWyzwuTInaVJErNAd+ZASCef1lN/jUYhjf7Xd+8k9X1VJZOKk3Bikx/F+HIsjcwj
yUBkuaGpSAMj0JilWnzwCE9p85mcZCYG2FA41FhkCWiGbPiquyyed60X0CXpG81B
nI6JNm2I3ngb8HTcRWHwtS86RFVh9q/6MQdoXEjnWCK5JmEqOy46xzqozFKycN1G
DQ6r5yCYe/WEXYzG9dpsZHF1AyVh2wfzkcB7tWtlmykm/+FR2Lev3h4i/nNtxtlD
yQfSgeFE2OPSa7Ts2xnsGy2YaKBR+rNaG1CEbv7pV9tjCwuDxGrJJVkKRAVA/IfU
NGxQ08LwBInLUY7VRx45asuZ1NoT+vVNArZZf3M5g70DhWTW8xWmf/ua8Bx4GWxD
vK2HC36GxrbGDXXYeu7LcwT+PsIB/goVkZtIVMwiTujhI3igwER1epEOaS/CjqnU
xju9Q2geEz2pyWM8jiXdl9YlJmpL9OuK+CP7Cj0wAzfbcRmbU9WkM9LzDlwd0EY2
+RnPt6HWxyD8ALTFhvn3v/JAnQgS53vstqTjI/wl3xDYUlR0UoorAjUJQkzZzl81
0ypYdt9Qkp5uJ2ZlP9L6dap12Hz4sT6q9DAlQREDIFl8pz03bJkEcBqSDgO9NzJQ
bRdttRuEw6SNc64rOWhQb+u3/BemizkZoTjFYMxwhB1q/ZiYtucg9SsVHsmuCyL2
Oif5b9cgBJWpe7oji0F3sv5DVK9pXWXgKGLuRWtAQgnaOnRya/7vYtkg0dIVt5h8
lqFtOHDPeyYf8Zv7t5JWdjCwctzm0Tn0Y7HuNsFbtaFd6vSXBbso6eY5WzRKGX6r
98/8/8wa3TsFMKqXdLYQ7FpzpgmL+nrqrum+Dq8r24LiG2/XM5n+lQiF/8psJwJ6
xuWZMiTQMQQnJBPlfa69vLiyuT9C37dp2QYGBWOBOUYQlhql5209ZZBV46WtAd9O
nBbqPdwnPFOJLs+WSVokAu+R58JdVzZvHTVyihpNMr8IugC4IuPpUsX1+bb4byRo
rqi8NW17tc1zzNWdD3pnkcbmb4O+qcsb7gb53QjDRrAlbQnwDWxV7ovgwnrF4sJW
BAoaPHZvwgzwszz2rcWy0naR1TVdiE9OhRKvJEhwKI/WNIFdwLnVM/c5xNEoeMqv
13oIZg7kuiPDFhosKOhlXNC0+KZIvOTFUJeMlZ/p03mxFGByW9Q4XXRVKTp0Ez+2
n5NXEKB6zGKuhpPxiaz5J0l3TRnIIYNHYAeF0iB3kTCbt21SILZ3e7EuSCVgN/bP
dgLCVClbTttRngclv1Z/75jclrI68Ea86L8X1ld5TiMIyTvnCoWuBTJmssm5vL3+
3ZHr+du2S/E0ghSDjZRKuKPzEtoHFBATYGXlIIAB6HZ9UoE1/KuPch3H+X6zPB0e
3yzRTe73lJ/MifGqSp0YlLXbHUeuxj896M006wjNib0yr0NYVM0zzrAiyObn4uwM
h4fmnWivYV//6yz+lo5QgJi4NiJ1CkbJevRmglBRSbhQkRF8Ve3q/wUgThl6QuyJ
w2Abx/FRdTRQhJpvIDvyMknsDbAQE0MIP8bBLX+8rSjTlSa+8rfZzmryqm99Trit
cX8ErsXHdbW+UziWmL48NYYdkE2WPrrLJ8SqxC5ZEg8K0liJgKA3y5CQm5Q9WhtK
5BpYFVMJQhXCmBldDhceYWCg6gTXRniTXtSJmZvQo2uG/CeKZUqrk8d4Ue/0pFEl
5y6xZnyHtBpxpYYfPe2NI1Liit2NvL4nczYbcAOWtFEpMrutqQc0A4h8TeVCvAG6
AsfGqHdKQI5p3OHNeRRASDOeJv0OjZYyk4a4zrVsMsgAm3whAZpH34Mod4PPYzWd
7wkIhuUvdZitGmfFfXJrACCTesqWrbT6PWipSU4DxOxdHTSFZmatjpue4fHiA2If
CBUwuyyjS0OmsYJfFgIub21vSh/h2mgIz3J2/Zc7lGrK9fKsHM+etaDAZ6JATqOK
mFNyNog2zZ0uSxOcu5JWDThxCsTLHjCUuqSJQjPtBuYbbcYa3NOOcBQAMsE9vCwL
X4Qu2ysVnGCWciHo2guIhV3u6zTZV+XAl4tNCHwyiADKv2zuTW6iczoxkwN9DjJm
8waHHV7mhku5MiCG9vyNBv1UsXIA42piFe7WvR/BVstKqNSdqkZKqmBuKXBKPmCr
AgO6rFI5xPxGhReeV9MFCblb9OwMj4U/l1keyfzfhQ5ubpbdbjbx5xRgtbD23+vi
6KBHcOho+Bpn3S5/K5sSqSsbYK5b9TQP5kKlgPLNDC7lu7g/1SgFBfZ0kckVIRs7
54K/a0Tj3ABqmE7NUq91j4d5qazEtytMWXXgRjbbJaKijN/lSlmWHrf40CmRShv/
iIo1kJmWZrxpmS08T7ePhu+TsrauU1mcpOpkv7oobHnAZBjFpBpdmpmkugWGB+h3
1gKZ6GEsta9h8OS6n6dRNfphRJOIc8fI3YGstIQBIcs91+YASPYsFUMG089y1KEF
QYWr+6oeNxSSR5D3f3ZsQ2Sd6ILUd9SpGzSQJ+0VMfLiFeLuzetp2VO5imIzmts3
859lW5XF4kJRHjpLR3/T8W4KgL8zBkfycBDdpZdh8YvVs/GRTRNCwylZMY8kqPmZ
orOPRDyPvAczJ4aSTyFQpi3x3gdo28Dp3wdhyZMzAlhapt5X/JAQ4BhB2EIBAnOd
WVnDi1qwBBBUS9xbsKFTwzMn4rzNj24A2AN61DulVOzrAHhvnMGf9zUm5vjCLde6
2sV0mmVo0m5XyeGj4Dzdvr53VsfCruPdgtgNESF14R3Vv1IY8N8/dW589HMEO04c
5FkYk37avIL7ZLCyfoDEQoMlt8tjwUZsOAba3+zQGaXSDJrU9ACqoUyOaKgk5w5/
rpgAa/Rd9sAQKJphIlZHdvGDqoV6LjXCYZMXheeKUNtCkg17vqRczb4CIGsqfe/y
R+aCujLyO6seXAaSBOHhAUgMNoeWCGZDPwS6y29EKQtBeawEMMKPhBwjyibWaEJ2
UmmUmg52bSW6YD4r8TWnLzfEO3YvSKS6cSUiEyLBBL9H4d98tXm7XmqoEzVWx3Qy
Rv2ip58P+m/UhI//ciTGLUunuF0gHTWA8DSbWdb4TZMpn7WDdQKqQ3SPkaY0C66f
KfHSKX7FaulsWEL5R4FUEhb9k8mZZlZylvpq0+9FKVyNfaCv/RZG3jXuLe2RlAHd
IbAVkRhxmf7R8bvU6iV0Uaa68kGCX/qfEQA5tpOgGonZYEFAqfmkt1vijcHLmNaU
2LPIEnoXfi2UgqxpkdFNPLxfifK2m8PZ1l/RZiyXtWcxxZCo9rkrbihy6Twqo067
CmuTBqHtXwrtMDkHNwoR1EgXQMpy6O9FCQ1swqovNBuXBCOBukzSxlKBuI0jg/84
4L1Qy90BDq2v8v7OiD6tpXyJGWx1we2KF8HR3T7py8oJ/NeXHcGwWHDdbZl/l+bX
8+DoKTTyCN4gFPgFU3IqZPb1P0k6+Iw0VVtjUSRtypxDu2Xx36GlFrwshTtumI9Z
Y5fW39UwGf/cA0DqS+tzp6ZUnDhLN98WApMem9SraznicA6JfSJ4y8DP/0of2LG/
pnOCZ873YFFQ4HuKVoWXOLXjYX0YeSIedoK7JAGUeeJzBm95+DPXGa4idqWSqRQ3
ZZa3z3+otbCIHYiTeNSL47eiIlzFG6V2sUqZqIQMZg931cP+Ews5P7mu1e+91o4x
/z4GE364WqGKyoE1zpKLO0EhP4kLIJ/Q7U7/W6TE+9Ixvp6+8r25TsZDlo7fbDR5
0gIRK8DjyhaB0B1eO2ruVdRMYVu0ma9hFPqKk3CQ/goBIuK+FMLy7Wa1f4MP9ikL
4BicHudU0RwfwAUvbmw33ZxpcHxFQzllsL9exDVN7pniT2weI8UUxx7aEO7Gegz0
3cEiW4lq8MhUMGceZe5UD+GI78UGDeBMUfzAP+594thtOVxf3cOFezgVhovUhGym
eF7mqbX0sWAgW53ZY2QjlZZ++93NX3hlgXlVy3LXs7sKtkAz2jp1iMPGWmADXWEy
Xd7KX9hhBJ1Hyc2PgXrkP9VRVYlQ+eeAE1B0qcpn2F8/UhI9pcMx2TG1H5ymprjH
OP6xnsS0Nzs7/egkddMqksVKW4FYk15GL6d3y1tON899Oz4qYhSwL/0G7e0s8CzK
rKnyOE3lPv9a9UoOY/pMFsl2qXBmhh0cQKf0dZHdUGR6+l5+m6sXMOjy1UU4MG9i
rS3GCiRDdmB8pQvEKMGMDNfF6g9OUxn1NioQuco0Seu6HJHmYfNK4net8YMJHmZ5
amsUffOl6MNt9xiJ7x0EREFhbFaA13VDtgAtx73w868Bv9JAKwmYWncB9lkFebaZ
Uv2bIAip+dIpf82qmNqOe/1zgjv1hwHezRjHtotz2XbNiFHGXvC0IkR5KUW4/3Q4
kfGf1ivtTUF+cT1ZWELdxNITIyhJhGTL6y2/4um2qac0IKuXYJqCKfEXAMtDP6Yn
q/kNSt2jNAug7t7BOjDt+nL+9FrCFs0nQAl72tdHjYKXMNEHBwGvz+Pg52m2gcVV
UO8yTUT97VZl5UFS5Y0zZYeQ7XBYz0+STvSZMUzYIt9Trvh/38AYsazM2m3pNNHp
xQubRF1XrX5fpNIWTSyFvQODxzcUFuVb30OqwynLBrsAk6vQrhAlgdZ18v7uptru
o0b+8ZWsEhTf58/My0gy1AYK13fYmfON3CHi0UxiFNBAjYeN5x6UCOnSdK99SOjv
TgI1phaxxRomADOwtT8kbL7q8YefyQGmKLqROMEJzFvsGHbWDCf9yvnvh7GgDAIY
PGrYESvQbwt280JiloOlHci9+3CubuXClnn+Z13wxklRA4LuqMcw3BWskD3Kl2VH
kGHwPEsRJ3uG1EUZ7Oy3uPTEkZs7OaXp/Wjh54FSeJcIzf+Lhic6o/a3E+PMDfyl
yjOcfmvoypjnjIoVDfrK9pNVi70jI181kp614ZM+A/1dBfFucg48OQoq7nBjZVav
GP31uLxAxBm7wThEaElRrowWHkDpp7NKUz/p97/rzHfwA65eT7ZaoYqb2H2Ei17V
T0Cpl4Oc8Tb64qMVsxJSssPyAlDpl/xcDRwgtEGy5dBnuQkNjJHpH5RUuikZYx4D
V+QkNc+kzxhWqRVV/evD1udvUMImX24ay4FKagueygO3SFV6b0YSEkPKY9OkngBm
Ajx70AZgU0gLY9h7kKxHREpi27M3SK7oHlg0Bb974y28lm1npZ/WBGL8yEOoikD1
YnRWQlfaJj9aS5JTRdvtdrENjOcSYX50CWHWxq3vXfj29jgix/F43nzcAcM2ieXE
dUIz3EdCpOb32xj1OqKuCqtCqo3AXFUsviq1zPlC1Nzryv6SA29WcJ6c+4CTzTNm
AM/kueNXcEfBsCqHKlzU5FUjjBdap241gCNJsk6EBNYh76eMbh7h4crjJ+LdWZyZ
Yb9FTBCTga199sMa6sCTNvLKhGejccW0RQqKd4t5GZ1/vXrjgBc5ura4L99eIKfc
r65wxTkT1Fu+pO5ywI+Pb+w0TFI4+2i00lFSSBq1xXvIFwBMwmWvM3ORg4X39453
hp3SXM2lrt0km+9so5lWH5rt7Xo2TNg7nzNirv6FlGZ9/+QJY/ptkuoYhWa5WMWp
RsjkSPTMQZIAvyEhHALLgwl1y8F3SqFiieFIaBw1mGDlwMM3FIBEStRkcvO6DCbe
/gqHSxRbr1uEGI/ljV0RSeLN97XLK3Ee8G5mp0f8tISd7KPKD8j19OQNkcxAZeL8
v2fBsOCQtD3TzcaBte1f+enoHl/qzIn97iuU2LT+xJ+jnPJFPi7/nKVLW/yR9o2s
fD2x2DOa5xn1zc4/TVXHuQUHjuQJktV9NwPxNLvURvmrZs4W+lmAj28UUGke+QvQ
VXHr6mL1RDkY6NKFBZaoVKx0SnmQYgNDPU8nbqGrzoUdS9lApetjgBEnOPpe/1Tz
mqKlqKsz7QPR5B277b5q17xblSeGT/HTsthNMSzb0BQizHdlo+PQ9yHtcyJZyq/m
d+/GKeltzvyX1H0S6XtI7Eq5OD/McKXy9AgYCnTuxC9An+/F+u2mQZbVM22L20cl
HPLdmnNVKwnSS5ft6dW0wwYxpDcuP/7FJcwkaO/u3y6vFR2I1ALV1IxN67izjhGg
xNbGL/Af4q0uTl7HQuFfjmJAQQ8TgJeE/iebmZECjA8bOO99uCV7InZWeWR2Kl+v
OlUqkB9ZuRK8KTP+zYvT5GebWVtUa//ZpORKXA8EH5knxqei0BCImop5msI/RzdP
f0d06ne/qHdwJuml3GzP6MFcXCpLm4oUfBvxuZT/MEbg1ttybPHFhuaE1TRwzdBU
l7HUYAtvK57D2M6QBE/3qMu2SgQ2zyt0Isz9u5O63OsGSH3gG3PmeC9EQ3rEIV7R
xfiB33vahQod3b+PXzkyqxxig/czL1HPpYanZRuF0fA6AkeXl2XJZ/4T1SVCWBBE
Ityz2vxWlpqh71Mr1c4NNNfA+LxqlwLUORhKbe0HnBDk36v0EJNAdrtkW0CRjSrc
IPB3wMLln68yU1ZeKykAaX4UNV/9RBXLOSZrFWVXt7p5UiitTAp6RPUv/BbKW0Zf
SLEJ62g8if6eIuZqXlYT8EdnBFQPLL6YLidovTjikaLJzBJ4rENcfF4b1qlYYoTO
dcGziAV04TPDKQNFb7BmGk32FYxSDI/nCanwBrLAohEifWtXgZ4v+rqG6l8aW6y+
VRCU2Fd4AYjDmxn3wBnjU/Rrcq+bAkMp6bsN+f5giGIopAY1GegG9SlmTyxJBNe/
pPKMrgt+e6I0+4oQSxwCWi7YGvgPm0pgnU8haL0f033s7sHqCR//SEXDVil8GVdO
tMJKhIOSBDZ0lyDys+ubnfzySFHfjzvYNaHbRjHZDNe6MtobYCzW9RWo8odaAmzx
YPgBkF4vc55qvvcH7j5VM/GWhcbbhJhjaUTy1XwHuGOiFAGrrFc1HP/qopzAKpQ9
hrOj0Z0eC2yAIvI3HEMEpdVyTncZRO1Ku7TIIOE6FI6goLDbLePqNxsTY6KL6jaW
emUARNoPpBRjR8+Q0CT7Iu0s54vt95+4Fyz8gdWX2udOn5Lh5Ta83QZBWbv+JiYj
M2mNWXkkUxJq6W3uzN2GGqOAbPuY01Z4UnVWvrQPWr1OcHwtDIpNQN5vgg3LpXSW
duyt9P+YYa19jkBvnXaMILOEHxj7Y6YNosbJi4MY8srljiPVJ73n11OrY7Z44+/k
nR78ODuATHjPH9/wYhUnunsjkT2Tn+15RCrn4P89lNW9H9aIRgOY5gFx5cTDQzPG
G6e/y7Nrbv+9Mxpz9vJH2U7t1I0M/GGPLsoVBRlD15C8ZHlOUsPmFfYIWHZBR9rg
5/sK1l2UZR9jHgvDqusSI3oSoscpb1R4LoRomgt10E+SIymyDX/OaMhfWBvnmwAi
1PgoSZ6kyuGMKg/x8L+CrlEPfmrR/0OXU7Y4akUg1b+t9iamRVpyPDvcIbC8MW+H
qIpVZ3rUmE8XMd/VUN5blxGB/jLHLHV/Y7UPNg+5i6dceA95ezNUlbZ0cIVZHtTM
snnTMIN6CYHVH0YPLewd3Q0Px5/5MUhZMgNdUmMnBYK26jd/78YdEPqRkPG1ApMl
TgeYcItA8AM0n56HpeEo+xRZPEh1yoomzjic9A9pOFeOPWg/Q/ykdhg+Do4ly14W
ACbqMlZUp/1zGtJ16BdJEOkRQzNUNhLLXgTTQKqpMzsVfz9D2Xm4wQaCMPIrqK3t
qUyGxbFT5zdzcc5cSD3Xe/YXcETyoaRnnt5f70uwaYh9pey437SosH8T2POlq/oI
WeOuOdspIFK/bnboGtPpnUqkezk/06RVm/uqM7o4p0MLrCD3OSg20sTAnbYUsK3J
Sd3ezzE19ujHWXRMQF2Wk0CSFvA+TsytefNKeAM9iHRYMT5budahD6MzzqRyj+gY
d8tV5n+Jco5TO3lMM78pZZl0sxm/jz2Mkd85p9qsXIwjK8cogbM/CQ8tb0P5xcUK
R09d0taDQO6QsXS/Syk64Ipl4ofrBp5C3nfsj2E5E48dtsxL5mfx4MqwaingFXS9
yWHrJc55nXpVnhoYcmL2MvTFFSuq4DAvUYgJ6PGjxLo6zn7nTHVxDEjzH5z+Zpd5
EaDR6GipPTkUYuCPQ5+QpNW4qLe/lDOzOArjXrVaRrP+uH+F3Ga0B90l1daN3Aw7
1qwM4Sj5TZscqAlEya3pkZ/8sSbRyU0fkUvr0iTaqdHqOJ/LCQtIZRJE4OZwgwOK
lUgF72u0xl9h7YE96kwGiVlGGORToE10OwJrOV2ht81zCNe7P4hwN7e5CI/IB1+C
OE9Z4b+MaR8fw0GeEPJezaKVOlCEj88Bj0C64DgtZO/sAx8F6Fp7tPcAO8HYhlT8
N2GZ3NJ7zW04r+vvy34E74TVN8klBFFUl4pgA8GmKSx4pieerrrHtYKG5w0hwPUZ
bIC4EEVDQzy5yyWJc0px4DwsscDTxDZbGFFZXcP2MicMCervm1UWVbxj4VBWE9pq
9jiDFWpAjVf6AHHGIsiZbjrrWyKeRHMtJb7miMVT2oy31JxJknGdRCMcJ1bYtXP+
RF68yMiMg+lFNs9Ca6uE0IsX5ybza+rWVYktgTlZYWUNQux+KhSW2YnPCUp3dSwA
7PQnLI3iIxHq2vlydr1SdBmxmYeXdLBnShPD3qY/8YnL9FPRSoMg0iiHUkJhQt6F
58CqTFMjT2gdZyjbZsmUN2IbeFM4o66Bp4HMWmdGnuI3TK8holQHntMTbKwjIPcs
rrjsu2g+k9UWi5f+18XZg0XrLuB6rL3Jzso5jh98wfCC/2CvaGfS4W4U7fIOsp+K
UyNpWxIkdE7b1TBlcHzQH+HmQimhyrR3z75LthNsIRoBN+FbmlWS3tro8qAX+u9b
d5pzL9qkuPeT+qUYs6Edi/SWdKYlqFCpy0Ikc0tYJp+aRBi8H7YMooIShixzXj5g
F+BqP9KqYJ2Q1bDOxQqAXQEUPMHBaWFuDhREsJb89l2ie13uXHKEJA7d4EEgIIDm
8EfGLqTo3rBD0Rjkju/kZO9XAezjITsXaCKPYyXFdJrE/w8NIEtprL70LNM4Rg3W
qETReoYVeWgvRYe/G7X8px0Vc7m3WGfyJkwUJqLfGRLmnZFm+bhYUQZtFe7MQeVJ
NOhWkVu+jxdy5djUt3QXl/WPfbdIEsmHYCOXBMAhWJjpTP1Z2/JXK7XzyIc12xZv
+vwa4b1cdXMzucHhp35rJpE9GgPEnPMPOJ4b+joHWzfxovc4qwuzhbzX3K333dhx
Ipw/qYfRMFcWY4fS7/+ozZ7ssmMiSVD83jReJPEs5TQLkXXOS2UikOci8DHA8E+b
7zJoKnohnsqDQC3xP6CLOdDe2h56Ii9LtLgbwiG0HySIzUmGX2TdEO20LgoVvGeC
lR5SABWU7GqrHOpH1haxdVULyPZhDsdmOxD9qGEJ+ZQox451GnpHtncdVvC8xdfh
68QlQ+hx8xtDuNf3IVoUsHbJ5DqJkHSWyICtG8BKwKzOm1ZLPIWbtlVwzSBp8yon
nSeMh4cneuoyPXUJT+xuhIJH+61MoV/CSJNLMQGTmbR4ThNASBXyb4c58Axb+fPI
vj56iUZvQG8hzpmlQDqdPbe6QHfBoXLb6JmFlyLJsVDmL6+Za+6ULTQYGZI0tGaV
yQMgBQ35IWFkqtxLuT8W2EpyfIl5uO9dLFDXtkDWRkBDszl6K2OoVnBINnrELfag
I+9FDL9eZnYxufB9WRkr1oQyiFW4H+rd7iYuAKy5UBZwXPUeXA54EcbxT/qvO2aN
V8DV3aU17lZSO7ZjUPwCZUz5vgiPEb92dehTw9NP2aDbaZqBJcTYggTs5oZ7X9Ff
J+XXMRbd9Mr8oSiBh0241+eBq9HN9VGL/Xupi5UlLokInOCCQrLE/1MUOfFuz1vd
ixnsuflxcvPdUQ+4HwGH4OcFCKfw1rmSzGtbSWaY/zRPIuZZAZmDZU5XkFJrMKgs
/BN0USiGhagv8GkEQdOJ9H7EkAklwNdJ/4W8n/Ur/liatR7fPjHQSbLj290SRFBy
8ndYpjKTjV/kOcZ7Hc+lhwnEu0baH0BY+hUeZoRxaEsoH+62RAeS9nyCNoHrI+Ak
m6/+lcyJYK7Xvlpt1cxMPyB76wd90Y9/y93Fnr9OTopS5P2FAcsWI1PMyoheq3ME
rPL4esgsHyHJKCPAAmwUJ1BgEz5CfnB8JFsRF73ofyvvnokt5aaI5whtPV9bD/dM
PErV3/jgTfCFAvyxMfgCCFSHEH2VOMI8M+esyIRt/VxCcHLRSXDURNQ35nrZ750W
+mpCP7+lmy2sShVWOMAdThrGELVzsh5tgDnyusZFnjNtBZNueZcyhf4P8PmGDkVp
5QRL46df6Wy3Fv6h3cxUXk3pSLDaWsMX1Up/gQlffyfanZzjqpFP6ulPT9HyN2i4
BqBhHieLdIPfeJl7navxOEvsMrhoBilbVylx6c19ujkXKfJavrr9bjo7QGuvmHZh
72mSZ9V1V+LMLaOIe+50bFr/+qgE+aSw5+z6+3hrgL4ELXqJpvsI3+D84WMkld42
oV2yFtyvtL6Ub5q/ncl8Yb9XeDQzzDnlLOeTsilu99Q/DecMTRpP6ShUEI+nbiSC
YTi8+MnNAtHxO1SoU7Oh/mU5AFOeiKmb6Nv/xSh0RRKaqgaQlF2o+SVce240uXSh
eA+o4pnW/HTJUuApwy5mCMwOYXiq6W/SqiIFKaek7vSboNOCGSutOFMHkvVQm9hr
n7rEq2zZ0uWfvYmdol16qYaQgbvn/HMUVCHTNoeJfZFRzJF37NM9gAiB9+LDuyl5
PAWbKTpurBCOXgjEe1Kzx1qkn+mGRAaJHdIYjXpPDbYNZHSmuIrcU5AeHc91Z8Nu
MxANSoeplLIOb/q6C3U+VHWoP1fP2Uu5E57+CURW4/y+omPmSUSpFGqj+MIlPm1x
k6VCn5ZygPT2hRUnOstq0c2jjNPAzVoQDNG+y7MA/UOoW6FSLIE25rrLbyv0ppYK
3rk3Xr96rHKYQQDJ1HfFWBLw4DkiJ3J6GIvtOfSfmV5M2NSUMIoZIgueD14ZHWoK
G1v58q+B/5D78H0lN8YYeZVfG0ZFVQbPs+XwJhhNsNy1XFMvAViC++1PM9N/sFrS
FlPdPhJWrvRD+lGn7efFVaamU6+U6CnKmHH4SrfIvkviZ2aclImfiZu2e+Ha/JIJ
BGZipZtHqNMJx7H6pS/MRR+uA8hvqAZuLRQ+p/vRBlgKA+gk8OZuzOGfV+6dw7R7
irK0E0lxCLw1a6w2Yih1ihirfWzhrgxy+0gm/ESAHAlKnvPW0e2nnkD8suZzNEfE
VU3Dm50FRZC+ARyc0ejvxv7PWgGg2uGMWEi2gkfLI2+dG3jkwb6N3A0amQpa2pIL
UHQH7eCHM2hnzcKP2kiBDnLL81P1vQH1Ayafy+pNSvOPkghm8b1bxze3eU0bBiU4
sAZ14+WdMhSvfrILSGWel8STn1oOYe4yNmN0Rc68iLpFQmyx+6zx1FREqnGLcQAQ
xnoTZGyVRfc3g3codWEIWZhcjUHXPAbIryQ/YwHaXRagax98OEgTXyNEO9G35m7d
ZIVNV93hGwqLhoOuHgl+IIptCL+gv0pp4pVJlgxg3UyNOX++Dr1bhG6pV0yP+8aB
RZFASmzMZUNfKBp53hFzA96cypqkSyE7YrFP6R05U4cXxdkUMJ6GVC1mC6CiRQYA
VKv2z6gf2YZ9uXrOgKZTWnR9crv3Xv3wIuQloJ5FgrSDjTjb5/QF4JNI+aJOiQZL
ViPgFTMoDs3IUBYOtzFQVjrOv2mcGf0Qphe1cG8BVBAOeiJcjk65uY6qhP+Tv85r
RK6Kd68O0yuByLOz3/I9QO0CSXyE/ddYbD5WQteq2FHuhYZ6UuI1cnq3TpsG/NME
AHYCXI9qlPat8p3GmlshoKWZbzMIkzP6riXce3nKLPQ1deUMH55BcdMce9S+0YKB
wnCE51GUq4RyHbZMKnFnAyrEQ4BnvrFbaawAEAfphFVOtQC8ObV/EEgiCZIB2WbC
mmZsjzCmgVfPTE6FvFYetHT9FT8lPYol5UaMlvgOLLE/E7kUCQG7mKZqX+1zMnJO
0fcmPtI/7SdNCEPP7tehQM0GSq19/4tAHF0SvF9JY0CoT7KTMDRC4OSL859/EVYy
AcBKweL7KBSDgnJnv5KRwt+Erd5rAKFK2f2jBIGuXUuvhZO92Dk2+AKkchgU8X7i
ru2iDsY9Qy5VOGfj6G8AghA8bggwSc81kcI4SOjlW+K5/jff1fWuXcLkVWEKb6fw
L8y3qTXMgcLgmL+1jePF/FdPauNcFZtyZGJVZpHphUg3MMke1GRevIyZOLDYmAfd
XcemqmtpNXJ1Zqs/RUadlTB+WBCc5FKPCbQUUqC2FSkUERnnxyzloiwqC7tUsMHh
v7IvJVVtozdUTl+ClFWM6j0AKLFML1ioeXymFB2jFCwaxWOhwpw/eS+Z7GE/OpAD
pKHBSIsrOV2ovrF7NvQ9RpHPaaX9E1EAm+a7zbLSnC3iaOBb3d7NhNm0Y7j98tXd
3qqsY693ruYlYk8syj0x475/MnPdN+xGsF/yjQ1BvMHm5XRB6JTelTLjYRRUgYyn
mm/lj/12atYUI5kjpDaEb2c5dgXGepSl0VmDyjRfGAbb0+ZMaoMXadu2NZ8SRpEz
RH3nTSrEbx3QgwSOVRPJg2IEXudOCb70ra+3dT+s/bxq2BNfaodfQpaIfHdQG6zP
SmMbYZVwtSksXa9z1JYPRqudyVgimvMycSQFfD8QQrdJSzOugMuSklkT5dpgt+A+
GK+1FB/rzzRPQSvTZUw1CeZgT22tFue5syE0J856i2Y6m09fuWGg4Pqa8QxUHfZm
4E//6LW9ZDjVRXC8IihZ80QnE1/Ixq9kYEg6+YrzR0PWUBwBmxQW0UtRmJjRKnSG
wQBPJXZnW9RDFt1EfBFT4zwIBZPZGotvsvYFaGsOWOPO5Nu6yhPGYPyx9+sXL1xT
rXElKUcDRZYLTXqN+S0yHGafrgnDnFtkdgR8VrqTKvQhF4gts9qXyDjuSs7vhy+r
cPZIkaV6S+eZXHgpYouQ5mey317LsHhSnOPG0FPkXfifMvGjxBaNXFiOoO0xjIFj
v41g5Hu/7COGUn5dPCqDUoZwSZdIfwwv7EeFygiHhuKjlB5Q2m5VDb9RtmX1U2iE
FZ7Mufip5p63+DtMXXbNSsJufmU0jHilM4t+kB0NeKOlG8EYnswjWNd6fcukx2K0
Vm2xni1MopRJODdALV0iUnUb+SVAwm0zj6wOPUP1o+n616jNXqh2MFcMl5erzlqv
0pHl5RAtFz/AzCG8evYqBTMAPNgenca9De8XV9wpr+qHSB1dlDRRYDfJ+DLFjmPA
7qkUQaejbUikPGVRMmjPPJ3DhH2Ks5nTQINsZ09mUixT+0qwe7FlJVLlOr/X5Vol
N/rJV/LMxunb2ZGMez8RXVVtbPH/1JD0ynnovL8LA4xC1fJoB23uUC/+BBFJoYEu
VmI8HM/QauWVVYuIgJm4d7XRmL17Dv1pgIOmLt79Ekno3lBjPeeK04sYuPCVrqyB
iAHiE9SFN+0tO4cY8ynTd+x3qiY3Bs2UusRUzdh3LzNfNz5+QPL6UScpz3gzGmwA
x0xa14EPR2geQO4UKOHneWhbvYZ+l9Q1U8znsyPpr8BjWiI3oKF9AqJAr3GSspSv
8MUmWH+9u0Y5h+zcDryZc52TVqftXDcegiqBRg1DQ3qyy+dJxlELsPvTv6cRNqXG
BHEcIWhQErO+uNbnYrUbH4ZSiX8blaHsVk+kBRFLvvTVXMZ4hO8Z5RyI34yxh4XU
a2zbCILPnRd0yGmvb9YOwT1B3ysZrIHSxiqAu7uCTnSWctxE2i+XG2jwansAIdKM
CT3+BZmE4u3DOfs/kxyRYkbib2ad9kIsGToWSu8lXc6kZ9wTISVm7pHT6fl5XTw6
oBwduDqzAK8ygCUuNa2w+udscXy+zkAOZ62tBQokb3HSaUUVzIYxFdI9EVxf+z8s
w8c02+0rpV9SfpRG0/hntkvN/2GX2aTxtp0iwukCGLiZuwju53UqfS2I4QzJYjMn
USmehufmPmvnKF1dWq0uoGv69AcsuM/3CuBF9wq/9plIUgwp7eDFNr6JAWr58xYT
ONxUa+s285oT+JzTf3J5blcGeGDKfqWDJ5WH4PIVJAB+Yf9ck2HpSe+/51IKlYbQ
ySfiq/gyc6tTo89TtQlbmPA7YNPtN6+XQHw0/QxzYMqcTuIksS65SBmo1vj6YuGN
JHZ/N4wEF0mO/xmP8GQRUWvBC9CWL64JnTaY3QghDg2g3OoDVMICzOdEXCT1HNQ3
3k/Fx7wiRfT6vkxUUpyZPOkJ5sVBNSFp5206RPeyTMTMaeD8QSNJaqACiG39WEg3
vBf9uDfPkHzby6yp3sMsgzm+TA0BDpM4dzaU7GtcPJoUtu4GRwS+0185eF4JB3Ec
h5QlD0tp1Hgdhw071Wgbw5XnJzfaygA0q47jS3Tx9UToJl8vBlJK74LgMw5f4UqE
jK6pEZtA7jNXOsu1/EstIXvudo+zborM0c/DbjtOO+m7m/CudUjJ2ATFw2Z+LAHu
4kBhx7syDySR85TXp+w/6CVovNw8GwjWlzeboqdL/x3oSi1YqHj5ttylXH9nbQQv
51zS19cmkDnnXb01W/HFOOgaat4uqCmcHMdOGfiB+8OrpL/90EOwA3gBYRQ4gqxX
SZ3U0muM8hjhKfah1QNqL5cQxQx9ZhXVkFGtpL1oPqbTNn61RA2Ejjr4KOJOLqH0
wULHKP5cw89ch9WWDe87/a3a79UtAuyy+/p0DBLarJF8+Mlx/bjEloWP2Rulk3eu
o6FsK5D8D8Rv9VTktQC3hGFGip4deQFsVrowUMoN8Az0Mp8o7oEWQRKgmzxo8yUY
GTI/fj/lzQ3L+1ZG0b+TKPrjSvU1OWi2oZLeqYj/je8Y03vXnYpksl3YqUS8FvKv
sdiOFBz/PED2Yrkc6iWLdk2CI0mwdMeTVCOqiwT+usy2bMhAndODlbmNCDWNE+dP
ooWcASOpbZkPA79nsET4PyckEbI4hJglkEbgoRIqCjHH9iOrH9eAhY12dbYfy7yt
AWSSXOUgEnV1C+bQsJ8je2buhM4cLf1Rh6eGk1aL4MClSKM4JwlirxSatU6dCM10
2+dpo6UA64/2d0WO0Pnzj/aEIRTUrHyn5zzZpRPIRh+G/Fe4HsjndCRIgNkq/9si
IajJdbbpqHaWTw31AftPqFTI2fhpxeof3txuKIrr3ag+gKx5v3Fht/uBnqkdJm+7
tbhgVAkrsQRVS69tulNvoJJYQQ0K01ZTY8m4l5A/UYL9FswPlgopSEmQGS9bJ5LO
fixYAn1FnfPSc8JTCTM4+qBNQk9qyClGYPN2kWlzT+Us8OBsjCnUJEYzCblJKVvW
4MomtOOc8SmBf2rFr/gD/HHYRBjNg7z2TxocbI9oGTPQbUldyKzXIz47jH/rPe/F
ndfcdUxVm1gd5wj+xQ1WJZMDtU3wGM+QQHQOCMiKTOnoXMJlBwFR1Ynw3VdC8hE5
HkT+kEWi21Yr1NeUhs4nwIcnEIPHOiBeq6RJBu4KDIh4c75yCesZgs0B6dnAICT8
ERFe7QKG4KOrwdJYkAbC9AMjcERkidQCQ//vshBSn7liaFLVrEuA0o9qr4jvAQQR
wxcg2/u0A99M0g9DZoKGa18L/qwoaFFBz8UcIxiEgrPwuTV28wgl6D1388aforNE
y0En3uvvo2ZJ4gSQhEqthOSnMqI/G4KvIW7vow4bD/OVMZnZSeu69IB8yZJzu6Ge
av1NCliwFgh7qLwklcCfX60c2NpjT/HwCNmH9Uv2g96NhL3NAUpsNIWMXVU23six
O3vhs2PkVDeY2HKGFWtCArWp1BVoy7I8zzzo3b4SBgJjV6Lq9rSCeDzQ2VyQI0sr
Bo+pNGZQrQddqKtQIa9u1vxj6KIpl8ABCFLx3LvyBUJXai83sEHfex4p3s9ePFbJ
EQOTWoQEjzqmFFfjcHz9pSHw8c7x8kUFG1LsGvrZw6KrOjh68/uR3w9mVJMaDXur
opzACvWePgjjFbzPeOxWnD/YxAvtOv++tQxr7kFFIDzDGCIkAX9eniKIy0jWTQCt
9LAgZo0O3pHVo7hzublla8y4CYKZrdTa5sR12NwzvzokPX92rB0Hzg2EemX3olXt
znlT07L6SnV5XUgx5qfBPVlKev5BvFdKoEsQ/9dI36DDpX2Cwq+QWcfVfAFL0HIm
N0PqHDsYKqvHAn1IHS1pKezZqeGUy2Rf9X5Mp+1hZib3TaFpsp+8kNjeH/ZmEk89
JC6+69njt2C7eDC0MaItjcNjrGoq2aA0ZzYSRUuxyezRpezKVm6E8VrhCszmWjqw
RfCZkORid8vqXT9cS987HKtqadCLNOTiWjiPWtycQZGAw2KHM6XerCKDrBY6LVQ9
pHLFfd5TlAxWo11gaHtJ4DeULT7Rpshj75hKhWJZBFf4sbj+vqrnCvJmktCE+uYY
RwPIWg8FgNivgIt5ycQovH3IBuV3PoVMZssZby6qhaAF+rJ2+6iyb/KgRy34E8cF
InU0/2Ki6fnyvLtBtjhC64wme2Q0Aag6m+R2jRamm6styA5Cq5EGoyGPLfOMIuyP
nElheP4hxjyT1YweV+eA+zu/2CFqrx/qAzpsbCa0mx0pOIjzcYtr9tPP30u0ARma
qQEzKt8d/ApDKHhVbqRu2Zl3s7qW2b1qXSnwC8kALeK0jOMMtMfaZ3+fB343L6fG
Pl8YdOir+vx+9dt5asPtxHkZpjLZ/uYctTVJmGYhKsYzU6AHorPOB9RXjL9WM/NB
0/PeibUVmQbZ/fBaIyHDve7vBRDAto2Z2MH1SUx2vS7eAttKSPKU7qfHwIPWNz4N
PQ6OFllBEcfmfvOwXTT6afZjT9XyXFPYB3wgaAss3uErGoecP90eikcE7uX6xUmI
35jmlnsATH5A3TTu6uhKkkKpkJ+CbDjndDayvL1Cs3juIiDexH/0xp4BcKzfj+Fs
mciRphUOYXOZwHNZ8I/29lCVZOyx0ReuUw/SCiNa2ETvjezsGPb3xS3zCzJzQ2m0
q640wGVvM51zaLHukC6YXnENJdt5NtIKs75Svm0NOz2F6MAD6rvvEQovWXXSa1BC
TlCScCRpNN6dEDMCWQi/ILMCgG5XkSET0A9c8Ztj2OOZ6WnnOPYtIz0MdSBFvelm
ARpexS3ACrfARK4LU/DdPOm5HJkc+kmn6oGmWlMNFSVZsDDislm9u/aGtZ2HyAfb
DIOWwq1IXmHUdzrtQV5VZYC1Le0ZQH3DKmdG1c+lfRo9D5TTAJ/E5sqmdu7gBB2B
QDtjgCPS4TpTuFRdLZO3dPB9oruATsRhRCmjIz/7p1QHLDwu7AxkkYn4ayaXz3k6
2V57P74Cc1htalsGefo2Jg8CDmwYxaQxdPzfxuVQqMn7avBQtvqihMnvJTXWRXC8
Yiyb9KH7Wl6qoQfeIn97Wzw8pq5g3BDwKeWZlF7/nVJWi+Oldrl64X2KAzyP8Bhp
AXFGlSovH8DvjlzZO757LlsTnRF5lx8vlL2kI8Ka5LMv53BVe4Sixt9cwPEcHIm8
IFBrDV1hh/T/JCoHjqgbmVOEImHJmKY2Re1E1t6kun/m/HTNqkkEvdVWX3XD+rln
VbJ6N7gbiNdEA2M26VuCzWpurWywJVYiP8V6VJQqqnzZHxmSvDfKc+Mqc8hCvHlA
i18hIiOqXAHvntfZmLGpZZs3z8a8lfCh0UtS+XyqTxB6HnxG2auhhGAseswc+snn
inV5jkj8csUGV0LVXMmSZVKOSgTzF/kEktBw6wQYUq9K1/pQVXiTKU8LSIWvoVIN
gZnhIVqsins5I5ID6Hsh9PIbA3Tg92qjgOJy0TcJ22lJy4Ur1oqdsCak0HXwG724
U004rS8yA++GnD5+O9Tbw/daT+SwM8PUMoqM5aHHGAg2/tDWr3mnn7iFMJ8Hr19/
Eg6ujXG8IlZ9lmTeS3C/TC9pif5Jv0f7ZOrBA74Q7kkjHlYrW/FqEnYg/2PjV+od
bZNiPUR0Ks2LlgpOq44f8psghw0g9PdjvanBAOmqh0ESpYQDey8sckIRR69bFJpO
x3klpTmseNwQo0lEXQM5RqEsP6MA37Dp0oPUOxpqxKSmWajGHzdF56poSK/g9Gfn
KHxwwMkJjJizqE9lsN+m0QP0Q7ZZ/22Pvw/dmFV9mJGv36b0SQCng6qanJqPl/XC
2+5KieO0tundzD17Fb/KIC/yENSBYDxeuwawZ86eozmPBXN+MZnKBmpBetkIghpO
Nc/wgbLB3AHsWdi4MSY/ZkmVZfjjNoOuy3inRQ78SrBbT7nYjYoEqBkoKgLyihuN
HtWmNDvnlgLW9x0nJ8Jv5bkupB6lJUFQ7wwA6SFv7H/rH7c0ipmBqBrH0LQdm3NC
sEY8TdVJynbSM00A83X2fESjhMasO3pXNlh5Qf73eNj8cvFDCH85eBsAvGy09R7i
1qmL+rrFgPGWTr1xO9etGKyP4VBxvkeeAGkqpPfKO1QS1y3l3ZR96zvNtAR3PEK4
3Bqo1flMMUg7eP0q7YMWBcbGEyx5C3aVGqEuC+2FiLhWlpgPkhQaf+58G/ymEdK2
hGbPVuMi5wWLmd0XH6bffBlaU0n7cpQWY06Hc8SQdsDlFsPAyyU/hTICK/NNoWUx
I5valF4PLcdv8/qAr0XYL3sHCxBcOCAHwBJaf140/ssJYp1ZUM2twXBrmJaq+X9C
pM5SJHpP/440wR7sQKP6ibJ9829oxBGdwT8Y1abFPfPifdm1Lg2/1WCEx4vIJly4
9cBPYvYdyuD3eItnzoKUfOoZbZD+80RpSal5AVlUas0nQHjdCW2A3mv/KB0Wbvf+
f3Zgn/674EzRWZo9aqlidwc27cWLFrcLl+ntN6Zv5R3tQjQokb1QbmyzIsZ94rOn
mNXYscEosZDNi/nKH+a1m5bUNJlf3n6+XEbskVPeatPW3/8t/Mre9h1BbG8YafU6
79qfosks2UaKQy76xz5wqJrsDyfE72rx5eVOxsxcrmEjeALF2dMZiIaW4phbb5Y5
tSjqX863R1kqmSGJSAXJ7bFSGGor+zmRWvxr93qMZhDkpwyHkX606rPAp1p9WUHQ
2yTF2iUDgFXzqBROIYPdHwpr8/IjK0DRrsJMQaH6sZV5pbhQdhl7l8ePSlNk6Kye
n3mHAhCBE8EMpTw9k+/4w8tKzNpeUqmEMiDQaPCvIWD/ZXv0ZCNzcT7Abem+LNRD
w33C2WYr051mV/AoUF1cKmH2A+8mnHDq9tw3T1/Mt3qrBtVvAivJG5KFRIHHueCz
L5mOnUpYI17H8C3oSS7W5qw+tfaNL168pJMdghV7AnNYrvgZmVPoP51wiN/+NS2e
Z2WYtiZ2FKOX4J5YjRJV1J/pxn+1B7VLqoTKGOGyNKjwKHf9S/aW7FM2MYeXDpA3
jU8psK/+Pls/UWkYHbeu05caZrFn5nPCMRFIYmfQpfjmNTXOzuEEh4mUkWNfxNAd
9mjqnUQD/B2jpSHS/ICbZbT+/LjO8HAg8oHA0PXGdbnSPNOy3r4N4P04DmaKkIp3
VVQsyOj7Zj20Jz83GA1fslow4pOEiBy1jQzOXRDZKqUNg23Svq3oXyaUoK8EaWFl
Xj/E4jg4nN9FKdLGTy0fqF7QNb1hi9CRJ24p8CLlvekJ/ahqIS33G2MbQRb4MxOF
ln/yaaxb0EghpCwNfBlZlHI6h4uZ0o7+XtaCbtuJjJ7fMuR958kmx8jDx32Xnltj
bLxl/TOOvpUqtRSsWyARqSPe+zTj8F50zk3ivgYAicb+PwS5jUgDfPNw7EkKMmBb
msRScaHfxhAaseINaJNudcQCRQD0ZFqH3UhQmmTbGOPdkZHGyoUbwxcLZule0kJu
cq6OuxqAANp9WU8Y8h4Phma4Zlf5cMZ0OXH1o/l/NCVYu6ZHxR6prfAkNrdZiu9r
zrw2LPW9TZ33X1bPhpWY7PuKWNQ+tyfwmbMTUWnAgG0Zz15fgHUwM9gpZDiklWyP
3UNhN7DUqshv4c+YhjvoBILFF0306TSfHG9PlscgyCg+l5+cPPxXwIe3oTpZo81T
Ufsyk9H0n96Rxjkl4+cHysxLAJoZwKpuXsQ3r1RkDXXY/rSyT1GzAzgTcqD6CPVq
lXEeNEPesaUpEQ+6fMbALlRhGCkIDbgRML4BIMu6Hl3CuBnekp/bevLiO0hBf6Js
VXPl+6h/iJg4uZK/Tv/mYApSFqAB/Q45TTfeToDYPCsBV/+M9h+Dv/8spsGNHlgA
LBOkkWtOPfaWTYLYPfKcfoLsivz2qzOp0l2RuYUxGMqhXh4kds0wPfnrKAyKzLak
CLfx2SruCmcCEVsfD55A9oTNoA8aBCdmVBZviofk6GBJoYitN/21bCwVuLH+bms9
mvpffFxhxgzsRttARHHTbyLrpQXvy2BAu7cXnr7LEEsPwglfCNAhWxPQe6YhgIJH
Bqj2q2O5D6JDICjI2JYn7/s7fG+LU3P5VFcQaIEvdJewYO8xCVB/EC9VjaUoK+rC
j93QD2bar+6sCgrprzFV/EQ0Q5CrP+9bA67ytwAbA2eLAC8IatrV67JaSWetiRYx
IX8O3duU8Xf8TR3LCzKs8Czf6r5lSAV9VnbrqejSVtnfogm1PuzN47poTMvqB3De
2QaMRV7BjlvOXbE8RkunPBdJPyg6LMou+9C0F/Lq/FS6N/38NjrZgOC+A7NmR2F7
yI/qL3pkjqoRvsFuTSKGlh86CeMC/r7PFvlieV73xIYoB0Ji6efvaW11ZqcOQgo5
6dP7pf4SqrEPJJoqwWLl8q+6XStIcYasLx3lAZGKIq9f8Sy+ud2z0ZlIJ6sKSMY2
xhdjsoeY/909DNcdDdJffgqZu5rM7tIVEMHWBll1Opj2k120TMuYiiab9G/JLBXZ
7GIQUfNRewKrFV9HyWJtIbs/9dy1WuHbr0CRq9NvzGrhoMez/yNcVnqvBDt3DQVO
BJNSFYdsMMPv8JeAaY+JgSH2gaL9DMeHeLs+mcgoH/iQgvkXeLcdr84Cf1igfnS2
aa9pv7I3nmYR3F/qDWyzKBCN2mgoJ3ouCavjLFhUicyMQ1KdnYe8gIloSde4izTd
b4YHsnzX+gIERCUQlykz/3w1Fdn1bH1m3gPbMss3VfONWN3hsTTt5htTXWBA6stK
u/vJemkk2pCoJ6OSnMJbpN6fgGw/+b1KvqHHy/BcNP6zySN/ecquI2aZJrDEyVle
sS/BjNO8aYTR4HI94ylvFtil5qmgXT+R0NUVpyl5miR4BOo7bdTc6j9UsvBeYzUS
VBuWWB+KZLVoaeevvAT6+++S00U6Wks9GHfQPcIPmUduveO3x75JhBTg/f0WLC+p
Flk4w8b/0KcEpPU+fZsZS5ISA+it7iSApylIJwaWY72fQGz7JeGwiNse3/dHbnr3
mLVGhB0Fqm/dTAxqy9I8RYdIDdGb1Ds0vAqZwvyB5TCjODkP3YOsUXprs9/HDJmr
tmLXQXO1nuYh0m+DraCgCONl657jMnbVeTzH2LrkO/bf5+EDQIzwwjXOUm5UG6ec
uFz5JGs1bpIMxfjh4/Sbf3fNc3Kfe2XD2SuDp4AOu5Ohq86cR3HV8bLvPYVCo7U8
FsluNrihwmMXOEfk9hpM/iteDQpOalL1Z42PdCmXuPwJG/Utnle+t2ev1uVDeTZR
Y+0bJLmsrprV5XPLQg2GvwlYuR+et3d5SvD49KtWx81l9ab9GB1/beYcTuKYx8hn
dF+1rtZPyfLc4dRfeV7TbrZM1DZp5DAXz3e+CQxE7CodqhJ0GWXu9w+dzL93ZLEJ
NHdKmQQX2y0MsrGWV2Fy20CJmZCKyx5oldvHnRHvDaU/HkKTteXQS6HttYmctlK3
bH7l1LgZ3GgPSXj1zXyRytaHSsY+nqTRGcwppNNQxFzRy2pBB+5S3EQU5klpCZ5l
N/iqCEBZKvC0cMlNM/+SYEL0dkA2Nqsg/DpR4LtVC9rWEdoPu6g3iuhT6r3ZYVWz
VoPIMqfRzYhoRSAv/w+vM5dJSvJaxHDG4IZ6ZGyZ8X/3ksfIsmTZlxriA4Okn2Mj
YCyjYBy6FxWwJiTmT3q53UlOE9WlMUpyuKVE3e+hw+S/i5YGx8foumzpYb4wA50J
unCC0bx/ipMmq69KlYDBWZUQdqI/PxLvxndCzCoGj6HD6YdK7oTwesCPUqjfSCDn
gVG5eR2BuWLe7mZXqMiLxOm5ccMyrlZdlYU51Rn2dvrP3hcRfx8oOEVf72PcsAqj
WAUBnq5LQ8cFadCQtxMFYfCzJdjrepuPwMcYVQnjxrl84FhRwwFndeK7xqdQpdVX
uPklwIZL891PewPO0IIgptgRZHc0qGl/VghBmLPSg4fcUSbi+s+9akkoFNoQwl5S
tVGudnS94sGUEIUvcCnD7xg8b4CykMs0Hqkm7xinYyPn0yQ/6ELSgnEFV31hZRRU
P1Lo48gmF1e+zQm0CNeMcdN+JF9XWaQyrjn+TBiKqJBSdYayZXnQxqf+vvkv/jww
ZmOS0dcdLB+Wij5dSe6FwVJO+67miZ3IZIXabFbMaOhTuxolpuXQ1RauovqzgFG8
M1OxKno1Dg+FJmVLjIYLYsoDyX3gZppnGrzJbOtDYuolfZAReG54PUBOFPHGG6LS
pbLflCnS7l1GgIlvLi3dMGGOeK3m/dh+MbFH+fRATdtFGf9UW9Ishsele5FgIFIL
svFyXbi0PJIGSeLUFtAbul/cKumDGEGLm7Va1EIETALbiqYFMjNgWddx1w8AFcNd
H8aGC2JNe0sn3a4s+RQj11IQm249oJdoG4wr+dlDQmT3T6JKhKwkXEt44uXON9g3
U1YEvy6dqHfD6svu+8Ei1Yv00GuBC/ZY+9vH0gcgISD4UmJDVdkkwKlqOVo6/9lb
yrBDBx0qJeBppzr74YwuZou01o6hqBYX5NvAjuunBAN0kNkSqgIi1WfIMxiT5SCJ
Qsmom+MBMVz1TqPv06odItrfftimD6d7kDjNqL5dQnzbLGkM0dB0hefmuyhEVYbu
rI2FvERADdYEioQF0FU5XsKP212Pur5NrU9yxJJMJNdPSpQr0E92Xgwsxey/cLVW
AVBHmJFBEPpR/DpGVhKAeT2ttXYhx7QFXoflUI4OgoctonPvf8CLoG0xxUzXsnaM
bs08eHMZfKQoWFbq8d69H0cseljpyYaJPjAJu+hZz9/cx3IfXixaInLmTap1o1+Y
SZeYxQU4g8MiNyN5P4r5w6OFmZpytoUsOUjxERxHJGArFpcGfDH7L1+ihp5rAsQs
aq3yDNIlfn+P67SCA8xnQ1tSX7e0gckraG7JzWACIKvySnFpJDr34lYQZyEhgmZA
nDXV5rssPa20Xng4aVMVUF5wFmN3rn0U9lga8QNNMnqYq9oCGy0I1NYHbGnSRTe9
FkEqW5Qza/IRQyzaYotEA8A/K8JWSG5RjB6TiY1sEGpDEGprrd+xFjTQhoEDqbcv
bcytJDgcW7fx2+ur49CxGs+QTyK4/1jT64I3RwHttPkGGivfjwW8EJ2ReYOny/w5
u3541sOouHsK2eDH0GIHMrBrzKGMzFQk/3jo52hajXQwj+1d/ycvqvzFskp2hOkZ
KGWN0xW2DM0K/HScfFQVjvdmCJ5TdyTw1sXW2Z5KVEEVXttmNaVw4BltXeA1a7G/
V+egD6n0lCxNx2uQKYHe/Ehn6mhXAaYl3XSA8Cjzk0NxBoS1mfKjdg8JveynVDuy
591X3m1mSWxn6tWAuSPf97PXSVoYSY4q03ueBC1Gof51p0xY0XjB8L556TFDnObf
Fix5IngKDQCqQqwlQj4c6yCEgkFfN/Vq/BfmKxjKrZVEi1b/pQrERNhEURDQXFWs
fzwWalHD8+vWGk1KtOSwwHPfRQ1KRdNC5B93Ojxnxp262PbC2zY+NbHqEs6NOJ1C
TOV8duGgPnOAi8JUe2ZWbno6SKoxgrlF5YBV/4nTgq7wENKAAVihJjYTQNt0rO6L
2YSp2OcV19OcZ5uqUI3a3m/nLgegu45JPQFxkkr7bCt2h5Hg/8cU9JWmV2od+zC3
rF+CGM7GKPcv/CdXIZB1WYvepTS0bOJgiITOIxoqbtEvY02AeBJDRSZzNDVdOfut
ddoHcBPut3AfjB1gGkAmQoWnhVurXNYgo1/y5PCskjs1PuTCfZsSpNYyzV6iyOuF
2Rm0TSpRD2aR0s7taSP4xRw/wyxmRBTtpYLUefVJrMx/5luR03berB00dYMr9Vv8
5bkg+oHTyG6o7U9GUfu8dwbnvuK51qRatAhxJo1BKrVZX0SfUzMWFcFMbmh/ZZe3
Bxe3cxcQz5b2tJERq7988SikVafTqa3NBlgRCuwHfZ/gSo/5brkszj2HwoKq1qtX
DkX88YIfLRIklx4O7mtvbNNldmySI/JzHwJvKDlqq3HSCMn2G2hraC/S6UImj3n4
XxnT0ei+50b3kSw3if84ot1rG9S2gyoVSnFQtNdywDV7i9gpekKUX77NwHdW0QUA
spxH+nco6zXErUSGoEQeGztlxaFnr18kSFl5RmiUTu78UzHKHLssi0nkeL4hznRI
3HBP2br4cjkUXzSZPFRYQln0ga10Gch2G0VxkAvLxUfguPHHRpcAnWXmE/PYoCNj
3nXcQOYYft6Ls+LMv4SJzEQ8nupz/yJnqIQjeM6SU6VTL4eIwojXYfAua4ERpFD8
yvff+FxfxDgWwA2BkmJS811ENIZlXoq55e6vhPP35IHEg930LfeyugFznOfu+HQ5
hOpcLMoLnv/lXGCmy2WFL2QUoUCfIfboUhbMlqoi6ohDoxFfzBUgi0R0GcV41311
s4sIjoWQLcSVeC3j6B6GPrvcTuTvqJRNyH+tlSJ76Hhg/Pppgxb/O54pbvF6m3KN
LxAHOkvJ8dnhjDW48QTsdu5yJhcG93SiwaATfUpCSKTMz9kSOeXDmQ1tOH7c7+5f
ZOW9mFb7Xjfkry+mu3yOa9gqLTehuZvjBpgro5qb1CZGrLJVGellaIjRpGPY+QtH
gAUomcmX8O0L7vYiFBxqILmji8v8byFaWYxDAdHD5vahEZd75Jr8atcSKZJGmvne
CVZlYjbAVh/NLZJc62SHHY6+/JCVSVCnztX40HFIBKq/JtFSVesWApmvlFqz1mth
0dDYM8/6w5P56dU3bNlCW2z1hV7N6acfBsTPvrBkQ0QPvpy2ShvwbG2VqB7Xddzz
rPY1dCwSmC8gqNCHcaNuIYyKoFc5kxBheC3GelVKLgFcMRExp9s5pnKEAd9ipGMs
nY5hqiksxlYOcJ//Bt3HgMSnn4tw9dhYNeMi4M5wEEZ2mxtl7dzO9WBHU2F/OH/C
3otW3Q8N+j1N+20A3WljJ8GRSHy2YeBdlF7CkqjF4jxFYPNdqeDGih8MReeN0CXJ
hUverzJkANckJyEdJgBw4qwx0XFwu5ehjSIVxco2ZtT2/Cwg73OU7m7emARCLiMC
mbyVHGIwWGFn7NjnhfYOeh2xHI7l80Yrit70y8IEl19NHJR7dtJpFVGFM7ci4YX/
rc30LtM5k5rTW+Cl0JEyaGx+QqRP+GZvpLst/O4y/NcinePm7aLlUPyiDUnXW19j
esUZay93vDu57yBzNFEkmhS3f3LUCcUhJ8+2Cn1/wR+v8bwOucc7vlkhNPaKTAxA
tHrYoCTh+ZuXVO9vNyALku8oBaZY+O8Ip7LLZszUqlJxM5Ff9rvpBK/tipbhnCB+
BD9KugJFlAsS7zfF1YCu2GYWuPTaJz480EKvTZM208A6biviycJYnuvTL1TARRHm
BuxI0MWM0xSeApWW62+xGDnsetQQ0yQjzHKitpUpZvPj+iFa+HcxY+gK/vCu2iIh
RZQlXsc73o0sU6SiVqSz+5Lsnbf7pvVEPHFZhdxbRWXvh1fkleR0pHXf4Wc12FG0
JBOTEZoS0wJDscW84dojm2p64Iet0mf+4iK7/shQuNieSeswtZhv7pwIbF2awTa9
hwDi7F2513/Z0bCW7/6OJR7f/JLkLhUY3ztUYzOPHuPvUfomceMUUAewjgXFd7kr
QNZHFByINkntSNcflu06r5IGW57Xs315EMLAGtZMp2eVwUL0JWp2f9hFdtji0Rls
t8xWm6WHWDzzcjO8cxcoYcH3A4sGlQc1fow81B1qy6x2fac7V69ZbOiGv0tTMeRa
EPl9tDSHOgTr+JyoCSlz9+CQtY5JLkHWAkfXDVkKgLbHjsatOn2gWdzqGw3ttpB2
ffovG8kkDcSJ2j3F3YnyED+/ZoOXor3umtLajpNB5YQLN0LuMUWODxoUKUkvvT0L
FH6emutv0eZZe0Qu0blQUY6+h/LMUe+/3MeI/SQg4A3AK3FL79wn/7RFNLAFeD34
Fy/5CWwjMtlldMddQvO4gdqIam/4NURnYCI4uRLuBKYm/so871EyMzBMg45R2jRB
pvgBtszWz7gHWG8I7UPFAnndVQfwJvZFJWYTBdOj4Apl0s4/sUIwVtItKr4vD+Sj
2hRni1AL0qC0g7wl+XbNL8RINsLadS21RiSrcYb7riAuKJe7SxsVlyf387Qxj3f9
+CrCP7yGy5BIj5pngq1KS3VRCCTSN88rsqw8Tss9pthOgDnx6CQiNjQArgBm4T60
4dD6QdN8V7KDiqe8RT1QzEEcMXEoeVlhgI0mKJ7sJC1Bn/+hfchQgAd1/GFZGUit
w8VIfLlOguwXJ1YGAJlJWRAx38kx4KssQXZuVN8kO2BdYKT39yOJ50PCDNYQm8Yl
AKls9xlOJzZzcM6GGq12jda0etVCtzRF8+7cV4PCs9H+qhm/2DYuiSU3oyXFV5XM
cMZO8aVTf/OVV8a3nc4MC9fhxmrhJ7l96+iciCY0t2lm7xDEyBHJwgQ3R1KV3G1C
mIwi7z4xj3ulDyShTOj0VOTIqnFQ6eCskiTv/RCkfaOfO7vUiYOj0AcPPrtMVNPc
EHY095bBCJ3pUAnXanDW11sPm28m08bwHEbY+vHxlHi4S+A5J/Hfz63/RfIAlSAW
wKlwFvk0pdbzdsR3+9p46fbtHv3PDA30WTcge7d18yWbHuw6kAG9wWJUc9GQ8RwE
Mg3kHMR8sR52dtnAg6OoD+ixmAaD6Itlp3IzTNOoY0N/9oR8IzRDjKqqpmrXEs36
l4EkYBw3vndrytQonzOGbUDrrvApz/V1nhNYyU83Zr8HarEz4Mp9QzRA+SwjoDD0
6A61O3iDTMVNZXVyJBVUifjZu01b5s49s4r1Jm2Qush69xOEV0rjfX01PI9o7twe
dluhsfbojEjWx4SaeH/xqQnx29WrvwI/dpWYsK4D+R492UhgRTo9ZSjSdYNz0im9
5lk5Z7t19lokVX2ku2wimoco6uTwn8Xi3DfbHoIVdqv06VRdUgy7aBCccYobBcYq
MUuCljpwCOQAhdDbnyvuWKUCdbY+FjqAC1uv30CWPrKXQ60B/jYW4Kx/d7W/qna9
X78yu1jRM3s4YhFGRvvKVjtaT9VzyS4XR/1aVBJF8S8W/0x51CFMJhBr0FoqyYZ1
Q23S9h8wj3Z+4pqBDrkt3sX3hEozcy7PgPwrwOs2uk9gDhPd8pTUkZFgMLLqCl6x
P1fmmydOEXSwjtSR/R0uT7tjM/kMKefOE5vd5rGkKXai1+XorjNngJ9iDdMdB7+s
1HaQbkOFSZdALa+Y7mmIgx6LcLzLYPJGuDRN3MbLDdYeujLnSyg5lL0W3I3ixTTe
YdEXcVMX6Wh7vOntox/W8wsnx++Zfz6r0i5gj7Fb921H4c4v7pr4KqZ6ZBaTM1Tn
oFCY9HeKl196kDpUh6C85gUspP8VRStUlGz8adPCMlCaObYH2V0co3zgf6Tpz18K
Pej1bAtK0gMN9dXqwd3LFKjz7ZdXl2hb1OhzQM/BkPFQntDcqgPhbkzZ/7sKwx/n
DYelCaVULh1uPbeePR1Qxux0pF+pzln5QMu65IKJpB2rxGqcRjJVbnl374tkLHQd
8i2pt1yFEzawpvUo6+VXC+HXYwJcZi/09WU5kid2ajMA8Ju5ut7jKO74v0yJdtio
FhLlBR7f60LQeda4EiVbo6hxdArhIQ9FTuVQV+RvibbfgVRlyFbWGVNIr6PcnPes
JafuTcGwn92VjbwBR+fQ0mPutq+q5XjcTXNIOkHggw6TWnG3emarLeeOkgDCRRVs
W1LzCky5bN2hFz63xQ2bwfhszOfZM6hsflP+FDxYhPjvkSoKtYEW/gqlZBO0M2k3
c1kN3NszH+hVwgkd6u7oMlcvXfUmHH1tBGK2uxv7K1iC/e2HhcT2nOB2T1iob6kL
DimPWiblJnYSfoy299Sg/1gykdxI3CpwEKlpoy3VSEqgNySZr4AhiMwAKrT1QDZ0
qP0YIQqpN86Tc2UWxF2/znh3FVNy5IGF/MkLFdFk+cnlFgW1FTs7fwf/4OpHnO9H
ZR+uGlGS7QKn/OVyo6jWWID7hKAO66023WueMBsRcWC38/Y7gHJGtBCNcqKNL3Hy
bwa/2JH9NuXbxE9V3BFXLpsMKTLLNKO3Sn9+wu/i6CbqAb16nazHD5PCyCMEkREt
h5ypQExzw6b70dWeLZ4nkZyfd+qSY45KK/vfGl+RaF9UQASbHrHxZTMHBcpLvr0w
898gWOIALCvyJKRKGCFatXXLSaZx8DVT2tvdzVdEb8oIGVwJ/mOTMP1y1fdAb/pL
wUu2s3+bmV3bkLjIaxZB9U2wGUdiRTPs9Dtx+3uaz6PoaV511+wDD768Lq3esk/R
//5+nu7cYPLMF7TBsZtWJHnLbT6b8fE1b8MzzeSe258PxHv0UN3amBUxr2bKiGWB
Z/zO7l9cKeujZEwHrU8SQ+SmEAVX1/K+EN8wQGATQRg/hWh2ju6m9X1HQu+ZU2yU
asyTcDIp6MwT4ceRnKnmpkALFWAInYZxcaE4TV3VV7Lylo/Sw8lf/upgKu1P9rx0
HxP9mAIMg75q2zHe33RnKg5HEPvRgoVWHc69Wk2EQUtZaTv7UuS0khZH08tKUsXd
Z48iFhJmu6b1UbWGwG1d8Gi31APFJdGIXdg6fRULCYRZ3TP6Z59FFdAUPePCnQql
cUZL3Pdp/QZEKd68fkzXoL53RsNDpPDQTCZQauvcGn5nU6T6EMnd6yLPoDMFQyLE
l7FbvgwuWOOC5hJ5htVHESvQz08VnGERoC2t3NwY0mswCCAsOniVaRUnrSwmwU0L
vJ6jd3yhjo5CxKzBXYXTUyvGxZMyyMHve5JRy7aLgMVgv3yZAQW7rR1h21f1+yNW
zchDAQDfnVjkonk+ugAfybt1lSS6CPgN4FUgX2RO76B4cMQzj8uV7J8v8fSqaRbD
Fg+OYRZ6BN9MCl9cFVz7HHPfD1OZn+KOxn8rmqqVAJ1oL5wYghCG6dz/BP83oYUe
SoR1Qwl97kdBEjW0VmGFT4HZsEYij2KxORy4CYuMfEhCvSMY/+cEvdk8In6R3A0d
89utiqxERi19xFJpZ5xaOI2HV8FnlxLeeUsm8S1XrYDlOqs08JLp4oMAjmBrRhGA
bQ08XkdRY+sN1OHdznZRyUDQ97p5L4ga118zF2+TMRq7kb/Mhf6Q2aHKrGgeW9Cz
YPTrUCxCB33nOADOtyyvu8xzSbq8kELjK7FQ/zRyvNEnU5kIS6+FDAqYFWcK82b7
W7Bp+wZP4cOVk5Fesq5Pv6vnrMZSaqnNX4pFbZV92ihLpV6f1dDhwliSwMV+kh0e
wEexN2UpmgFoVGgyCk8xOWicUJVC84Y86lZzjLaky1XZUEJ4KwOrpK9HzqQzk/ks
FniXk0FBGVMgMd0k6xc45jNU5KkzcLMcvIGW9wH/0pONsmZDySIC3ixZHklvSpRA
rDSNyn506rlOlEOFUuDytVFh76O2xGPz5ixRnh/0QdYxjuwgAK45ipiEpRV2F3Cb
/Ow3rYT9WKp7a+8yEsHnEXsUfhXH1PauO55gLcptiEuIKMPLkkxrerrfGak8QotY
FBnW5tVoBx71SOgNqIUTQ2qjGOAup1+oPjTbsX6LrxBAEn7OsV5SIZhhgIr3CmwG
T3hFPaPL9ZCErIeP7N01T3xl9MjZwRS8XnM8FH0C0b/0YpcHltYdpSKqs/QdODwN
SSVMetnPbDl8OM3YxTP93Yuuigsic+BSknmiaKGKSXKKHPH8gCPjNBBej6LI9lEv
+QNUJYeFDuJJ5AaIP91IWsWUl2mynon+hJnO5eSbD8IIHTkUA4CfuDevamAC/rud
t9G4hCRkLtKUWL/WqxPHaHp9gN/ybV3X8w0JBmPeafssVFb99YgZ64FgvTsXOTkV
aITcUy3EKh/d21tAs77BeV/tUBFgJ+tlMHCxycs8Sz2CwxQVJm+pCAQ+RNKO4Cq2
7VnA9VFguqdI5brB2ycwJNeXEFky9DilmXicQ5sG+H1XDm1GERCW0HdQD+yUIpbs
dCYkCJ7u301uRrG2FLYgK5ew5yHkFTeLWwcO1CJKv0n45IlTRKr/ziGm8Xl92YBH
XTVq85K+UxKOKNFC65/d7amtEUwCF3Cn0+ENYDNoYur88DvjwHeUwiUlhiWUZwat
wZFd++Ghwf0H8hOHaNziTkA6dZNHVxrgqu7+OwlIJRmAV/kDmUXTKn2iqnOhU9Ex
dGgUiZkikOtXp8lox0YgZLANUCE1pY64xCA2RyLPftWCZSruH6TljpJ7jKNJxW/C
Ka7HXURmHoWB7GA5FVXRoWD7liLeWpLy1DYJurfwKN5GCwojnQf7+P6TrdJBBmKo
wHuvrrBK2RC1hs0NSStZJI5g2ERm8j7jxyIosYlNsJPH2tNjjWIv8KG8WdO3u1yL
t5MsUwQ12Mo8QzbNdBGs47lxqJFle1hRCTmzK1ydfExdta77rsAN2FAhNemRiTy3
p0lITqtso4D4a/soJeF3jCUDnnuRpN12EZ9lKmuqhlVbvO2B9ZaZWBkWEmw2zjX1
iLOC4NSpkNaLcIBoJlkkyoEyx/ZkArANGV+2bfB9Y8lmERxNUxReath6+r9cvaYe
Vr2BqgO/xI57aWsxuGOksTR83UZ4UZXqQPu5asdCLvsfcX9JREnR9dC2AyRAHnQ5
LjuV+X09k7IV1KWuSy6KawKyLeOhadABvmZfof/Djg9o1V5THrBQLDvbYteNE4c/
QaCO+5NZP8IA0d2sK40G6DZU/e5rEadSgs9qfuVFcKDL+/kIFLiHX7NkRRJmTwLX
Wcleg3tIQbSNnFy8tyqaV6qhqUJWd9ofqkEl9TH9Xnlz99vVbIc2P3hYXBeTPgyD
azvcQNwYr1Cf0mcMj22qidf4BNYQXRKiBAtnkHaiLBbPFJr3UwC7Fwz8uKxyRuLI
dt/oMUrXxGeomLuoLMNEeuE3xOi1e2WR6efvqwOnX2vRBoolUq7F85eTHtg65ina
D0gz5mjDOhw7ju1RL82Wr8aQHQQNluXa0QkXdq6bZDFL7/hH0ZL/ho+XUfRuX8RT
j5rWcoeHoZqd2ijaRz/pv/N+aEAZa/v6LJBz28WHeRlTPgzCdz4z9z4ksqqOkAbE
aMFTtXswCVRjnqJtCYB5zZKFKeTJEjcw4vAE0gd8G6wQApwtM+j3EnJhKq8NGCNF
6y1TJXfQOM+QPLPx3bEjjSfodmbly4detz7xXK5NoO4+HzeBV8ZpSG/Z13JfDFpn
Pb1pZBnObOGOw77HiIkbPh7IXEox1uhhbUwSzfN5PwINIsUHdt36iurQ6zcHCF1A
27ioBgLhJuYt+yEPi5zG5SWGg6lLIOjIM6zbBLbtAOCFDZLCDwJXnGusUEXBx7MR
YPkquQSwhjOjvLL5pdOWo8P+Hdqr1h8H0N3tNk0EcfaQxnwljYS/MsXKBGesZ9de
65IivO5eWK8b3oUg4ca3v5DyqD3KeioitblJ7X4Vrjok/JYlWOLEDFDHKQ7vBlXe
nIPLq4ngzbyPSdrEtoi6yHbDui8uzz1zvrryRXGy9SKYFVLRxiV3peWvAirvPMXP
pfu4R2OfO2JWvj4G5proq5fKgXtUswdjGRJpP0PjJX3Vj9VTTbDOpAj4e+WGBsnC
84ePkCnajVAKECzDsGE163WSgZQu+8776NiQYS+XqSk5sO2/Md58fXYgdgO+p27K
H2H32wzT//qh65RrZHBaBqwPf94vEzGlkG56ZZd6yK/5BBy15wKOgv6ivNJKCOdm
E2mnp/uZ+2HuozTbAw6npVfWfI8s7nuwOg5ahfkIgj9IN46qw+IwJL6+Yn2Jjp0q
5g/J3r1tteyFafpeI1TtvFiylzdvXE0A/Qlj42xL1nW512YZnCYRwg2sv1QNyIl6
8bwrKQv5KbiEAtYvgUnjOo/8ilbZDKJQkNwcICsCNNwL05DH67KyQ1n8/TC2bs20
+n+36c3WIqEnvPPoBaOJG9f61xsNdv6XLmVauFgREv8MJomaKjl2yEQDD/rwKX+g
XkCuhwzNdk/GG583oCyLAHNs+gz32tUU0sx1nm+3yrcDlHixtCWOLkVeQH85Sjbi
u6Io3K+tbJPr1tq7u9b95stWz6IZUOA0MgtdXt2di8ProVnz8BH/WsK5vEf98QxK
j4/oYs77IApFblUkVY58Dzw+B5xEGXZQQ+Ubncp5KnAu2ixaqn0XVg23nRMHWQVc
m59zwM0fneI2TjfJ7rbW1SCEt4Z1mctGCUG1Eqt0lP2dLt3O3w4lXG+n95EjLV1a
7Exo2G7vYPm/9MNcsqHkwhGZuFGWi3CxOpb/8d42Yu7tY5njNbGGOk9R5xzAFd2o
iwpJAbYyD9TNmXdcCWNCI9r/MrlImGePTbojwQ+OoThtIfhi6vhIOeO4eds/VKmk
rWnPPrW8GuTcDLwzNVZiqmtrrMu+dq2EPiU3XX07btrLc8dhptdcERb71vxqANR1
Uy7MXYBhYUx8XguhpQGH+ndiyGGvP5IJrT8gOd81xyHs+UdnwyYM0u1D1b6sX3rn
wjDKtmcnKZJi6LvsxlIWt4U67g99juAD18wTh3wuAAcX+23MjtVRj9y3B1TM4jo5
s/6WfWYHjg+1e+BII3CUoTIAiqSGkfVX56aNcOgq8eDliujMd5CgHYxjX2lUISMT
nXTNsuNgDWJgJL6fs/+yc17k7AwO/ilr/tmIrvEBGoaXbLjtv5ni9LWyczg394fI
ehwN4ZWQMK9gR5rGdCDdSy/fzB1pVJoAy5PvM2wAj32coJPVQk9IHPDOmFgCzcT4
+Sx/AgrE4lvDHOeMhw/uLYMS5XUz9d+C47z5VLxk/rkCBM9LQ/zPr2rOvDCNyR0G
WLebxuH3PhqRS6D95AmmWKpIz0o2wIZXFMmbElYeuY6pMdBgFzfVkUMqZvgaTkF2
mrTqHYd6ZDoctSH2oOnshQiCkgvYwuilKL6jJL6Ga3hVFoIlHWqbTv69x3NeNZyq
Gnep/bjQX6/j3QPu/hHmW4PZMMEyLRh9CkW8w0GrVSKw0A5C9QwDc3dxTyOBs+Ai
eJBmOxPz8eQngxdDIeCTcr99ml2QsRnJGWYn/lq/NXRhUq8Dcvmo+39Wi+/8iJs3
/37dZEn2XmWRbHg4odtVvtqQ+o8NL1+kvNKJu8nBoRTPY96XOxl2X/9gG91eiEV3
onfbWJWu6Iu9RbghzvlsuByCG2J4/qUj8UqmBS1pEw2TNxsYfREeQqXTMontBt5y
U1diaBGqbs+kHgpjnfJ76KnPuZKybjK8gUunklRhpS6kvMYIs7eRiDX2Xbh6jAgN
e9vfovcKOwgQ8ZZjW9mpk7LglVLeZoMZINNci52mAYBoY7jO6cLk4mwpazD6/MdQ
63sOE2TJ7BZghBJoiv9juW0QcOG8XxAQZKiA4lG+P8HYYmWVlmSF3Dni0w/xT3Kd
Qjg3++pBkJKigaxgSsOEAU5jE2wuHk34kHeQQYCf31AFyhVxHsQnL4WJxapBoZS7
9iFd4F3CddgRghI9mmjpdLqHwlakAOEx2aFyjeH+jn/bpCsg82f+GKOb1mIiaZYT
uVn5fR7t/xt85nnhOIqAzwFpkfRaBLwy5+9oMSQ/BMFwDCareoldiSyvZWPcwLPl
sCxFku80GfprsJMUZbdxfqWEsqqPFagqjGHsUH1o3f7qHlIMR+e3ii56+N9LNlY9
k/iZvVcjAY/udRTjYBintV+NfBzlIKwEtisW6DlpvR1/uxyHWWX1aZFKYLbwUjA4
RNoxenxqqrJDCkCMAN1zZdAnty1p4V27AdVxuRIqA+BlP0PxzT2GYmHaCG6N8GPN
hDoaMTVB1JYJExw/Lwoz4njfEBm6uInznsG57yoJHRril9C+XQ29fO6nIp3QBWFF
JwgHsdNiiiuGyh0OZrMc3g76rVqeVD538TKff98ut0IFokD0JUPZVZgGgnMvfxK3
q5qVsrIEQfZZRikjhb4wwZeUHOCdMgPTnSEpJ4TKRW1e6NMx9Ur0knxCDtRvuS5J
ncwRITcJopLC/tURDOmNZ2d/e6YH8jta3PBQE9BgyyLOzXApowwnook8RNuG6spG
c+Znp0EejE+DItJCGHzEblMa2iXliFc5RLGO67ZqqG+UgixEEqc8AoNAa7rgVIzH
qe5QFFAtq1m79D0BrQsNZHYZ1aWGpRxpllnRnG3Fovyeo16UDMop+UiBI+04I4/k
Vx7QIOBegQUvFt5sqXaSZrxRJQpcEqrzYO5lRYFusFx1g9g5vau5Sd0teXAThDH6
v372RXyyOeFXAh7BeCxfOOcvXtn1XmF4wD44QKPPjvG+ci9lultYX9Exz7U3DgSv
dxi8TGKxH9OfkMK9p1tt16tvhP8MDIKHQaq8unIvbQqgXF5IEYwafKgzsL5RRZie
aso4wXAknpWmfo3iivnqYb6dDW/eAFIAO+5uOxpkPEkyM7dqSRcgrF5gO2citqw4
SHbINUwZGy6YZnjzxuLLJCUinCCVdJBDRbomFW14tmn1IiyEh2B8terGALPaSIB/
iOT9cd8rwpDx5mOJ/TT/oeVB+YopFxRYmBZDS9B7G9wCa3BZ1ccEqKJejRUurAjU
jneEx/38cKpxLbirkm3NUluItiBAUfgXj8XuS1mcH9t/0mX+AdfyB8rp6n/Dw29A
pEIPYoaUGN1c4TG4dmRSUw0o/ufuweMGhfWaFCNJ3zLt6n5Tyh1pE05OzT3BNuOd
HFQqnVtaElEw1O5njMvAHBz/12fvs4XiHu9pppRaNvIy8ometz6BHwHfOYb2xQH2
Osmqk/wgyJj1KuMZUWA4eDdF8vQXDdjuYjPrVOCFFIras3aiQM+bHXdGsN44vKvb
FZoBXxwK6qrc1TjxF7vTyK3YawCYQ1Cl7roEnjBfURH5/iv62Dum7hO5D6mMAvoy
xSKsuHQ3h+yyiloga32uSZzLIR3dC046jgCxHJUFlpNOtMCOLA813JI8KeoL+teP
t4OAX7ve50MBEARWMa6cznobaKnUJeDhHqB1tW1nS9EZ5xTEMMXtpPVA3UNvmVkK
BYTWCTh77m57MGjcDrFs+e5jGkupjeB9kfUWlkFVj14BH/993mchcskdkdPqttpQ
h8lqQtqeohlIUOiN2PPc99Rilgtt9/lsuuv1/OxGEf6gLiYGs//wWXdRwmO/hJaW
gxq50grLX6xvr0N9JbYaRcFC2ZHjxDAw6hSzTwnn/wcjkq9aX/pEANkNYVV5GZoR
7vj5O/+klI2fbIV/LAUho55N9sk82rYv+T9hEbpovhkmx4PwQ3Td3Ojdct9hxEBz
YAdgYI/T8xzflM6qYsoq45bvjlByoN/7Uj8D3NSsTOvn2wjoHGJZnGMpAMcxNANS
60TlKV8HeiANE/OB+wClWivguAB00KN5r/s02lrvEi4fFE3gfx2CIS0BibkWh1fW
ofhL1WKMkzxsdLy3y+dMAkmvJSwcpN3A2NgyOMhG8JMgAqezTcMUvTnXv0v2Y0ea
w58ldgGK10XPSM+TCWdnWNma7GHPo2Et2YGa2fjw+uGYwGBpC4LfqAJAFhnwwFyd
Y9IF8G7+k4rsrP0/OiBaHXVfsIpdrHv22z1TFAdaUAd8qg62eqUYEk7cBBG3qJWQ
2oslEv0T537tha14lMORMDW4mTXYjZMOUxjGZNWhWsqLIVT+mNw+I4cVfN/xdews
dCeQHVC5/wJOLhx/A+fMDYzb9Tcg/wsqP4rvIEYBRoCJnFRwQMfQOjzRKQ9fGHKR
mvEgfH28vsWAZfSZRjUTqFP5Semghwhm5Om3XX4/tQFmAZgX5sXSFq/7PDwP1V3N
CMrM8JAkFHvAMp6ulwarBdVAc+wFQhzFdc7zOiWFVXlzoNntnp3utKUDCL/1Mxfi
tc3CmxOW5aITDR2U/98hi1CHquX2NhBo5wSrEUYsD4j8w0eTwBLBGOKvp3DwoJK9
fPY8NGoMw7vmk8Q9MqEb6nUA3zUfQDWIv2bIc8YctVTHNxUBYSrlHUbdqDrIxthF
w8t411B3AAZsMfcvindOPbtVoaxdZRm+q8GKC47/y+IBXIJC/6wIQ5Qk0Fx0hn/p
Et5pK9WluOaEh7vuB8fGXt8FHC4zW3Xnwo//Lx2JSTfmqjQMbYOeIq9H88sQ1bkD
OWJrsgJNHZVGxhEoaylDpfbc9NOgctw7OVQVYeUI+1B1y3uob/driUnwhq76njfC
0CeRajkUu8BRnLjYc4V+YTZQxv4PIdMK/vgXbECcNdhebMqE9lnP04xa2xuLzGwT
NIgtZ1X0CiiGpgY572KYLIS41CwDWeco/nLGNYEYRId2S+1QmMzfM76zuDuBbbhL
5GOySkKn0mb2GtnkquByuVb+bIG1fd8FMSsHdu+VHFAe+eBSW6cTCcG1kPmDSoK+
TRZIZDZo5xoIf7EOkuzHd811l8zgaHS2GA3JrXXpMY+eiBaBMVhiLU2mItkZsCEj
VQIm5KHSp4e5XcZK2JUw5tCMUlaRlksGXJVa0pmGfu3GGvzRmJb5e6QBMnS6SE6q
OBKNzRO61vcOscugK7xtE/iYWrrRDjf7zEh2wVxNOfz3SJ5jUoHeR0pMdtEBcNLs
36EnxVyLMk0S1FvGul1HykOG74E5LkuS/S6zy6Uc9sItDhYTSh6SQSrTgnyaQ79n
So3KgqTeAPGY4XSl6TskWcM5lrX6qM7tXUajz/wR2EHeUQ+3vfL2tqrBCwR3Dont
XboyiRItzxktPoV0Bda93evSlJ5/CQ76UHKvGw5+X377YHdBee82pHU3p5cW311z
RFhFVCHywrtM+aW1EqpKKtLvdYsZhc1MannOZ3KU9+uVgIH0q3UGWhvzwqjCI32Z
ML6XYGQSuTWRF1X+PVyfOYeDmtJt56NNrn0XSZaVQIGqejdJFL2sRT0G+uYvIxz9
Ux8mVV9cYH5k58fGhApRxOipQWG5Fo3JccBULbTF3byKM0Vak+RjowE4nPWJgd+3
5WyIEYD1PHut7ASsFuqyx/LUZzT4wwwACOdk2dXUMMlv7YzpFJYO5skFSxj7PJ4O
0BZK6rSRxlpjLrSqUoUOL2kQgnPlOh8MKBIX/VOWyBAkj1N/mNm3KLvwTGFoIWAo
crXUnIDRb+zKDzKcb6fZ3yyv1wdv4HS53cbaODod6J1vH/YAda9zk9/3xkINVuuA
BHY2xAvkohtT1WNi++nuKAsZAmV/DWYLP1TwOaBCva2aJ4/qqmngpmWgbv3URfD4
Vg3JNvuov+rsu9lPo51hyea0wpfce7wfaaMRmkiefli++MbwBm8hlkz7Wvak+8HP
wBfj1ppCBvwWMEURGvWX4vM7JJeRfz5mMiv9OOPx26ghF+wIUoz2nyvYKcB+OMpR
s/7XCfemfiXNFTTElAQjN8Dlaru+O2FMRnzx/OZauiGloxA+xUgPSV/Gu8RpkbRA
dLHFkrKQvPTFySLJPwm3OYq/t7cceZK9I8yBNz49xlGC9UxyOaLd8KwSipIzOaSE
TTay+u+/1UKzLh10d5MI5gMXub+/Ws6dXYpJIzE95gQR7beK6xvjiJTjgMiHCzgn
Oj7Gd+bxExsZ0ZLRRvTV6QBENDORSGoXcr8j/Zr3fX1fGNYFhk/4NtmmuMqhbJmT
GBVapOOuZ+5E195F2i0UUl0bKszZ94sTz1sXJ4QrVVYu8JLfmqNI4ArWLP3ne0mp
pHvdKzhLL+zeM1k1/nHHGEGeeOcHVUhOt8p7KtvYAhn/TI/77Y5gqeRYnQ40ykct
bAbLIR/0zgzl2g4h/W/g3Ok24abW3c0wOXpm7EEeP0I2AzxGYZvA4jD0ZUEmlEfw
iaZrS4SVJm5iqv1n8tO3lMcgbDMfbZ0pxtJHOG5kryxEkjS6adw6YIvq7si4IPlZ
2VtvDS9W3jIrhqNFyQJSRjKehTYXEQ/Eg6TsTIgDuS3DfblWW5eZDApxth7FESOC
9bPXrL1IuwC47WCwGm+LnrJHEKVvOucPtyRdXYez8v1Xs+dMjfqRHTJCIEzB+wJh
QuukbyPMaWAf392xBJS0gSNQLr8XggkYTSQrqsrHNrVroPpsP5qXIp4XmJUl4o8B
dgYCKT+6ZXjF5MHspXXEEmvESbHIMVYurfcYHNAVyyi43OCjGLL6Jv9TSayzTpS3
WgGAmX4gYXOb6UVcqZ0HZfvd09/k4BROk3SjwTtnGU2B9v9Ton2Rqe2KSgaSee3n
6cUXDCPuwvmFauZQTGqmnOKsvzGqoBf7KDNToK/WnOjfsX1X9ncOvo5O9xKonOzu
WE37gT8YY1TrqdX0MsRciMr+g5oO8QYFhf6i4enyEHKhPMIN1l0lrLalI1FQ5d1+
FoFziVGzPjaqHu/Q2aLzYfSijkAGk+jcu+BQj3b7p4MaVZ14JEcuMbulKiwYRycV
iy5dLz4tydwf7ra0hd9Nu0WG98+q7Lqgjb4ei20LhafRl3b8AHr1Db9UEioSun8z
3HS6oYSvmtYultTymRYXhgXOYSh8qcXsJ3TDEY9bR8q0iJOjYok4dB2vUiuuXf0K
NGDiodKnTbPqtpaW68cWRKGg8hwF/lHto+VfQxkRvevAye9cos4m889Vl+dvGyLW
+871mDJP7e+6wpXPnTHCYR5iX2fyW+sBATYCtytvx03gcoMO3SbONZ5KhmaUSVW7
ygtcPzCgsN8UHAscjfA3Y/I5GQD0Fk/rKTBMaAZ+if/URipTSy/DRr8WW2jLcUtN
N0n2uKJLsgYuor8QDrpJMi7Uody5GCuFX3QfYzrXtwoVos+uOzPwUYukz/NXdt6W
CizenXHjq8TZn/mxbZIxDnb4upkcMx2sy+cMI/kxkdOMzJj180DVVXWeRS0S+t4Z
IsioVQ3yB4MUiw1ClKYVRa42RSFb9KKFaHltY21tcpFxZRpYan7uv+DAbi6dGgQI
dwCnIM1mFwviKr+ui+AGrjE97eoUcMmUjqUsJ1zOIbmx3OKvvYIgQoDDYuDcuFWC
ancFTVkOxfgH15UnDWKJgJKS2NxsYkoMdUzUoDop3in7IOWbOiHlTKB7sa/mE2DD
kWGlzyTKexCzo/a2bimXX0SmEBGi9WH5g7CwaeQiXSOM3K3ksDjiizA3z5XDTqDh
rAOjhgCN8AsYJZ85elXWSGF0Qp+mM/Qs3Ux1DFjIl4lmLXiHqDb/zWQmNlFBbniv
Gi5Hi7f4lXzU5McJvLuT42/wd1nX/65OHAIXZWTI57FMbGB/O2c/8Z+spOtPgBRe
pcU0Nh/O0WU2mibDRUSOzULPpMirJRCnv+jur+J0Ql88sSZ4nHnazaKzzxx7Iazt
iBpfdXIfcbYgL0O6M9DPVhEcjZwLeXSxFKkCPig6GVONSonAmT0w7mbtB8r16K2Y
zDU+ea2EcXU0jNZNkr7RJhTjCG4yJs88Ra27ey8Bpr9wSCRih7JvLiNXmIXygOop
EegQcc4YefPYn/U7ZP8UHGm9Xxcbf/+H9o21jDqlWI99oGnKmEIfGUJWWxP4vFIv
FpveHFiJ8fqi/EeiizFuG1GIMzbyTdMf3yQvj+/Pho2QqKuAO85CZMZMNfz6mB6m
74C4cEG4L1MzR8j1HD0ki6JrjSmVhfsqNMVqRMPtRRSV8StY7OxKmSBBVgHxeUqz
YbvZzSFSXLd6MYUAk773bQsjSHDYEqKjqI8B4l1BlzCBAyoOL4lmqNoZQDUQ37BU
3ETeWwy9O/FS+2eTWf8qw6I0vU8nkCLk89hF9K13niHr0GJpkS10+B/mvqFTYCJt
omvCWkW4oD81x8LdnEkPpwaNhNCTGpFFAwujL5NqZCYOhxU0zDaUMPCBPbSaLguT
hoSsi2pdU9U1dcwscmMr0W3YETkWdxWTN/VVPgSrNLDkxv5Nf3ryxgPeRYvD/Fes
6jrzqu3zh9Sh5wLzeWJPT13sMhoHx+a/gB+W7RY9wO0cWA8gg46O30H2vTNvAN5L
UKW8nekcdKjMUzezIBINYpZZisUfzAgQtc4+I2qbDmV7XegjzsGMW0iYahoF5co/
P6PFy9ZeiyiPNwBzTdcPRjdNhT3oLCjhmE1u3KjgIf5cLtTcXeX+v0brFvgWb8pC
MXMi0NPMCfrbvp33JHm0qitBWPoyDnAOmNcibDVYHHwGD17VALy0V8XnxGYoOTZB
nWK+nFWf4udCChlzkQadI8ogeurtA+AFpRNCGHYf5t57TpOsNmBo6TLl7y9AhX1j
exMeuXHFgCk/fAuvbM0tWiNAIwgj9g6Jw7lI+FQQCZhlHTlwXV4l1O5k/89xGYY3
jvBasVKJ8DCe03PvUEM/NTPI4JoV3u8OxMOcb0ZkWTsEJ+tRah61PPWAkBpvT0ny
GtpdBGiB8QGiCYBrzwukI/o0lkPMc8QI+sv8Nfq1LMqdcxnRSIcS4Smo8x7YLMKy
hRaSeO+ZXfG3HxRwg7CAy6jT3KHO39ZQm8FmYAOJY3uctghhuozmOx+DraEjDR/1
vONcp65G5OF0RCyMRMQDaCYHtdocYeWT0AgkI5s0ZiRyPWBEWz+PwKMPrW96HG2X
RRnHtnpH/15smayD/105XcXgqq8sYrMISqkS2T7oAPI5gEvcstKzrfXDrtlN7efE
AcjhQXFpjGAOe8QkSPRs7kf3JF2ULyTq0BtionIT9qYUiWGYSdRGacPWsDX5pW05
3z3mkGADVRY5Jd2mDuREWKKW91kvA4ai6OlwaMQ60terG7fjAEAnadPRlPbGex3l
50+KaHFGdprRpDgz0VgdZbS0azsxOuXC3YB0QSUSKLj2dOTO1TXAirIB98poqLSW
g8lRi/7DZEMpe3+pr6/6r5Zw+y0aVgPynlTMYvJ02HYw/j3JDYmu08Ys08ZsruOD
ur/0cSMcek06IUVHd59bHI6wRn9j6pQOk0jc3xEdNfzrjP0KJSPDZBRpF/Udd50/
UrTnr7SiEJ6ozeXUUyGipQ19qUicrWFhQNF+M4vbwyjfPTdQv/zOF95n1e+FIzFy
S3Gvs+oyHZ3AOSKsfR41jOUfFcpifv0di+33f1AZ2hy91q3F8goAYFHaxDE53cBp
oKdK6Ki6P6tUYrKknRTy7FtJsxixD42EffMJ1ZIhXOn4GwhMC7mrFcF42NTi2fRU
qDcea5Mv578odORaY1MVS5+j3dxSb+eW59FXZkeZs0GYzkrTMQy0enQO5hP0aedd
AjjDTk38h2xxbGuaQhgDpGzHqsbhKAKgMpLvXHjT8HMHuEC45cVIle1z5k19/We/
55D9Ikp0cn9tul7W0eI0UuxN9+Z/SQTTxn6rp0YSErF32Gt39ASCJvi2Q3AGjMOg
+yahx2gN7OvDi87BkvL1ZKDe+FK7fi6uiUkv1zOfE0c3C6h+NwsAanOVOyYbbOff
soLLDpd27sk1hydF7zKVcbWg7PArjA4xCHXqFL7U1CdyYUlKEruSpVGi4ZlHSE0M
CwT61hBH29UVolk+cvhkYeV2j7GmCCnG8siK2Ar9Cnh7HMfIy3s5k+FcLGt8bEuX
/OEBAcCa3I4M8sDjKISK44oZ+b9a0G6KGGQ4UiwVRjr6+KisgRbwRZaN3+xRzry3
dccwHoa2sbpWeMearV5mEy567KGPLA3VDRUcEmysw5WOlKHek8hm5XvIDM6dLy9w
XhqkI9cMs/1hMI3pGHssPJySdMV+/6UhL0pdHgpsQfMgi9ihBt63YSU0CvNXk94i
wjB1sHjyAe+DP3PP3buLNb8XMAEQ6xB7vb+yk+gC46oyVpiWB8CQgb4AxGSGYxDf
JB59rBV9ANFVoHbyD7ITSN4N0/nfCw6KhpAVE9D8FbawkefK/mRjWDIB1WvniYjR
UhayfGBqN4gbHH2SexBAChNBWymOqwSDmMAtCi4T2Cy+vjXLMYmK9qrp1CIEzZli
fDLr2Mj+QXg4aj4dw/etsmIbfs386xGJHmbeWpNU0fZq/TV4iB4+FltAB87peGTr
AVmySwo5Ihf5MaP7Y93C+GPjh5VpFeW8r1aH7usVqD3QHHtSbivDLorSpN2EH/6L
j2Lj+usd05uwtqkoTyGXFj9G4u44Ox5JoubiBOLyhw4AsIZ6r0PomTwXqfUHkt9V
n5txMfvd7+UssGGKoWsSuzDX2zCXzMxYeO5VEncKQsDSFyoElySAtLiiChw/AGcr
h0QT+kDIyDsHJmXtCBXoNae0qWocdAWDOFHmvMyLLyETMAUD9M/N2WHLxmy03b8d
35jEjl2fJYPyYk6riLcX4Ztgv+fETurtmH7G6wvpbVpJn+QeI+EZDG147FlfV1lR
zOARrJEmALjRprkrnDTpqL/7Kd6wmCeSvVEOmfAx/RkL/iJjlYiRWxBuoY2/RIML
D1Qf/S1SbUhorETnjiGgZGVqlx4c5+6vXxraR3wmfNYWD3zzaYJu0rTFGPBZOVlj
x9dA2HLyJS9x+pzI6MyW7ZTmoLFzIFrA6nsqTlL0+HVsdX8pRrbeUIsA9czubjzS
adKSg/IGatoEpRm8qOnpeW7Co4z9+tl/5Rw0e+4agylNxS4rJcCYE8DDkxXjpi6V
gx1VJJ9iHH2zfErh9pWP6E28J8liJmMPhmjTjSwT7pSTriKM6pmZShrJM2SL4866
D3OvrpExLZxCl7dS1uAAII4ZY7elvY7OEpOGXXMlXLJt/qDqtMQt+aLcqYYeMHaa
Xh12r36+Un0GAXKQV7dGWpNzgJPwArzQ5tTswdKT2uv52fE3dXJ38v0+czedjs5r
VTG0tgFgET3oBVlbQnjDMEkrUUdjjBuyDgd5MhElZ6rzPMIT7MbYu3qhHjDyJVQt
O+HiDd3UYkOxKz6HxmeIZateASaAV/n3eNjJBvF0FxPUvmbyzRp6oTFjpC1omDYI
okqWyuDP8sSdmx8UksL4KeAFNWD4DKIEAdPkKNL30CXeXCTpy8WuhafzqTov5lPI
8ufxHocAxQm8BXDo05ew24Bf7lNXskI+p8+1XLbo0lb93AhVqSuqcZS5CzDFsCM5
ITilioqpUMvqPS17hzfeNij7XwvR/4u+aEGbCBKK0yoBe6SsufcfBwFVAbNDbWHZ
lUxhNiA6NFlWkHEOKpaPjWl35PLtG6XFFz4+11npDnRxEmB6zp+hSXhcNPYh1szh
/9zkpYEuoFZUUAiUz9PKmEVm0mrYt7AMa11qPLlspamx6l/xLOHajygw3qPZCmCF
hceEtKt4msnbARAx3F9QpdRQVSUPTH0LLvFX2j3liAOJR/zDa9V1yjJrzHB+v7y3
myDWjdfK4JCYE5k68xAALVDsTtx18nFbh/sCjvLwvPPTff68+6Kl/2vu5MB7YMiA
Rb7RaJFoytniDinwRdTlSMETANWy5hJK5ojpfyRTvG4JM4nuGQa/2Wn2BRcN9KVt
pK8efqIlPPH3MlAjvJog+3YATDUTvoTSF1kcn00qcEv+Sq6zP6eeWI0vS74fig9V
MuLA6jW/3pLGQTwH/58zZwW3LD5PhyTY3xR06PksfTw7+oNQhlc1BFOn8XujALAG
mJ/Sbsabodif9FGyXZtNbpBAQ498tA9+zAH75xhc751mApC+tzKOk4R2VLR/LlRQ
oWwD6HrGeuupkzKqN2Mhnizy66BIln7OdnyB5x/6aAaCfN8/VPSsqHHOSCJtnRjl
CltI/qQTLLHh/3dBAuGzBMCvDUXUpGYLOKznzPDwXwyPYW5SAOfj8IrSUzTLD3/B
TVw3lPcwVIlaBYZhNKGaNJcshYfhlt8RXwg0z17PEfGPYWVn4eEWmKlmwr6Mdtf/
u27EbdZLR4/sRthX5u3UE2gKcanOpe+beeecyMOh56VUX2O2PkRfuRbGQvpzJzDN
zFuPuvDITMSw5NMhZHPGcY0jIV5pamoPbtyepWj4SYQsuZcAvydzh0CIzIAxx0q3
14gDQxdYfjotxR99Z0/E0tfggFSn1pe8QH52PxDVJPAjvGBCq7KUj3A0BYssf2K+
YS98mvCIF4MRrps54u561aIMm7359SrQc0iaxo9wvcn1O4F6VxlXxe7nWCevgajv
K4Bk7gBy6vzy6nRZBsYWt2ugbX25p+1YR8OqcJzYTp7HOIITJMDuOAyEE5+e/mGx
JuRzZxGGl4ge9rL5rh/L21X9Q8FMFH53Yw1zwOVSTsf2fVCn18LftYmNhVxe21ua
4fIjK664UQrlq3nI2HTZfPjDHpdMwXrxlH5LlylbTLHI/uoJNlRpnd4DaPG4cxQO
a69k9oiIQ9fNqieOYbpitwPNkIKzZZ7XwbjeqJ2Rp4QipLUpVOTScaPtjnOYtvp1
YhqD5IbagzdH5X0kh2w5LZMXAsliTIXLFrCpbKGKvcTAFG37d4p5k7VkUHV6Yvvp
pZpInwH2gm8CaBJzQGa0jKy5OrhJi1z19RNP9NIh/HXSKDU+vtyBUiPt6w9w9O27
GH+7G+C4J7OWS+EU2VsiuuflElQ4uTrKXDGVGU8Ic3npApOicMbmk3HBQ5GxwqEY
ulEGGp+f0h1aZHurVJRu11+2PlaPktvu04xgHLc6vHDVxfjxieV6AqdtTz+GjeH8
eNURTHWsyfwbDQGSuxKkBbNxGuZoskHRDBY986w71VG1ueOdYX4NdQ9GvuR06j/3
iw5AOCd15p9uasEXcEXkrC8YccPT8fO08/RrvJZwzoMxS8Zv3zEzpvTbDT/3vQZs
LRI01Cz8goCkv9HUBoUq/HOGgmmXFv4lZa6ooE3agl7pXdFioMR43hLvpRYWbiK2
AxldEw5nlxn0I2Bbi4UXofJs/mxvRUmXoMZitQB/IM3JKzpgk/mrJeEfTdz3D0B5
oysHsoFX2+uNaqBU9BxmR71brzsFKeWGsotyRP06HaQ1FLAQheAYl3ID/yt73fiG
hCFKmAg0jdEAvJmhbfj5VAVwUpVrosTnA1sUmZ7FlzZdbE/7Ui/HBuKjaKBCt8jF
Fnv1ySFstxmmpaC+z/S7QE93NUJFIP4pwGng+k1kzny7/Qve5u8jjP+nefuBMo5c
EI8qwQZSVQqRzfiXv+syCCqQGJJvA3/z+82y+0iWC3tyz0uPzg7cXQzLBs5OEFSX
j7jDTIec+hCffoYZiSmWUYOAzARDrUniUkQc6fhXCvRfBNPvnchW97vmFSnQXToz
2e233v/8mRZdLcyYOk7cTTdztT+SQkQJFdu/b+2gfmn5Sj07+MRyFqE7SlBKNx2B
jZI/P9zURdxQxSIX5oCY5YubRihLTZ06neHfBL9gRz1oNGMfV4JSAh3BpwICV69q
ErBcpLB8IQQqAHKbKHqyF3g6wafi7A0+tT+39Vq3W89jchmdbUQbL5XfmkStSBcL
wxgqDObLFfky9PMaj7W+O8C6xbAU2puoje4ezoUofDno2wVFg/ESVVaNUteZrRKk
O33Vq9MQdnwfN7jfxLg8YmCI3k4JmKl52nypnWJwJypVh/KSNCLCQwshlUox/8WJ
/cNB6jYyWv13abb2r9j2MUr4nbJ0MKbGhWZweR3x3zYubh6B2OcQsY8nhOTt+7OH
MNDnjtRpbmnvVAK6LFdLeambEq6ig0EPQ1zl3/Kb5uP+hCU4NB9CqIJs+Jc1htYH
pt802cBzGeisJ8pbekVX7/o0y/4JJ3HywL86k8XycZM2VvHCuORD3BkkRRTXfUMl
RIDB9b0yoWc5bxBEyR0hLgGtFrYmWp1iaWBautQph31Xw6qnwz1RnxzvwdTDOtCO
0K4SkdBmI9qQA1moSAaHUq2iPNVL9v4ImtcKeiKM/5LLfycsCEILNY9uhZ96d7cy
/r/tTrt6+ZG7n7xU3X4+E/QLfdUpakC44vLG4AUJ1yETO6CAHdHXxBAp/u3GQY+s
Vl6yeliknkmMKkzvXol1DNW19HcsUDNQDiFIU/YdUAc=
>>>>>>> main
`protect end_protected