`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yuiAF2djpiMVQLjverTUdFCFIYXCBmhYgTqYKX8jtGWEyoPysnKDHMmDo1SxI1oS
q7jVQyFtflTFBlUE01M52Qh4Adrz06pzXMEsdNa8oMxcoL+NaQw9Iqp3TmMJmh7L
N6SnhVmXe3rYitUM2DH+h5pP5UPInkfLy1hfDJUP2m6Bet3lVK4gWQY04Cn0On3k
gY0fDabph/q76MNdOjPEPmd/zd9LUYmISqt/DQoGuG9kp4jJQhvcJVosXUs6kSzu
m7iDSy91YjfBo6wOFs++vNiS6mkSjhuQCQYXYvwK6R8qds7w3E4wmfOTpxiD618n
o5doeWcNB9XT2lGhFTOq1XqAgp4XKcdIJaj4Lu3ccYo9SYng5qZU/8IK0KoKRvLU
wmoYxJD8Haeqb332DD0BF/lOku5fhCkKeJ7tWYXSxMQ6wP7q9UDGt+fGnBis/VRn
QKM22bht04yjpudWpc2TH1GjGhTdWWnYRHgM6OG2H8CiIgwnipqAskLJdAokC8j8
1DfbcrxeSQiBSEn9YGvvYZihdtRmBOsdz8EdZEk89XswT4Bgs5kT0AKxUFg0i/NU
YS+pIz1F9EkvxOcveEM+o823FhUHjFxWkKTmWR9Mma91q5D23TSwzwxamAui1Uud
77W2aYvAfaHttXq+UIqRVwiiWPd+UU2W15VkO+fbE7uPFRnd2zEDi4hb81ep3xi2
FjTXXpA6htGgIi14rV5YNrrK+EhH6WGEmVLXDlnDIW0Kdhystlivt8vXujBEx/D1
uvYO8w1fgVmX6ro7gOKI3ebgiSICxf8FHpGDiYFeWcBYjjkBIBWpd2h4wayRghbl
6VWxcIjfVI4yrACJbcsQaIAajvAT40K+Z4Kk7R4JI3xOmFMWQBu5hEan/B50uBrG
CXspG2XuD1t5KJuGWoe8bo2Oz0zHTgaaFzyXyqNlf/h84pQ3xeDhuU2dJtx7YqHg
YpLLp5+3316dJXhT3Kvdd8fiw2nXdaBViqzhjNYbeLUGuhkJw0N8ea6epwFZpWCT
1lcEqcUHHECqIwA6SI5DTtth0yy4PcyCIm5KJlJANW6bfgFf8z8XHlz4yKZNUom3
ecEv2tywY5UJdo7IK5qEiT1wIATk9KRsoB2uKDDuXKMt3WyYQMCKKu2dZjBCpX6g
kJLicwn/7U6WA7amPE0VlgaXs0JCk0IpgTv053WNmiNq58Ljuy4qsFAzGqe6sVGq
8zsBvgGeCT8kTB+vjPwTDQRXzsOKTXgSPdQg75IkVFuxGV4ELi9pIa9MqogyHs8V
xlU1Wr2XEL0fqDHelOB3QbifCVnYbJ+6C9DbOWMBZ1VEvH2GK9fldmDwYKApAso0
NEu+2KCZ4U0exgmILnqe9jffvdKV74a309FQEH87Stg0rv6zSY7gDt2SJC6Slm3T
CHziQSUp/iAgJXsFZ0Ws1aDSymbOuoL8H3izgl5mOYebwuFxx3y43uPv9Cl4P5tc
cZFIDYxQF2oAfMnKM0lghe0UIm+zTnREEngahcmmvTRf3KxG5NAagBDdBuyp7C4W
qAmb754rnaSuDh1vTA0tFnRzA3ntKrKCDXmPDC8CJXR4Lute0wdyWqGFm3zNslLx
ArQWBpgHXvgmwa1utkpc9hZObSriExHFnS0renLV6JhqS2viTXHkoAFSOummNajh
IzPIDSFNqCoXRmlDu/eSRrgi7QFNym4/szoJbj24YvTotyOQ/j6ovj+FXTwYrSN+
APKz6McGX/w3kqwt2Zbt/c0LHToqiBEiGnN4p9cUy2rRSlJYjXp0iDwGNOZKwFsE
YUWrA1gOXcrIcgehIWReFMVnGUd2BIDYKotRzI5qKUA3hyB8osgTGUKricJXyBnD
tQ9fsDNWdt9tspLGn2Xd3S3Fbt+lYZSG9Ceupx97dsdgcj4I3X0Ry3CYeTHLTX8y
djlSMOVy/S5v5e/FIlxs1pGX1+bWGyRLCvGPZRbJBbPIdjvpi5gxNGDI9jkcAieE
FpRELQ2uayrgYc+Bguq4m5O30xAHhlFxztLW78kKfiWJ+OV2nJOBH/NlzvJ+hbrD
0McLRMHZJrbmO+2/AGBlQT2f/cdjJ0TWMaS+HN1Ew9U9awYNOwJB3k0T/mhGblMC
qMz2Gpldzw9FrxH+uKcFfn77Jj4PscsbdjR20QDhlDT7hGghr+13pFRMIUVKHt/G
EHD5bOzgTo+3HoNznjG3DYaBGep3EqY0ya9wOrURq9aj/CDwTZPwGkLHYZlw4lvF
OrbXytDlzotPxkxESoDXWx134Vkwuwmju/Wx/abi7IMaQp4H/ed5PJqzyZuv8Ltu
TEpXUHMvoD0LbrR4LalmTRz8lO0/UMiSBbLOBTZXpTrgTl5kbuIQUtaVdwfQ3eSc
z2RNw5Y8WxJ1K51P+uLtBVqCaeaUAxrPsurRCex4RCrevFS5R1dYDLLW33bq154/
aY3dP4wyFftYZ14f3iHqjNrhA8oJ4feU/6F+lk9u2BPdmHlosviQnv7Y4Wuppmmc
nlR4Qh7jBzc7q80M/cJsjlS2kddYMiISXlVbLoxUjUan644Wo8AuOQlNbxwT8eFW
sUu0GKKFfnj3tToMIZ7plKyFkEUgGaIp7ekBjXMPUvzD/ApDPlexN3XW4Hu46+09
J8iKM5Qnmfspr4zXJ7RXaUBUGuckHVo3Z22/IiIkPKJjRiscUrVGND8FBvdh3RPq
/dPdScR/fLSwdA8Fy/KdrZYjXI0bZE5xoIV5R9XqscZcSDM7u162V0WbEXeLePn9
o8Q2E4erWqZsovJyBYrqskC0/j+Kto+GeFcOLQpa5Fc2/3TiZSYNTknnC4zRgCC9
5k3NklnWXB2Y6aQRG7YTIAeZ1Qk7zVkHUI611t+DGPt2rHl9i4/xTQJ0mfiw2NMm
J1wgbSe3g0DhZIukM78qCfQfnVeRB7Nbw5wisxRVcl+uQBn/djp7x/XTkoM7tLeR
XElWt2jlOJK/LZpLP15EgiCuVlfJ18Gux3lO6kGBX3Og7LXZNHQhbaBwm5cfwHvK
Zy5hLr5iFzizM2oI3/15/iBRhHQ3xzGA9C56BUgikANxJzdvAuspoytve17V/Yid
KyDDYXuwsl461/p4FlreA65DunNKubw2aTB5Yv4YbnF6JoazSzY2G+HJdkMaNP9g
u7A9Wz2wra9b+/zSgqegU4Jd7yxjLd7xfJCJ0B4iJh+YsrT3Sq592FTrMWcBav41
OyHcXZBYftBnMVnAZmN5f1dig19F1QFd597xL93lbZCDySfOxOdCDCVXCUM5ybVj
A1FUM+grdTPEPAp3P6U9Or/O2rxGXhXy35ySSGTtd0SRIe4TJpZbhrLA6nTkCbmE
6uqLqFBTTqhaHVMmWkPtNHshBQf4BnL4QdSiHrVVqBdIg9ZmdTAE8hBcH46NxcAZ
kkaGraPjqU6uOzYTRMNK32DRg0A+6DrPuCMA6m3aSg17x3hN7v/NKECYPovxFQI8
LFqQgvlBsbg1YDXL7dSZxclcBQN0ukahmaJB+FSJS8yveU3WvIAmANhc7fujgkBy
YdriWayRjMlVzSJLxDvGB1ea9JfXACDaZqhAikvHL3dO7RZcNdP5WlEsp3CLmCUV
ZmUcmpcGT/rKQBrQBtdeSGrGSD31CIHrKAnGPCGlFobiEQNJdsq2xbHZmkllC32X
PxqGbrYVvJOAn2B2vFK8XHs4TQxkmGxQRFEPE4hc+h5NJjDsJjd6A0mM4aiasXDq
fbx7KMc2T9dzqpLZdD7m4/HPE6uK3TzjaFKXTEaX6RxyaLYej6IcGha0rJGTtfoa
Y6wJeaaWLYEUTgMgYmcterom4ow2TwYPC+IlCrBILEaNLt2NoQgkIqhqXrLw34zO
0jeBAWy0FqcEejo0VjuTmpCQz2sRiz5mdoyJt3mz45QDKVL6ynK17zHZxk3XdU+z
ZtRnsUewFXpDeWa4faemfbJNpTpxDtXn627Dr1JQGZt4Xa7bCIZAA/9NF/rWiCiF
c/F3sUD28DoWVE8sW7kyyMzV7nOw72goIy3cwQQPhbqIuIPlrwRde/pg75GoNvNt
JkWOVGaYtBhjDlkFiZDSH17q+isocwhopwTuZTo81OSBnrodPmBcFOGLztWKQYi+
HqYlvonb97Iav9/N0MQUnh1z3X5pifEEmLWK9OUfRempUGl/HEo/PLJ/sOjeQQpV
Ls5qjCGYJRU4a8fyHucfPB3jyd0UYmwGAPfok371dKN+0N6vfg1k9Be1uyDs0NZy
GCgqRrb6b4VtrV9/eVlSjWHiBo9oEpDkMi7tFDD4U4a7KKLEyltKyBLEVye62tYE
dlVW4/gb5k99Q/t00L7W9AFzWH6McwsD/C25VtAHanDA74stnP2YCbfaORb6Iia6
D67vYp6IoqgCfHV2J4hyB0x068kgPUn8cZQ571ngmapTsymaYaLwBqTa6PmYDvDd
e3lvxzzn6/5Y1nJbKBuXGg6KfnBSrfC/Tq9BNE06wme/mUqXxSDAenofmaa39/jY
/Z0dB0TxfLfKWpD6sjdnU2ad+4p34KSqXXRB6sFpxOJEEIiadrM1kk6w6ekysrsr
Uzq2BYLVdpI4JvwPfRixFx1DzvX3qBbs6AGFjPhsDW3O0BElL5LIhY/soIDWmQYv
vsxJbYxuhKsOPVKm910JriN6Wb31q5JGi6chIIEzrL8vS/4qhZOF5G4O/FCLasQT
7f1D1hABx2r0mdy+NPdYGHHP+5n3ANR8Hp5SQUs790FBzPbx8Thnd3d/fHMVwglE
AMYDmhx9UQTrA/WQKaWse//wPRK1tsjpra5r4mEyJkHUOu6lT9LQ1wO8D3Ta7HeA
LAJObBG3hJUWGkQUZMGDruydlyYvoJLtMlJBQ0YW8TN+6zp305BBQu/esw+zqKPo
5uouZQGlsGceVxOHDxspbP44NiyvYtzaYsazFNCAu8nApq1bSLE/tSF16fzMubqF
`protect end_protected