`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
7d1aayJWrMXzpB8QUg69LEGhkdg8kTVcSgErrhWC9h5ktvf28mB+Fzkz7OFSzaZs
80IyvnCzp+zC2zh8fwuHo4COAY6oRjnq/LP6i3+HDMDH54Poimqpv1cbnyOG/d8p
h7FEnApMTB0Na6uLXNCyFr+/j0RVPLBRnvBaJgy/IIdLIqplmbefsjGGV6h18FkB
8LcV/KXBQ6YigTcr+36rpFlgYqD3a5TOUXWPkd5uzGE3Vp2ho1T4C9FFaS0Gc9hU
v/z9pTs0tGrsLBTSpvyLQUtOKmYtT2PYoq5mL13dhf5c9O8Sbd6GtDp3MnSpFu1/
iPlP+DSDf4wZTrkhclS3eJBzDXz/FtSlL9ti2ZNdSOvQ/5OIMJoJ9wg21DWvRB7w
2glXJ3Qv5itZJgdpYCTYa+WwI5558A2aCMrmWqhMkPR+vNU+WvZAH/J+Z0Qm5/oZ
1xI3Dzme+JIOEnpdnDhpKL77zgixAO2m+8C+6YasAB9Z2OW1pUP8dfreah8I7XLz
bSQqyXrDR8H6Qvj9XpGJm4CzTcALDqK8f+5IMc+Pwe8WbmT2YCLPcOdd+w9z99TL
vKgv+6IYBwDnFUGWKkS9t9e81ESbHHIBJCwy+Bhi7OSZK03KrV4KmqXRTX/Oglrt
7MHih1HY/pAitWT2zBBNjaRDx8EfBrBT36IAe5sV22D00rtBUIR2HSu2FDa4e/DI
50Kg9bR0ZsHFx2qG57cA7qpYNF7zpr+46JOle6Hes/Sj0bRZFw3Lbs1/b4idkhJl
7PwwplxpMQMH8+RAMknJr6ZIIIZ8BJGa7BIN48NJbPS+E4owMmLXYAVW5ecUf+Zn
k8xUzXulfvboFX/T3d9UVA3/ahpabTbH4+91Zj0wjqIDSaJwfXvUc/1O1adsWfcl
NSFSjEA8WOSHjapxYwVcAYiTeV/fiY/5twNcGvLZ2UUPodGaATyHNr4tuH4YFA68
9SrTFTp2wffDTKVd3z5zS65IRdXY/U2U/9wqMih9PWLuZgFK0fIELEnjThhJAY9M
tge6ZWPFLqHmvQt3aOdclNbp2EvsuZ2teoduVMAY7GdVtxq4HxzRgkfsVlbZ8ffD
xMuMJtXwXxPkRwzAETL34hkl/cNcINhhFQJLbiASE+RtRAaxupsLAGz46uUk0ZXE
iFCRbanBiT37cHMeyJGIqkyGjT1jOvsDao84LK8bfjdNiUUz4C/r5K/b0lqHQ6I3
WKrZzLl6aRcTDLTNS33yx+DnBWC+roZ3n+Bu9GPD8ZI8tfAE86dpZTorlelstNpb
KVxeZ4fdace/rx6LLVmNz9r+J60MwJAiFdiQzbn3nwE+kPN02J+xjQLQ1JIysRUR
dFWrrZDAWhDCVKLe03/wpwXTGitKpwKlSE0BV12113uvwDNJz/ueTvJHq6gkzgZG
DEvRc2xOvmvcDi458mkIHcDoCN4JoXJVXUyPsVe2c9rWSnvDv/VACyKnIcfQ66fl
+4khvbRKSO0LleMP9ECFT9PDET+TqIfCQXi89ijYa1GNvpFPGAGxPAhJ7ZIJeQqx
twzF6G9gQsYhVb7If/O8MHpMvOWTe9fyFnhmgHvFzbHocHiOm0hkzt5i3PsokWt4
4SNeV/k+axGTmmnDm75OqOvPv2e2zGIpaPVnXMxeFQLjCmvWjoT1o0jGZtNJitXC
IpgH211ML9GbEFt6JMecQW1TmR+yjWq9Hkq20v4NB47Q7Rs3XUtGyYIlwWl7NKWI
X8d+y23eE9LvIu0fUtsWa9Tts7hAOrgOxWME5hKRw6PbK5fmVRC65tUMVXWdEoSt
GU6ndhOXbfd3rM3c2yYCM97gvHxA/OVfIhRVc2sbA/rxow0A+8wO7Xb+k7g+dl6M
ZW1GAouIFAMzQnzMaH61u0HDrT3o+S73bTOytzfnRRfgaT6mjlnkd/e1TMnSnDpG
1slbRdA66mSuN467uLNSXbRpdy3PHk7A2/XcQqAIeekHjJgPjblZBZy0r+r3K+0U
pJ9mTL0bsf7IC0XFHhWzSnmr23ZFa28MR9ww3M66io2vuqr2X1459FzlzpchUeVP
CJLDyvIFnYJcLjV/bZXM6Ps0MppHGiB7pcvmPomfPhwAdLb/XgYbrs+YpWM/KhfJ
pQrNjsdsi0liraU48WMhp895Y17lOtrbDGuWQTjbqNhE2YErwYpyywmy3lt4TQtO
dn+9qtrDgvDhFBTo+TWbb4pbTtFHNlQhsy8GY02/032hvW+xsx17mJ8xPqnjIbC7
o+EyroqDD50vKSx9VLrn77YatOfPiSnamJJoYYwzv5ZALnKrzPan1iJUmNqTeG21
/yNA/fTN0/8Ecq2M4vYXNl8c57JXOq4/I9R8jwF2DIQH/RNiRRlj67yReggJkeKD
7vnju2UaHWM/kAzAJzn1SFgSw32gBJF6GT90JU/owtWdRbKyolexx4H4IHTlXnnk
b0gl9/d4qtLwoFZYt3tPHBe+W4Y2D2z6i6UTyr7n7xgxfsjk5SZaMYG734Xpik2n
Z00WGBFc7ArTTWG/Lg05xngBLRF/aFWv//BrAusZ8SdVnffWS6MqaNNp0CiU5iEo
vnwaFtCPIORmWfv+1dbx4z4cEdxC4dQ86Gre+25XtpeS9SNQAlEFRPucUF2ns0Eu
K6GUQKWEyTjpejSgezGlsSWHToD4FVGKcUGGolHiFR9+GGuehEBvySmnxt+Bj8Mr
FsIzRX4PtLSRMlRdTLxbyOhjc5UapZF3Cy//0jNWNufdhLXZI64p17F9R5UDqGMw
tvsObbU+nKq0i0sT2btyW0EKdAMSMGmw1dkuSM04H09p04FjZ42VwB7H+Eu+2nGt
v2HEVXZobpxFRbC6RA/Bx/jyzz7bsBCA/c7wZ9QNbwMq0B1q4qxo6WKACkxTmr8x
q1XADKUM9KIzaXMgD26FEtC3vBNCjxmJBjhmZTvEUwo46rOhcJSCmpLXeyMs4tVx
o4Q2T9AtrDZyEDGFqBSw4p8EhUjIUDVTB9c+8TpBjrZwne6iq2nVQaqqdfbHnSzn
uFBTZWb7P5xJXMqB/EoWhRps2c74gjx0T6QrVHygtjJRmQidc/7w1/1AL5VH6nph
VyYYgM/NRxu2ynLOTTdoN7y/RKmR2eV+jQyQDhEjdo7wZa7eCMVoHoi/k6ftLS3D
cqZsDvg6lfZujHEWCr5i+ThoTYWMsy1SvZBRRPfHxOCwNLc926Kt+8UDfDQoY26M
iPiACsfqaNHI94Nb0jiFwUU9xZj3Y0armBFZuMHWlsFstcxddRVQq1njP2VC8L/r
O3hVyx3eCjk+HCMVSg4p/an6d2TZ+ViSL6ustkBKxvMFyVsCWSX4qWYaWda4dAbD
0ByH16mtsiUbTRmRU0vnciHPIDyODQHXRKugk1uk6T008clD5EOy+IOT9TEPaqTV
GqwcmBRE8/eTN927ktl6UpyKCq4EnYf8jr1bKrVWmzbSh0N3CinUcUgzlIUr7IqG
sLEtxeHr30FhV0YLuxPqlgr+jE9CJXhU8nODqGrs3ClBG1LVv5fbjI4k+gNxMBcc
5Jul2oDbWxsO4NZ4vSw4E0RKgoFRtSi1DC615ASUPZ8CISAfjy5eZBc+75uGREVV
sln5T3ig/EH6PdC91jDDsVVWLlSRTGEKyS1DInbNfzyB2c5IwZFdEMdtqPWrwa0m
VwNJdtCIjDMdVSZPKdn3dDFJGSnp316bLWsW4p6Xq9kWpI3dNTRXM4+vV5UqXBpQ
mph0qzx33wp50ISaXRb0KzP5pduV4Tfsu9RW4GN8/gs5z/EJMwlR3TAC9FHWDEQN
1LrI1LnDDhuILZwP2qwVHVkpeoCj+GdpwsRLJn7tdqnYeJeq2/9nZHRfPmZ303O1
AC4PbRqgAyo4BpYh/OhPXH+L0/Yz/qfnqMNz5kirWqUdtQ7nndiC6pRHjvKY2vm7
H+yuou9C6hx9FKE7DqY+BNeXzL/yiy7c2hPADfRZI+Gknpknhhya2T3T9RceeJlg
JY5JPFRqU6XhQVEUmYIyVsr7AqJv1LAKtdgcPb/Xz6ObAP53tdgO9aTk3mJt9sn8
8cqXm2Xmi1xObRVG+9tTfOmk1gPgkdMHVZXdRYX1pA03AXjEFZqUwLw0v1i2mzBW
edCq4N2B5ESwNmYvRxzNbNVjceC7Hf2T85UYRebN0e36bHC4+ZCEwF3zvmtz+yeO
xFoFMQ01usxzd29L7VYcr/3OAZ8GdPjdWfm3k6Zw4oh9mDbcN6t+39CtQ28hulPW
5z3Q68e31BNAuKMrJX7izOOQxV0RaO7+8m+AcsqGO0kd0/lyNH7C9Og2rX7PPI6D
x+H6OKPsB1TulHhZ2sHe0cDZMCKW3+VNPnMJ0T9IuA7XnUk+XDSJDIrUokouN4Gj
BOLGTngcUiJyaQ/DQc95aE3Zr5a+f1zw5JX9azXsTsu9nPM+lC7BiWgII9IQS7qm
JPan4t/iGT2QAH+u7PFcfaRrr2AMHfKOee5dKJg/4kpmgj4FPuAWaKi+kCxO8Q6A
/j0/yEluYJKDRCN3hYXRADit2iSfYF66TB44NhDo7dLlI58OoFf3Vi+/bVrD2LET
XUW4sT78qY9hA9I7Q4kxkNpyKZxzA5JzmY7KDZBk1DRiatVkY3+MhQdr/esG5zql
6QBz6GbzsNsCpTzZmGnOxeXLTNS8aW/4ZKUCj8UlsXE0qvHZvN+Kj96veJSMg/Rw
EbJT10b6bfNrtL4Sn7kxCJozvxwek8POwPBPAGvTtR6AqlmhYCL7or27AYdKJrAH
Tv8I4JLuxYCfcIfG9IoWeoCNlWnbMTznNfH8G2BpUk5UYCoyXbwR4whXf0yN9vVE
buAtUns+QsMQBrfZrB8P5Ed6kBFDRNMCssFQmTaB8GNZmJzZIDVYgfNnwtMIViAC
hgSGQ9GfLAU97LHSLJTnPiSH3sXd0768nahL9dXmSbGWJOu1XA8nj8nyrWFQce4W
MbKJ86hXqWXpeh5fvX/d/ZQlk2+9UPkDpQIRGeEZs0QXXAUaHwAv15v5/4l9OkmV
gyFEKsBSoFVn6miVO2bcQiNVI1ANfoULj7VqZJki3zL68p/mhz+yerBZbV4VOL2R
OigeNdbMlsZop7I67WFD+3u7+VcZTrgnn4CzZ4vJKe2Tn99A06T5GflJRgDrhUYt
Kfkzfgqo9D4zLMlaT1Gs5VMRbM9ku0zMGko1/gJ08JEFgB5Taq3BXWsGIE/XGQNe
qKQmELsdUeEfePT3t4QxEad01VAVSL9KwKuCbxgm/GtHjG/AqA/P8JZPhrtMyh94
xbs8mV/mHke1J97JYR7anygsl/J1XgyBmfQy5WgSMXoKTksQzgs1HbL/S2NPiwki
PyEDPkzT8p9yy5B82X/cyTjbLXteF+fu3T5r5RVAPOpuGC+Mavksz/Famyx9gnMH
s+9Cjf1BNrXofuob4Nv8qWWYa0cgxkUhB8DD5+KUhG8hSazxqdYzlRYyi+V7N7GI
6Zb7YsIg/OYRLxnOa2pvVoml2gvJBl/jnjd2maQn0BqAEU0yNk7xw1MFKY/mK3OC
F1XRJt1WiKSUxZYyj4QpnLsOodUUylhcu6dXrXQ5arbhU+zNUzkEkFbPWH8+09Tm
gckNgs12VcdfdkW8nAvWnBlKXDDoCtnmmIEY6HAoPO22xcA4OV1WNk2EDBmEESTL
i1C+T6AksrYwl+g8eBSnDkqjSz0OTiO84XhINUjPtkFQu+xUw7exKfgbwvvHPE3T
8b1HdchPzBCCCuh6ItCLk3bDNNLNMlMpDDlIt0Uvxg35Fe1gqyzA7zezx7pmXlqE
07k2Op7cEFGbUFKzyqlEMuSNvezLUI5ORkVszOXx4w07lsoJj5z8PDihDh73Ii92
mGAbKFFyXglLAr90THA3PALMT//z6vVaAkJKCrV1YrErp+P3Hp79GcUPuRS4Fq+H
RRMv3bzK7HNHIfZsioV4OcBCGHwW6oqqktpBs+DUhI9M7cem6gwB8xelcmm1oFTb
fkXnvkqavmMs/IycFnbbCRdqeHKjCQDoC1YMFOr58pMTfa0QLOKTJP0zHI1uFHXH
ge9/IS4IFscYy8VX30Vom60Wzr4V9L5q1wvir1yB/jT8PIQCB3HQ9sIHhlzKMusP
oQZlItIejNff+kVKoHFXGkZFmCL9wgMKQpERS7MchUrwkSg8aersJvUnzaRHzfrC
GvKCdhXCL7mEVI/t47LQi0ajv5LlHCvMkkjnZjQR3QvrTHFSEZXfnZZmPsmV9BFn
wyP2QMriydVtTtGq+QUxcKtSjsWcbS35qf/hRKALBd3XFVKzhpZcYmB/LyOvyUP1
pmFJ/U0BoxY7bLMD5nwkyAlPyqsYofo0aHuQLRbj1HPebyjeGZMgfwl4MwnjyF6k
p1BGNUjmHXUotIFw9j3mEYZveNd1PSE3Wg53Yo7+ipG3KzG+9sKLSsxD3Of02iPn
qbo6/w1Q8pI4zlctaKqnL7P36M2Ze7iIyTP0+7L/jMAXPprKao8PwDjtBMucIoOd
b9BqdnbrJ3S9/Y7yPoRPamCG4PyMD0R8S6KWGxSuVKr+VIZCsVZ4g5yf3NouHyVg
etOEazW11iprw7JfTPr8gn7kJjXp34TC7WLjbiLWiNrrLkE0b1SM3zKcCjIeBFNx
kAbycMf71PErH3y2sISGb8Jba8GD2G2ru7VKBnWoOpKDBRQWt1RkT/9OmfGiJD0/
FNFMSgb7w1KWNOnZi5PnAaB2S9WGU+z55/YMinLGDarIifg6sWxiq4AEkrUfn/pA
6ER6YJIXjzuU1XIaDh3KWEQPOpjd3kRHbcM68X5RdiTDFH1rJzZLbe8MXKd4GHZd
5viPRpTOL96blXtdef08vuqhd7yY5PVVkjIE5CkSFwy4vUIJZ8y2wkiRcQt2G/Lv
PNRXVpO58N3IzmLtxQSyamNVJx1b/bO2wxaefagwgwi72SCkqkZ4c5IuEwAR0F7o
2Y74UlOkrpRSXez9fezDDsaCpZTQpaf1H+pUJTFaNrNaW/QWZYc6bpcdXuIiFl4N
blZLM41AC+o9ZlRvDXcZjMh4UIwTmKkEDSF3bULTobqEQfVtniMwMKbp0g8k1vdW
LaAbsqRwr8nxqMtuqAShT3FSwqtN4+cG6SSazXrocSOWe5UpgT+OLVikNdU0fkpk
XOZwk7xxnnppvtsw9gCRBH5FOp78xnyc+bpwaoh1lMmfY1vvRHTJeorseP2ycaYY
00oZtTr/LWf1FN4V63ZFFWRuyK0elCqRPGi7h21kX3uelRauCxasaz/RKaYZImca
n4QwFAwUf8EWGkK4/HCteMNyBfh05/z6I+dUUdWeKSQ9CXNf1dxosqjTdN3/EZt+
Yc1rE1kQYl6XSyf3caSzYf0Ua8DAkjzBmcGNTXyqWpNxyCh1ty1A22ASU6jhs8fy
bP59p/9IBD6WtN115hcgOBKWUjqHrG7P3+QuCht+08YatZPH1y3/04QgRbp8xQMH
w/cIY5ZzDMNJJNu9ByA9WFeSiA0YZNDEclUfgMfqb0IP4/+EdcJaUgA2N/vyt9k+
9xNEaHLfupUbLMyzH8fefbF1J1MZsYxOscjkX7wPcv+68B81EAfJ2hRYZfwbFvf4
LtqmXgMlUPwQ5IoGCU5cGoWxpfiycRZ4F937gVLOo4eW4Sn+07L3LFOCBpF13kC7
JhKrt5annlgTMjz16DrTW3jUb3SwOf5bxUZ5+6AZh9TTtDitur+pX9SYBVEI8apD
LnHsrajYB9kiyTz4L0/0OMU61cjU/iGd78WAn/n3TmYWOSPUmamHoLrIdW+zMSZQ
ixgYSqqk1UINH3uB4mXRLkXI5OaLrwYJts10OmioTW6P9kPjHf6CfRImn0jFvLzL
+ktbFfe9Tt1cRLrTzkKLgGPq87FtiJIs3DmOprFsjH7HurPjq1brL+CSJV70qsHB
EbRCrJrL8ON+lB6nFCY4pqZC4eeXjFMtvzGJgcnN7injmd1IaN7iSaU+Qt/JU7eh
6ogvHRT8FIuuyus37LBYwupMG2rOIe1UH5stGzaKhr7Ud1XFNEE8sX3DJ//DpDsw
sj+6Y4yyJUSClmmW28fWRU7YCMoSDoeLz5BokiK6juN/pR+qYd87Ps/H+loVZIDX
uVSAilgmb8Qc1QdiWI8B3M1r7DoiZsjonRLD8TKxfTi3VYYu3zmSVaCzFJC099DC
vIiGEqz4QDxW0Jqx28s6DT+LqkSeqznnXtoEZDAI4Zjw1FCT5j6VlZoxmFkS0S2L
Zud92/3b1vIUjhvqcp6xtbsuXCNyOYuwEvJYMAZ5X09PNdnemmDLZ7LQ0VQim5nD
Ngpl4PJjxlGgTG5+3FS7r5xjQhBGqqe2dFLFzY1gwK/2SMAU8/CfSPTlbo0Pt0SN
X9Lf3eFOWa3xkoour/PLQKzYjUc9kNnZWGova/3YHKMgSu9oO3hlodelFShSTDHn
Zh1buM5pu1tju/qIlrpt10KoUqZHonmNSx8lURlnRaoy/3yD8tA8zmNIN37HwW0j
d1bc7RGEH2bqkUouMUhXZvFOWRXkpfPeEbbX4sdBssWqmteDnkf1fO3n/5u+qOSm
kqZMDyNtxBVPNxcaLzmarNnx45R2AoGJ1P2YkvTYNXb93UB1/1eCcOHE0SwnF5Ds
iNemwr7RvkaLAgtdw2jZAXYGMmTdtYkHeW68P2D/3G4/UQAR6SNorM9es5v0QDdY
sPj7EIu8YZcdE3bhyi2Zb0h3uFx39fR+UAvZbVxj95NUnRsh49++p3eXogUYkdma
M2idLbCR8juVm9C/HARPDmJXriRizRKhFMRev9nyeALL49OBkm9Np55YmCkUNKHq
FPMB3XGXIrOwbp7j4bRs2Dpv16SXtV+Ft09pWmd5lox8OK1jtNJ/cXtGxqvXCkv4
8fEwaU8WWnDV2Xc9s38I04pMcFK27fwu+i8oqdnieA7Ftcva/EebE1pohomFbhCu
8d07FdA74Tt4+R0qzIz/+04hwN+wqlhgAqWJYbT3u2cl+ko5p2XUoWq7YsBhz/8S
syltBMox3NnGHWozY7DeW8Uf3nvCxHtYqh4izVVr5jzRdGJx5kF2rjA5q8RuhVfd
6PnW133uSzEei9jre+Gzt9L+Ozz5xYPTI59RUOkpe/111pX1neL8BjD1N+kol5gR
aTYKeHwtUrF4u8kDk1JHL6umDBGELToi4tQ6xq1r32PK+zia03r2/u4xixIOhcTW
YojNKt+xlrr3bH7PpT96eZ6dmXyc7VAwUqufHjV1X9U1hKqw5FqPs7prbTrYUZDx
urtVIkxbq4m2OafQxraju7XV0NEN2qDT1zaJ4Elypwbc9FIRKP0ybsqfEpSPV3Li
rr/XFp75+f6zsjVBNtVxYUr+/rCkKjSeyup7fvBkh7PMte4j19qHW9uoozCZEBm1
FBm39nHrbreZ536voudB+AO+u7sGVIeO63GwOzr0Awv6z0dIMHubX6iu4Og1rzKS
U9rzE2NjQz9uh2PsjtvsPSMul6ecf2557PbIWcIPurQxnHJcyWuZB8xL7sy9UiEI
mLPaARqKyvBonZwB7v9/Ryq0EJU/TojzxRxPW9K5I3/r1Lisck6T01GbqgYzK/Xc
3R8TKF/Ttbu9dnsV42+T8DIlbcXRtEX3gBOt3JtQ7js9UH4q3GJBsqhp3Y2Qi2y+
1TTtwBQxUtRVoPsDNOaOQhRsMktA6tzxtrcIBmD4KMh19kmEO9twSNN6ziV1nUvN
K9iYxxc7KYbj8frhxLQsxcsyCn+qfyu+6w7tS5KYMZHdn47U0yhbFKS9vMao5RSo
NZDKnH5DZmWY7aDQrvQY5auMmNZNCoLWplo1vRWKvZNvUdD1SF6tmvTwNMP4IE96
6CjvjHB2opzw0M83a0m1PgwvdgSDw9MHXoJK5drHadhMzT2N2e3weItv8yWupVTi
oAUVogtP2F2sjD2wn447XN+sU542iF6Nq+W+NYgPv4I/nBQsWI60BFYdgGNqz22G
30y17SCCEwsE9mZ0QfVjZx2BudUpFHebQUnRQWZxMdNt1nI9xYWQd7hhXHKQbrd9
ubXeQnMGrWpq98EW9pVLayP3bJmJWAsbBSNgQsnGeufkyCH9StMYKaotkb8Gzmrh
AYB+eAIRydd64GI4rJ+ONKx0K7qmo6csgWo3CjnsokrSy1Zk9ykGeVNjlFtxLDAl
RcS+aRP8Uo3iXp6pVLdFviSd0JSdcQUOgPMXYxQ/ms+vMcO1ZDnmJoEftGBdegWi
q12KKnbA4VZ1ndjunFBEYA+QMz0YmIEJ5EHL7lyMBHQB+mwNYDIqsnMtMADVbYx+
zd2toLCTHWWy5Q/zs8YK4ala573nA1yvB2OXttmqzbqlby0XDX1JUMsQuNOEsPx6
kGyR0I33JIABb1xkgZPjvanzM16r9P8/PYfwfV6iVifrKKWGkNkEIUNouHTStM8E
a+E4FcQWid69XIEVMz5mm+Es3+OSJwBAKca5seI8P52MUZeHRRnH2RJZhbuxwsi0
KWsLHB1AWwOUOLFLPKM8caIdgBOuoUmPh8PLSM1UpWJnx31xkWcHAEv/QUDChSR4
QFhaLynvjVfKzAncOZzsr4WsByE0GWFdfqSsc+Hs6DA5PemmUpScTMtwPa9PQflF
2Ofg/7Ot0iTHwJikgzpDVBtSqZOKONc2QVnCiOrab3/cq6pKwHH59vTdKH7aDytK
OaEyfur9A8n9WZZ0pm/wAbS2ePXLgL28Dcu6JeXQVBebmfdlUfY2XN5rX5F+2GTa
PsvGZEuE+FPxT29KaZaIIGPhBBefwGKwb492UZBNu3+8xT/bckKTu40osHOhTy4z
Wu9Z8z45UYeApF5gE9jak9NWXAeyCebrLWHnQHKKl9hUwfAgXSVOizVA3UNih9iY
mFFbx7Da0Y2n2ufpkgpdpS4xduglVUQvfUryRqi/gZu8n5DC+7MDD7kPxSM1nKY5
9ju0Ef6JwQMCzBku2zbhbB0hRwRpHEfTJ7sPNsWIp7Pmjt410smx/oiOJ3c+UhFp
7bzu5dRagtVwy7b/BlVZSJvk8AV6ILt2M+DocfK52g7rOC8O3aJVMeq8eF5e0IaC
2tIXCv5vsaYEzrQT7b+KkX8IlSBEyuiH/x+Wh4dn82hxa/SIu0MBwxlaNfF8D69P
oi1IYATmU5E5pcRlhCezTXIWFxS6XrCJsyRj0paQXtWAQPI6ttWw9VBkTm06lzfn
1kuvDSqqQpw8pnFwRcQR+aWDP6o4+Sp7Mpycm5spVoWW0Ad1Rks+06G2463P+eNm
becTWsNEpT8ZBCexoCBBuKlhJn35ijDjs5E42fit+mhBPRXqBmo1t7O1qHsG3MiB
M6pmSp2+52+8toN1ijK5U6fKeodwHnTIdR+mbwGQJQiceEcNwOPCPoqYykyHAEyZ
nMTPccDBuMME8+NdLHKULC5P8tBBiNQXPKt8GJPogh3dqOa67IE90/fKB/QeiuCa
CW+Caf2yB4IZfKFG3YQw6wqYLNyG3Wyl7yZ8tNNh070fEwKmTUA9+VYTTt7iWxZa
TbS9R2uNJuVljqC7z0VF3+o3K1Ywc4Mg2QK5cA68lSazKGLLN24rdm9Q4PAJJNqm
iLTC6EAAPmZ/dfB2jjXTNMn0H+v+4O4LqH1/8I3WaJOqNjaDY8B1gnlmYQxJaC/I
bEQjIyeKfuITd3zUy2IiSz3B0IPMMNukTlf/VpZWF2WxN+tGbA2SyTkzymM6oLSM
S3TQduWBg2Srd9Am8yK3mnmpJcJvhsYuYJT/KJVME/Z52S4ddBd24lvuENGG/ZHI
hCbUmhDGI+aZqgTtnRrUgpndMQA68a+Aq23MHgP0HI4dKam/u9jZY+1tDSFJxCEV
nZs7XbNQ+tI3kWafPBsn/lT7E3VR1xnNVm3YPXNqnpVgw1O0wAjZ2yfRkxn+iS7S
fEX3Hu6U7czLTcX1n88EDdfHYyK9gd2Xto2iBlnbJpNrW9C0728rgPJx3eZ3hhD/
WacZCHgYlCylygdXuPM09I9f80WFxoRsWjCFsTexgHyTaZw+LadmMr2ob8VlgUnP
K2wMrBih486XyNLhxk71VH5UyCYzPd6pTKM7n18ngvHY1VZtOY82eIJXgt8pLaK9
4ATTlhGGE+eHajRBD9CMEidR/jvrIQqNqcnl1BLUg5Ei1tUKWD/mTZoZi79tRMVM
Uq0VoKFo/yoVKF9GCy/ZykkYNv2anEJ9Y3HOj2MXB/fKs4tffBm9vTsprjLzuW3r
IgJZvhkltPYduqk4YArednb0EFaVLRgDdSjgJEHh7BixUOyVwkhMtrUObDMOKWVO
pu2eEOLESg3ng/Bmer+nDLch+epo4i7MnqYqbHiFNVR9fcBGtsR/FgFu0hcgV2oE
q6js29BdENb+JC+z5p/yS93PSZSQVhVqMjhMlQztuH6jVaNtDCDQ3QfqqFmm89d4
lEq5ushyMP9ukm8tT2+wseeSkFvRt47Seg9iFsov0On04d2P7c5yO24a4e6qhtE1
0Z2Ap9JMfsvkvyJQ89gh/n/CbgQco6D7E0oD0HZIMdVp/EUHxfiAfsYVXvsIpy9m
HLEZjLg63hXbDNYnJm8Y4iNFPASmMpvnyTbxL5MHaVZX4wdLZs/s6lIpb+QjiEES
HpuPqcpu3HntZoPOaFWALCNqgZdSJR0ndEerJLQIhcQ7W9d+O0yansxyHztl1fIC
vFeV6geRXvWWFgCUQm7JCnLFI5p48JF0F2YcSafHHGgmhhGEsEVvubd2LecDMwll
dlo32fY3UJ/rgg5Sx63B8Y2sS3ar2V4ndp95M4xMkbgVqM/OhktQui3nJGYDcTAA
uCwjnyvTV2ZIOXV/Zje50UyGO2LdIZzIPelVNLRlkGlca6eaJeQ2sjM13g15jeFc
QmibEFAKpp5GzaR3X3liG/LNwG1jOZ88EketKauFbNhCcdNG8mEsic5kPtILOoTE
UHREiauIm3FdeIx9azPRHUBZmz8fyRuiNKKMM5lYoHTqQcHJtn/XgPC5x9V1tHFJ
3Gbsrx/RlyXl8wiPJTV4uyFWjNRQGpLwxWOK8fI0wgUJi9Rnea17UxteuYX0F9Es
TpdSdKbTlKj/+CYiCTQMlg1b6UHyL7Z0i6b2UTJUttvwDx4HxFGojbIkoJZW86sE
eU3KEc84O4uw5rNgfmbfF1s2+1o0JlZwK93OUa9Q2CNp+uxGcx6wBNVihlq5DvQF
6CRX1WFCP+Lzr8UY15WnCgh4pVz6bft2/LuaTWmS2e8TQ8xXVx1jNK74zROSdCpp
ZnFjie0Jjao7liuM5NFM1HpEb9qD8K2KCy34eCAD3w2cfgrTQAFlN8E45NyXnVKk
6o/l2R5fELJBANvgPHBOJqPVmK7z93CAjAlNpPdkQ4qqwXe+OpucmB9qUDQzaPH0
KmNKBBrv+bLxTNJbCC9HX+YWDmfNrhcDqDnNdslpRxN8Lc74EV0iivzg8LJWflcV
nuUphR5zUTZBuENvn16U/rIRLoTWxphCE3clx8ARySZZnNUW98FhByONk/qZcV6s
P6S4hAl3SRsac3kAeH7pLGHUtyTBG23/ak/zsibQFb7Tsg/B46CJ5Qy+BA9afvQ4
NYdtEgvz8jRWqZM9KUF3IPZAwWedUWkmZghksqbr2Dkfxcma1M9acyYFblq3WgRc
yyS75GT/ChWMAt8+2sWg2Jwyw5ke2AzyyRUk5+6DHv8ERQY+72H/lj5dJbtImiGJ
1fSXXk1D8luEwhOvmE2FFq2clgHvT81gsYQTTtDoyWtTk50PBXTAS7OQgjHwbhXc
BAD0zLNGn8C3KaU59uB91NNCpXBAD2/1wMxSaC0XZelM/kFu3Gkfj4udSCMXDIlw
b9HcSJ+4jeyxMaNTEqdLdhafOoR1G8eVSngzVs70I7lF7yPkPLTLcZCavGzkKMkY
kydH9szIKPyhbOsTP3vCLX9eEV0cEZjx9i8hODkduNTFp3YKQlIMUXPO/EedzDUs
M5yDAC3BsVYt6z0FCA7a+aX1UzRYQJtan3pQk9fFvAyPqs11dT0UUFzsyBncmX0q
9ucp9OCrfkPXbz46Y5Bv0W0Lbdc0pHpkIJ3jUMFVWE4UAV4N9YAHKo5NGts4E3PE
aaZIaWMd5bFEMv10C/Bf6NyLkDUqqY5Kskkul7rRzbyfKPyMaQ8N9vBrLXt19A2I
K5IWbgzDwVmrr34WmvtowAP1ciQpijjlzkQQwWWFAykEWFiq3DKH0xZw3gMdOSX0
BaY9ojmnPlqlAs2j+nQ6xbvEJu3Ru0DZ9uzw3u2/gzskD4JxuL6kFNgCLgbFMWtg
QSjMMq4ccNLIJKuS8AiGu6/03PImmbspinrnfj6pK65SVT3rXJFYog9FyEBWc6Wq
YipTONrX22nXiJlduHC+9bNd0kVYL0D7+uq2tUmy35RSmckE+fbmGJoaDrooCyem
My1JFKvRi2tPxOyxFCv41ezK1xB57hq4RKM7UQ7E2hhzNJZhB/yuj5/RumBMUTNO
t+yDQV6mLiEWnnzPd6kb8yjHhiP0e2MNx8V/T+J86IxIxtpalvFuMXWLraquA7Yp
Hp5OmRL525CXYXGDNGLVxJVHZwizq3kwbVeAx5+wubidQPYGzrylsXI+zF7s+DBx
nAr9r8Znulf20x89ZVaa+jRNV2bkMs5M35zGPF/3f/jFaKrZnX6NX/7lUX7j8gE6
6+DZdGUC7MCd7276B4xxlloxZlEgPlp79tNrEcQqFp098uuUa1NsXwqITQlFrS3+
zb53cOKI357wXq0GUu8RJW2WYaMecVd3FN5otyDuGy/AMexc7IVRXhQZecz9OA6g
DA5toTb/+LvMUSJz6OuuLZYiGBHdg9vekrkIQnwWsFcAFxrnzVbqPcKkWCoBNddA
Se/EI8thJvKdI86g1DlXE23g8p6J13UiaBm0/yGaTieoG1DRgxasunveI+7RtGe1
WA+QYkLgIWshbSui9f6VP7TyoOXk0Wsxel922U+pVOmLaqnJZnO6+OH6D+MnXEAY
vnkv8Tr/EzHJfB7yUM+n4C7CdnckYEAU1+fMmh2C098LYNwWQfedw+JNIiOPaFj4
HqnLPLG/OtP1d18dnQEF5MWlxKbRM+DDHIt99O2r+NUquMT4ZfUQ5UdujDBbeK/C
CFVEy3X6HU4/MUfsEo1ImnDPPtWYmUundL0BXJpLK5ueMHZBp00+9l6Pc+2qIqXx
IVHxMWVELDEN6rKx4eMEzkBKfzjQzjRd8R9YgUeE4VWJDZHyJIUiE3souho7vRZc
f7KuhoSWtUwzZGBkiZgkPWH981+I1/NgVaNpq2SPxCAiSLWSA3iCZVaex8iIN9Gr
3CZBSiCNjfBBAMEUPbP/PqXx6XOUuV9B8kdWdW9mzuchtpRJUCYLjf+/GnC8+kay
sgGueIy9x8TmnLA7v23TBbTr5XiquFAEzClN9PYeGRcwLihVQpbfPNt8I+tYFYbb
Y+ciZbPqLUDdM689tREj+eckaMA8cli24a4DVPLVHAsV1gefy8j+nbxN8TxsPNcl
6aQW+sWRnwWPCDlw+YsS0MBH3vQ6HXOZ+4EA1krtfCZdiyuaAYYio9do6G4hDFvv
nQUjSxblSPgVjvh+0TUQiHn+PVPlQjyuz4mXdz9vQxO5SkIL9PX+ZMABJnwY9KnW
QGWM5mx6iqBLLC6P3SP3kH9ioelKx5aQFr22DbR2E76uNxIHxTbKw8iwN/z0ti+p
BO1nr5Q9RynJW2uw5CCafGuoW7F9q67YSM8nVtyj9ShaEjURId7VFS8oxv2+RI0p
SNQ+CGj9iKzKO+Q87hFP2slRxMf/YxDT9kLzQoIiu7cJeYMbSWEssRbgA2e0sunw
BRNJpCv2nWx42P3a/RVCLsPJQ07gqL62Lzq3WtUTM7zxuH91yBBDR3m9neIxFK75
vI5Dznwnaaq9aKFzBNF7ip5Mvm72rpM1cmTP2SDsrRqHTTfbAt+N2MRtHqCSs83v
Po4JDzK6LJSvTgG7B+28N+tU8fr1jCJ2+x/hzC2su2D67TYlZYJLpozZuJRcfi2i
4K6akMfapdNbUnjrIcnca2JRZ+uchn7PXNuB3sE0Js7ohG1fMVIevE2ijeV8Oejy
Wit7a+SwwshIS5s6nMT1c74nw15piI2cjEA539h70tROtPamzzaUlfDBxe3wcSqX
Y0/5XmCjSaxyugtKx+I5RBXjsyv6eOqtLtWlY1AloHZuGzAHtd4GmugQvxPCO/bv
BLBDH74YT7SqUzgBZMZqAfOvMg3e16z57Ax4htLJJVisib7rroOyDn5gVso4Szog
HZVySZ/ShzMfvZUSFxNAtOkqoM3KfAKZ9MB3UG3PMbo6KDPF2MHa9F//2PW38VFr
CvsT42Df65D0KkDoP27nmrKfyliD1MUwulJFRJiaC9B58lge93FBiqvW9682nhBH
jjPAdwEH8XyhhbzN6F1HQS9cMEqCYR2dVLwer+CsBBgRvC/KgtDc0LQwCB6L72hT
f/wvOSgircFj6ebjwNN2daHFQbGjME35LEHQJwJ4MIb3bLMmkKMXNpSzjqExUZcw
66gZzQtzv4x7PBFafg/1ge4vaTQNGh2iNcJEPaYucKgR+KfB0p/snnnBfnUbjxCx
s5Kw88oo26Pyk+3cQlJkSIbqHaw7OKASfrQ3PDKICVg5vjQ1959uFdKzCYvder2O
uv1vBVaVV9Hdd8Dz2OpBSKgtLOXFEKO6AItSX8WdldC6b5ip22bh3JOjAbd2JotK
R9LYI6B22EHsOaoN8Dvif8AuBPARKPSKthcz9KmmLkRLs6BZ9bB0OjE2dGpzKt/o
h6bN8vppXoOwU61v5rdMPkD7PZ6altBvnuZ1YrIbb1v4pA6845NZGaTePJVdoVG9
NZm0EU9xRjycVZTebgcUkAAE8/Z0p1OfDlrSYol4Fl6I5XVJe0eD/h/wukiNA3ko
wbY7APKpwX25LYO+0CPH/++WgvmBQaPEINuN8gccGrr9UkvQ3SCB9tk5p6Wwgb4V
qQxzmuKe+P6q/ZV2xXH1SApLNA973FuXqOmpScTubapJe7zZ6RzyP8pTsHBu2+gI
4PiUe19dmCooy0XdJoLOXXZsXCX4UkH0dA54T7dC4w434twwoMSDdbb43vggSkQe
CmQEUcsZRvrDBYNPv8VFyQCkKJPM6iLpb7CpQZXPziuVy7L4j2Hnif8BfPGDqrxs
gc+/Hu0d6hadn0gA0v2R6xnz/PD1rnLoqUysHT3x78OW8Pwav5qH2K1AzsjExnWl
PCBv+ha1gdBTG005MOMin1HIAZy8V6v3LumsfTKIWV0yqk/yBOVdeYl21GwKNYIL
AjAIvUSIy3BDSuTd/ZC7QkXU/jXk8LaRuFOH3Y1eOCvlspnWZ6aedgyH8xqwkDz6
Y0VNEADUqvvNyoKFCGIGDpKH6a/7F/nwnENliExiR0/bSqUqPq8qagwlH4Z6tPBv
bPFL/+2auOhuhI9dyK5Xgi1kAc2pZZ6EtRSxKAiKwKS7DS2TnEHHsA0sJPeJYCaH
jL2O19pTuUbIozjv4pPo0RYEkvkIfTIwse57/K2e/6GnNZ6nt5rldVLHaPFru3Pr
oCZz9Zq8pSI//UH2d1KT5nhgRVcqTY5FGZHHfMcitLB7sAvmGe4A71UAKiH58oI5
AqEIEdU7O3hyaIKreeQEJCPzY8CVSQ2L16yJjsdE5giMFjweMhY+I7ueLjgXD35h
f6oIc3FbA+PIQDSoOyQCbyT46wV/QRJrHQ4txneLY0xj3V0adApbUlstAoDcsYxI
wYGZdRMYNibeupcTUtFGbck0c/nO8tiUmFX9RCcEUQjyY6JBmPTY1JkB2VshSNwc
g+UAF167wwRpLnTahfa43dyM8QqxgfF2iawnjHNx2u3jV9ykJxtD7H2vY57dru51
+RPT6NU4u72lSZMoQJ5Vo8jR5UxXRU0bcOwwbo2fWQL6rJBfduToNkECnKUuico6
JvgRQT9yyRHI5HjsB2eHQPnug2jk1U6Mbp15nLt4R9Zk+oTdqD3mC/XlTgxyXjrk
faQpTf7gZ9bxQpPpGJhKTEZZ/NB2ktsp1brkARLFkZldvCfU0lqtruRMJj5tDjin
nt3GRnL6td/qNRuit9WUVK4mM/KmIVEbo2h3hnqaPzLrTvZGLtmxwq7jUvnlVE7k
/Fgn2niC8kVA/0rkDNzPqjQRbvSR8JaOHtA3Qp1AsIyic6pjKL3ZfZqpT7vITxSE
3RfzKReIjE2TRb/2M7t3IVZVBcS8yp1p8UP4V0ZFy5HGkv0aUqDiaV+2Gxe82LpS
qMtJ2b//akdHt+4pqIMmlPYFkN8AhEuIsVBLLz8A5kVFuJl+6E8LcxVrZX0ZxQ5I
Gr4A+jJ9Yy8OPaumwYGsVA0cnJnFBSTzuO0+d8nW92w7VYmE7xHiSGPbcdx6LiEa
MaIJVmf6NBi2eTWz0MgvXUPfY2+qGSbKdaJsdx/6mGkGswqWGXQZmN0oWTO1hvJh
Z3Vot3QeAotIIVRhG2cZySd0B2SUeAGDBPjLFtuYywn+Kpa1lsmhemSANet0OpVf
ucfqmha/m13gMBgV6crXVNVUEw1nSLs2b2hJXyDvNTBkrU84nRWu0uWAYTQO4nPS
F3+tZqkRtl0R4NG8ADknGw5A7mDVknpbpZitcd+ZirDpn0cseUCcJ57gpKvo+I+l
ghce6MqTs4oLqG6lPe3z5ZTxzoVVMdb9G7zedZ6qXU6MUEnDsulPOTyZrO8O9+X5
UYHIJ5ya3doLAQMSKsEYoU1jF5YMe2coIEJKxJRNiFfAZsgenpUsTyTK3Z2YnXP8
h8Aeu5qnFXwdlWDd8IkQvrb9oYBnZNQao3a3CmNGBqL8GlULVvA79spoKqvVbdX8
vK4yz8WmO65DFQ9+s14PTeFZB2DWVdZJ5C4QYUectiZ+Q3qDaotNxV0YyF5+qMUd
ELuiHzQmTMfKKPorXIA79NSA5dIltVcJpi0y/op8zkULm4b+C1zTZs7KvxWvBS6P
tJm8IUQDgJayRyd2+6zspZRzK9cqtdBp5UHP6N7fCSAHDh9tZMAV+A5grPWOExAE
uue/vBsE1jU/rFNrz33eTTojKz2mUpFOKEUWt9NFcPwvCW917ZhkpceP4QFfiBQp
UB7Y9dVOxTENOHE1hf4yFfa+sJ9vp9aJnNi1XaAjh+uQrVtMCTxtwm1GiSGZLF6j
JTNxix5Z55UGkeIdcgnqT+XJKV4HC8jOrXnxIa6RvpZ9LvIXUnLtyToUK6Ze572J
1mC7xl7HIfcXyRVf5J6RJv6i7oo4R01lPtUO+RAk1D7hlO/Tg98Gy8SNGa/HpNJR
POIhg+7uy+WdtOinS1AEQzyvG50X6pGpdrpENz1d3eWnl/E6k+Rm0QQhGvXHLCos
Fj9Y+ybEloSL2eBlRAwGIQlT/Q+EOn+fvQb2u4bVY1UdTwRjse3qaA8E/llsKkF/
PlP2nRwFTSWBSeJb4XcdewyTUyynKBw/4yI0yXN4iBO/M4pv7V3sLFZrqrFqFpX4
/TbtB/tyJtjRRclF8A9mu4TA9VQlP30A9AiFD2SubX0LbbyOI7Rzlj8YPADvs7ZC
LlKxHl9ZMyJyiIhH2RTD3wKKhMb3D5PVWm+97ZaV5g+PxPAKNGNOfQFox466MOKe
P2TQ8aujHThHT0iaPmDhSYNJIuzt46Fw9kx8xL3g05RYXkt/HYN8n6eYjs4gzPXu
g0dgMdQ5q969igkiwnLgUdVeMmkyx67x4yi0duhgHgRh+l5JXQlbkaSxlfu4K3FT
iWTw0ukiJwSd8DBIEEs1DM7TFA2XDXuhk3AQZDdeNzynYR3O9RP+93cPoF8vKg98
pwR0UfpKR1WYepeTysQQXHfQFAfTMl58zCXfaLPhykKvTjQ/TK7Vo/fL8x794EjE
ewBD0FG7GzL/OB3aACEUVVjyriJQQGBv2D88JpkpAJnjM7mjR0YMFqviVJO8lE1D
wetw9stKsVOKmanYweDwWBJCLQJDCSloLbOq+LXkWHgDwn+XERUXX5Nn+9HMe9do
+ltVdmD+EiB/gkqvyAsU2E1uGcx6JxOhOMCbIkHIZDGm+HaBEmn65WJ1x5XQ+e4Z
8YGlRtww15NbLJZz+wCkF67KqLeLLsfEwbcC+Zp+idAKEWfEcHs59+laXANJc9kU
aqfv78mFnaxIj13OLcalkqbiHc5oEiJI7vnftFAKAwz89HrmsZum84SKFOJNZ/40
Uj1sFFcajON4AjciW+yV7MNXRRuwSh2DyQ5pVlHM0NKAUkGGvX1XAkH/XhwPB0KA
rBvqm54lPygDxJg/C7N7jOcI4gCQFent9HqaMNnLsBhAJWVx54JQyqF4gVimF8Bi
GpEOjx1o/Lu+J3KfYRI1TRs+lxp/GVBKoHdvakEqFSdgIUmnpGwpZIizhPnYfpcV
9t05uF+J5yZ13Z2T3SjPTBJaL37mCe5wznvfq3g0LsvDutkAbkwXXjozC1vZLHUo
SXBbFG310Pq7YS0u+fEikWWe4aEKWK1mGcGugLPtfVfhShJDGNf/uAEabU4eci/O
nS0Lrwf1A7NDE4ed8apOtgZY+AdJDWkd19tNm5AXr73I5UH4/MrxLa1EBGY/ZxOK
FvnYRerQgWgXXdYl6zYlirsiiFLCRJtYD1fH8S4aZz97+RoQ6H/mVPYxKYjC/N1n
WE+TiT3pUP0Zg3M13JTfajujFG3r3PTXYUyt1ZGbJm1W/ViK6it0VbuRq4oAlbO2
pYjuTu21jsoIVftcWaceJheZjdaXiqkU9KuIr3xl2w22N6COFZLhUc0OHb/uaRZu
Iq/SvPw0FF0e4rgPIQf1eth0gv/K9vZFY9WYboi0js9CS+4YeeDTinYSSt9RwfsM
Rds/b5oqNkESgLRNQewyAN/QpnainlLRFfKQrxkpD0H28ulJjHHmYzppCsQaOogR
9diT/kUEXGb2QaLASoAPtnSZWvMy2RU/1njZnP7B4dOGYsdIJnEj46adFgtJEaWO
9mNAb52IFA9XrT9/I3JhApZAcOyuzoQgOXZ1dWO0fffct0ZL7ZkcSVka1AH92pY+
WAhMEp3952e0hfu/nULTVRP5AcBZRClqvaMdHgI8hxfpNRuMQhWQ4gfd7WP7dDCZ
WNzIaGsrpnR+Ul2XYmp0GMAJyMa3G/qFzPidMuslee7zr1Vs5V/5QA2o9Gq/NlGX
LcbqhUABhMo7RyQsvmp5sr9eaDdlyp+fdYjU3KXTzDIGbYIL/TwDS7s0EqYZR2dU
1hEOLNBrE9+GUyRS7KSwhFVWQ6XM1E0vFhbO4d0kvKcjYc4K1FQUvy76Vtk2HB4T
h+bDR/7XapYHgFiBIFS9altAsxF+u1jJQNqmItf7t5upu+lDDDWwLxhCGiV15C8o
LPnTGuqc88NI0F5W+TbcNSc8VT1ljIjfz5QVTOMiJBV05g/q/2j12nrPAQ/1QIiE
pjTwP5LXZ8xQSREOYJoFRoTs6I2MvC2zCmb0lmIET6rHanFQxzfk5UJEi5HEJ7Q/
8Ro+zVYDch6h46Vuf0rYTIsgccMNt+0ZVBTygolPJA2xxqAHHt7as0o+0BfoRL1k
RMi6hnjBNmCliqjwS04u0jQQ+4jT2Is6XnKla+Chgdc9Y01xv2eNVUcTFDdbKxG8
+vK4GE09zScsCzrsMbVeEPDaKa53Crqjy7YTDHGvRh4gU7YDxFgFO1JLzN9vxqsi
PUWtlCgc5y/CIDta8oZKUf+YZHf3u7yACAXOfr/aaXHAGHyGqZ2VmU6ZOWUhBlLU
14qsGG7A/Pid70JWb9C+kvRJ9ISobj946bBteNZMJpYHzb5647GaSh1VSOjqa5cs
os0QsyeFW22XFDzhNlUZdouDOfrxQwMs5E9ovCyDOsvZj94/0N6p5oU2Y4U6Efmw
YcD/pSFeCUXSlSxaihPxK19FkWM1qIpOjXf3m1gSCFJ2qnYMGJf/NH2p59ef11/X
ZF3l141PKAtMDRZXu4TfBAm+fpit42iGzFCM2qpr035CABwpzKYnO7/zsTPAsPPK
XkxfnhkRGTkS95gbBKJ3fcsy3zyDctFFziiis+FVEO8SC84ze4mZf+++XzarHqSJ
7TtfhrmE6neSq4YeAzChukQN9uDRNb4QnzdXFJSKRvar9ncWD4mmGqA+/Xl+XbMy
rRwVBQU/4T9LtNIB4aRzn6ub088hXyqUex0NMq2Ze6TB2n96aSkb/eTu7oOy5lDz
6yrMdgarkp+ObuYB66Vh1aV33sAFtFmbCAhKqVNtg/0+65RGUJqu5nlGau+E9tWx
pDtFRSQDfmVOsbi6Vly0IUzI/51B8i2gL9tZuTPTGBm363VFeS5ZcNE8BgcguubS
2jAvBUem7QB1LkabO6IiiCvs/FSIb8d6n01ykcBIq2gyUpQACOQaj3Tss+wFx9iH
5pdq7r5V5fvu2pqjVP84wQ+DjGcEklKDgbB2Gqbt/lrf5h3xW+4AoujEblelZP+D
GNhEiWbzqRxeC+ZV4dSaaHlnUucN/4XOiQtIj+Bt94ugxLVifvr2mT9tQ7r1Net6
Aj8iTAEZ/mwyolaP9kMJPMx7oj1kstvPFqokjHLuGKmbdikerVkONXgwStaR1cGr
DYcqzWNrBibKnOy7SNS+XEHrgKgAssQeYmD9jW0/frzrxtsC9B2/MI4gRzDaBMxF
YZYYZ4sC9V5EHJ/wf8jesAjC1Vw1K633CDktVkAADcTWVrJ3ndveUJ2/AsBnejYM
zbRpOdmuXCpRd19MoTtzwTLg9NSfvhH+wGAU36m+C2oC/vsGbQ/RpdBjhU5S90lF
TKFGIbIdBQ/lEmy1SMIM0gVAc54XQbax2AJxgHo2ClkBy2TdtoHoQ/L507mecoyI
OanczY4dNwhl2H6hkdpLZ58pOFNdDjMXZ5ONxY+dp2o1cd/z76XQoqpFst7RAdAM
q10Uen4Rfrt0mrktUJbcMiTM/h88tYtWKtzXbmaFsxVn5uPj6dXRcfWnRfV8Sp1W
tf1U+uHRA2PYVv+womTjMPyAUHKyocGCmNbvL/4GDlB5/jirD67Wb8r4PPNozyvG
FhLAFt9FFbkaJBiFUhUrxYfJogEmL1RCX0IWVetB2Dulz+4bCfQWb/dIM0KrihEP
BPBibkOS0AiXcY5PKO0Zn9iUpGQFGPy0nlyeBWjUc+CFhWhDcXFJHsdrnWoTZ6F0
iR5+DgDZWnflvQeW/tv8dbh7nG4czZmettNHW2xTzqHHuQh7crdfdKMlNgRKZTYi
hUOILtqvSsXF3RcHTFVEWFoh43SzMXfovFykv2th+yyCwotMNYbh255PaHEShJCb
G+WYTWkvWkkYbrujHzmSEHx4L78Kj6zHUAmfLR57cbGE0dj8/p7vqj560lFMlmkU
7YqWyrsVbmYGVqeul1h/sABSfV1S6NwkQNi85QjgxAgwpgrq8joSl2D8jM+Zr17G
EBlSW3Wjo6iAF/Gq5p4VUY64jdnGvzjgEfK4jmvo7jtwwDZ51ZKLWMONqVs7hqxK
Yg2qExxdmMyTWnUOsjnUwVT8x8n8SJbebVakJJXg9AjhCaiHFdgV0F8jPJ2HbnWm
8tJbd4mDd1AJf5mNiApbFmepVtBxEnV8tFdU5EFh+n2vp3Nrg9HRlzpyLxINOs8u
BvqFV/WLJcEBNtZHrbJGY8Yy9bdS6JpL9nkveNc1MOIIVmDvlzvNIlyy2xSvfq9o
OxKWbpnpTUuJ5p2tNVtYtxdWXikErJGL7Qe7nzeA3AOAqbOwVCoPVS5Y9uki+Sqw
EN7cK9pFI0T2OHNqP2ENkZyeTQhuFn7ixaQ0EqbHIqOG5zrE+9Z4eEfSjWAyZyw5
iQgeJrjFuO3a1AvNKELtYWl+2tv7ogWN7CPYLhLTUwYJSXCZSG0MKMpnIYmtxhuF
F34ulJM0ou0MTn7kZybKhc3UF76s2Z8r+OE0IQLwW5+dcnYbEzD+1kKgs+0CaOqK
32awK4lIkUFvSb8CbkZfzA0wfu5NBKFKsEFPsqXH9RK3nY5yAzfyDpRtfdcOQ/FS
ZcnPvR99Eoq1BsfwXsdB5UXYdD+zxgmMKnlP/qoStV7C8g7e3vqzKuL/HwTZJAJ7
srm2QVpXe6zGk4u9lQWFWqKb8DZ2pKKecKu1WGfJGQsKKatQPeZCd9MckpRGgDI6
CldBEAG4LDvu4oUQA5dOwQ686pr7sE3xyB1m044LaEFoM28KWGjEZLeZI34sKKPt
IdlUF5dQ4qCiiZRCjpDxmpBxPCvpgrS9hJzGT6J5QOIhVdJWPT9l9FPNHQE5jGul
5BTVQkGVVKq0PG8nEoDcu7YWHltoD0JabryuADiPJOdw2xDLwL8h8/rLYTzOM1LM
daqp4EcJb+rxD6VqXtCVEariS5LhwQOhMp6lzfmYU+5i9Oo80HZ9CMYAIKFMN/bJ
0UpUQjfNeCzgHu5j3LkEHmskrnFsq+64D65CjxC0zgP5uXBzeMXDCy9dxDeozqdS
5Pdfaf92jKJlNe545ftta/xw637lXFkzKytCsihJqh3yUYvg8Dfxc9EuQHabg/0c
s5p9FyiTTaZnUnt9dSPFujKAkm5bfiRImCGERDn/UOJ2aNvwYkES6GAGQQpO8P9f
MhQZXPkG/9oTtAzKHwAJTgdpf7LQFCAB2Q9wJr85Dn7r7PaiizcuizN29B/YsX44
0dt4utltYdzxdJ4GWW+G1caAmr2NMpZLiPerKNmH8DkWug100sVb7kX9a2AiLiPl
krWT3m26xe2zGoR/fzlX+MKkpB7SmH2mU1XajeHvKHvXrLMasIKwQ9EAxmdVobdS
P3idlTI6HVHoPZ53lhEsQKGxRaMdxiZFCsqno2Bhnv6wfZPvQd6vRbAXoE1y9WRK
ZgvHX4wOJbHVC7352whNJjVCih3vZStf40JYoJivAKkrGQqZfdWM6M7vsC5/5nYI
ikFss7w+ACr1ZKynsXgMUcm6TUBV5LfrNnrc9PPEcRicrQc5H9EAASVaubIQnAym
sUpgISLnGJnj4o0DrHChkg/1rBFgMvYxZ5Y19LhSTxXaBUB5/lR/SgdE85Agubpl
496NO7V5BVc7jTEBqDJaRokX10NKL1jnnzcB/jk5XaxIhTLexCjmPOWgYLBch4jB
TXuMHFl3LUUcDYR1nii+X2dh8DALFGVQdy8eo235TLoBLvftiAziDtlq3DCfp6sI
V3DSLOCHlgw7ID0T7tetlN0M2anb96MYBPmKdLIY3RtkaGsIIHM9v3Ywj9uM/a4R
RsLuSLpDB926EkgwNbdAoiClYU0CoSD369iSLLmk4OjC1YYjOEkEBlp/7hcKiLHM
FxhXWbnRHIR+3+0R66CNk0gAYdO6ow0lwyX0UsM+lXJxPJnaEbZEvd2YESYyHJy5
AglnNEtIF1PjjWUfq44jHAuW7hlcS63B87KWQcV41jCRxORLVpHvmU+ca2VbmwaH
JXQtoi/55s+WIfECMCJLZV5DI/TkNE4hsitC7jYpiw0u7L0O6sEv1JNcc6dvhX5n
c3EziGR+pBx4HkSf7MDSCl9SNd+oHhbhfVAX0vKO2FtFr2KcQ8MKoGs38agRf3DZ
Cq7VRcgT7BrifPyy3QQZZDDjVGrbAd9xpz3F7l511e1+taf4iLviFQ8igjJfbv3N
329PAoQl1RVQfCde7FcnYevU7uAmgEd/T/AKY7oK9xoyuxwTUqNyAYIYt2gs8xrQ
2kkM6TzF2bBNqESQMR6r8lnK6fmlIO0XvWQjy5TQ7nnVqq3DpWCEK9mnbTGGLCzL
WFzyTmvRBOallHDBySI/XwtKXsyWnGczbRaluUtz2yb3Mf/y+LKtAzxEnY+12Kl0
3fdCESrx45mDdIXA7bqFciAaYUDT2LpzGQlB7dvy9ew7VKxd2vtvsYvIR2r718yK
IWywmJcqweVnnUohO4EHS2eE+nhI2ke7IQlLihLwB+uQOpYQUd4QNPHGC8QfDcH+
GOGmaBWh0mUw0PHeeoTYfwJE9UYCcFLKBNR55O2MbJR7VI34jojZey70qE/Rsoro
cwuc7sXkn0FvHB7S8zGx+cbVWm6RuZ9V6/s19Z054QSYbM9i4BNJPcXpKTY6DB0p
ADM0Y3iY+rP3KZ62/WxMLG6RKyX74uVQYdLQ26dD0ZYB//iv5MjrmW40rLt20ra8
LQH52suoCgqxrqujPzPCGsF+GV9v1TGcNq+k2aC2BO+mrwf/Mq7gzcuZhmF8dil+
pxeMsUN7tOxIs9pAMf3L6/Q1lHgcQY6HpdztRnNy/pTAkHLCbzYSxmzcMSy44dLt
NHOL7/hAjzl0Jr6nnPm+2/SltaV9tQNV0moStmw/Jr+0+1HIRq8hQxrPEbORKiDQ
dZajoPMQFCwTRxpwTzvTbEMIP2fwVqySMAsWflcStoU6rcYPuWMVOG0zpnx0cJiQ
dAGfkNjTuTxzvlYfwq7a2Do5uTd5CT07BfpcLo7/Gk/PNO/33X+lLpDsas1wwa9Q
c4XxdQ/LV89dbRNVgx6XHD+xc5ITMxw+GezYOa8g+QiuJR62uLraulTcQDWKjacD
gbx8Ugxr5aBWm8eIsAwkRfEwd1jjsI217ddcbEFNopWnyjbu32ul5fU+0dJ4kstm
drZAAeyfb0nMwrx481YohkJb2IRmZAgUGYc/NulMKlukA9B8Aciqvcbj8tsZvotU
F03ZdhKwd8CV/bD8hljgWtfyFioHalNDs9XVIXMFAZDTHHfGN/FNE2bzSmrv/qTo
sCmadS+rM1g3etnr1mRyVTJvIQYDZC30Ri230/rMMLiMqrM1C4L1wfcRCpQhMbaq
WKZRwfehvWMVdCmcl/ymbEgeq/FQ8sqOE8Z0AakmM4yZq96PPcr1Io8h/PGutStV
uH6dxI3U4gSoXDExDwYEy4ljxcOB7t/82eN1qWUPO1rHNsYJVT+R6biGF6ufES8U
wmSWPDDWjTJd6F/qXAlTtEqKIGwmYRDein8coNWbeeNF9esais/jMmBqTGZ8q210
vxj9gmJfBmvjHXxjc6yqhmbvnZgKANSVHvLwFLEbmmmoRAy8K+RiWDlQNZOMvBKK
wTIMGa/p2/k2CXUgstCBb8d4uyJxmOybECNVBoBW7UT+WvAtiXzzplL3bs3v9qg4
fkMWa76Zq+0kM+eqF2rBLXpQlZm1cznLKMzEEhOr1MNFalUcNjBkONHuFmz2IaJg
6x420v/Boh1XMfOu2f4p+KH68zPtfQtOEdBJOLhTKpA/9A3yVe5vfma8yNioTRsj
0h+itN5CqyD1U1yGSyfllXbLrwQfu/dktd1LlCnc7ud9eYxmYMXd8y5lnCJWsk73
iIbVljCEav4tBEAEpyMf8QtihWEO0wF0gW+zByrKUEJqo4LHH/VHeKDn0DyxJ2Vu
ZAs8c1begOM83pN7UPdx3PurguhDE2h1/WitYnNWEJUFGMlY1xKuEcR90LaYdpQT
YKHSJ/GPETfu36Aw7PMSV3bSK6srrAs826fx+wHjuS3otb//DUpx8oAm5SemQOPZ
DGVtg7AAPD1kXtGA6MHWhR9eUydinl/TesSnhzKd9+urT2HH4JMRw9waWKQOOeqI
jbr5xU27qeL4zKt0E3SARIN04m6Jw9sGllmQYLUK+PpKaaOaLAdiRa+MrPtO1jRL
hdzJITy1vI0GIz4YuSd3OeQcERwoICEAxeufafUJ+9JBzx0isRQ8PMn/ffAprQ65
Gzn+z21bexs5P3888zmpBqsMRB/+5FCmtai2K0ZkzarERSkOvViotT/L1tDq0Ct6
hh5nVyvVv0P3mv97+5U9b9535kHL03IYrHZ83uJf5ZO8ucMmBbEnYJTkwCe6lw1X
qh0Rq+oRVrld8UbF3WMJVs4NhCp+smsOIRtJhSb1WG1+99+suHcykxYFZtbu10xR
JdFX0A5jfjLuvFxU63yG7enyJt2a2s3rktUr+1luSNVZ861lYgHWncD+u0OaHJi+
evouAw68VKO0yigPeoCUzOFjEJsmXn9vArnA+zjiQ7i0TfafVjBz28iX+bY9rUJj
soyLMU9iANtBcCjmbWask4jmYN3VkhBMyN26ZfFiGdOfBnB1tmfEhzjzXMD2dd0A
ar+yhpgxLMlGjiw5CzYPtVDleDyUj0bPm3RS0jInbioZKM+Ed9ZxONrixF5Levq8
WBVQUkWSH++8l0L4+nHrbnz+BHfSFAyKjfhiKu/LiASOWE/nJHHWpKLfcRW3cmQK
I0/8iFXdU+aNm/whioI32Fs0dLbQq9zCQQvInwV+MaBi2d8xu970YJIuGxddgIpP
MPRdKzmjUkNQYNdBdqQJwxAXDcZppG2fUNDHDims3BDtndP8aBgNYCezhxVns+1o
RPoO2MdnEhn4tg3m5bj8uggxIqTjCbuC11lmJfM1Nqt+UKqaFfiimvfzNbkXGZX4
Nr9eqsMWzcyTCg8jQ6RMdpHw+KJzZIFjYmYfldYpmX1UsebxM0MOSZWB37oPn7sF
Irj+C0pMgR4CoIPUpyXQ4tvTUzbkJQR/NJHyhT5zTG9SY37D4JpGznIybChfaMIi
hW9CtfqrQllOTyul1RuE1rp2YZFN/0md2azTTlFZmLEAzUaF0jpxkp7dYLSeITe4
cFHspzniMQDYZTRZx2fAM/YvRGqOKtjvDb8dIGY6ve3vQppVMYJndemljfbFSPut
+p29NLroEP5TRv/JLJSNmVqFXglXwRmzp7yMZ5p+XhuXh58GGExwkhuoLny1Ir3Y
MN72MW6diAOuDa6Rp2SHJjQp7SP0A94YQuUSepgL0xfgh1i9aD5yMiqk9LTVo2BG
lWHxV5wgpvS/+nbNhTUavnyBJEItezWshehK/IW6NCgGQN82/X17RHE1WeoeQjsv
p8Fm7d6zJ/il/8gtu5XJ0hdm6uCRXpcqNc8rzXFZit03FJhUBPnpMY/qm+v67VRm
iqPlf6lM4lNpPv+DvW/0F+y8A/4ZwT2q5Utx/CzpC3U0mYhDLZcWBTo7vInjJb15
Dfsy8xI6VIjvlfLj7oNS1lWxYrGRjPcbvPL6A6/yeK6BE4uCXgLWIfeNK6Hh5CDP
/HJYKxtZzpXpZYjOf8ICm8XqF2pVXVBfCFbhWeXOJvuFgKKIhbiNy36DoMg9kjV1
DBo//ihbr80Yt8TREw6trpRWRRINuV6cFlP/7fljJy/WkPHc6yoH7vLI2RugTjYj
AmyWTZyTGs6fxb7WVdZvPD7DdkPKXcwXxVlDFoEiOJ7/IrUG9MFUDGEpx7PtpS1J
WtCCUm3G0PmQwgvG3S14F8oUjAWjgKeaXI10FA9QvplvOJ1eluuAhXkiSsdDkaU6
CZOWhw3Obhq47v1qwUnDAfEWQXF+TKD9pCk6xXmcG+DpKyD1IBNgi9UTXydqpk3O
zpQHjROyMZjgcbpOOyt5zJfrWmY7ZdsdyWXQXXSWnYZHr7CoV/WqqaR6RG5UZt7Z
EYlAc25Fk6POkWFsPnEozkSOMQARdSDH+iwaENIT/oATEj9LZm2OAcVYDL66jnkH
Wa+BcS1pisUaTT8ls/Tmkhmbg2Ex0ulUla2TTJDqJ71cVPmJXtfO4oW0yQEPvAjd
6appAtD8S/bVjSx1cXh8G7N5/jM0nqsG8LdK7O631fti9UdUYDJph59wjVHIeHOj
Hv36G5f9leEbjAL9jUaZPwHVTloc6atis1EavgZ3R3SqpmPFPAd4kVPUWEZ8Z1Yp
ieDn3lZidw5K/s9R816jEUrPFq0Q2ty1A8V5wiNMpkHYyp9UIZXeYSn2Rw77FZdx
QFALn2q1AmkFQH7/RwOPvcCPsBGnYtDq0YCupDGj6l9EY3tRPSJkhjlZKCFOrXbk
aNWxsZbcYguWOKchIiOzB4uhDZvaK8P8WLS6GS8PFpbqd2jY+yym90+hzDiIAqj6
NWQ2DQjo49F9uxE1qjuNwI4rVdt7oTaPFjD80xK7waLfhGrja2vbxaiwU044gKcA
7ncOr3enSO0/jFzdeZsVoE9wwoXvSZlJsjAgvKaFRESkWd5X6oZhUBvMp+lru7Up
9f4L9aQo7pDsELPYYQll17nYjGhHSa36f8MfHNLCn+vPLJ2qJmNy3UtjFhzE0cHb
XeGTwvwwJeXssrfEpNUY2GLy40Bb4fzKBN0fqlugYAHaF/Tf5FK2nfm23tSh5KcT
zQDVdo2HteGb0z7W/JG/ALESqtOOEvLvRRAqVCZOrXOxEa66S2ejOrOdmWhUzMIb
2CE1xTpSUFIooLk7vSUT2Wcy3JOMdxaujnTFSBfusegsLiB2AfIYykFMXlKdL3dy
1H5YygEVKyd2IcwRBjjvwytjPmOsLR+Ak/PyR8Oa0DuHnIcVI0u3qaIpSB8w1FiO
OKOguLIqnaAcjXvVfPTncps2iBmpHtnuzvevKDECsmHvPAgvjTr2CuXSoloT4U5N
nznFhjgEycLY503GvqW1JTfTlyfJQ7MKDutY0LDcPJq2wveaQy/5zuJZtaKfvmkR
YzHi0L8RTfqmLGduXkSetxd4s6uIEv8lAlIPzYcmfWpu0DanxIYFNTnwevuNLQSy
CmZ/YP98gvNpD/jML6qt6Dr87O6YREY6jmHld5ruZJ/ay/sWz5iD9gr/BKylNaB8
f4hRjBZclBSnPS9dQvagqb0SKcPZU00qVAi6T3ncWj1TZE3JLVdkBB9apoTQhOGg
Q8gL7SunvufcgjU3aABb8XpderUfyQM0m4s6K/ShWhcCih6bEuighDhVlTYyEgYM
svs+WrfmRak0umB0svvoOV16YUCcHzRshFxkWzwyEDfm5UPgEG+PI/f5sF2GWGsr
B12pJuUUHBkrKIuOLAnD2d9Kh1WNjD4C+bWGtFUCvZ7MTACeKlG/U0Mi6/C75S6i
SOsQMWBpATnGvgDAtVg697W4kAbjp+Z3OsdCVgfqZAib3EzrKSxmGW0pBA3v0H61
rVSQtGjGENr5DBMDj8ZarWBBjK4YXak0bS4/oQFWkd18TEJPQxSlnFFdhlaDgZO7
NcwMCVsLLIrDDd/50dkhQYbyv39uPzFRO63rV98QBrkhSjM9JUy7wHa0wUoa2mYy
4yWhCrbMcTsHRmei/0llOtlD3TnfOlp8Qsn3l6/GiRFHMEkb7uOHmMN+hyAZgUtm
IugbdHDmhdDQpVrn7vtrAoKUr1v6VHcOv0p4jwUJGjnAlTdl3hnbomwPEpxcLZio
/Z20XRi5uY8QUeccJiDP+RB/z1pDwA9ZqGPEQui/YWhQ4Pm4SerMb7g2TOMFX2qk
zYwJ8FABdThsPFyYRf2Qp09WaKNV+N5AqeKXxPLE0hvtqPPTZymGWERv24zwm4NR
ayC5QOOX3NCAVKiSHm8f/jQingweKOWrwEBQTT/XodEiBSpbL6CuUtbzjHVRrVh6
iJL9PxmwGeqWt+uzGqWFbJATqbYlCKHtMAVQVoPaMXmpXkk5+fDveeX3AGYdC8Hc
W4yVYJLdnQ/t1yEKILUM8SQGfC9PmWeuXwdGu0Z3ZAUnhbnp7l4LQzmmduXMRitt
VzmynRd0S0U0ljwIauQjFR59M7JyoLs1tCGlIsDk+cDFPtHk1UB0AQwkyI/OxAZx
jyzBeN39XskY9/BtasfH25A0gilSFm/9xUajh0WtgUrE7khYvipFcwtwZ/a1xPJS
TsAgSjHSCm7de2qdqp5Fohf67ZYg3Zts5ocWvLEoCUcfqfgxTOoq8Ho+vDt4uOHe
DCz/Me7pTluqTQasClE4mOX6bu1s9JOWF2xKPsJLlPyqpluFZZB8GVAYCR9wJ1UR
znaFmk2mjee5iECy0HFYHqNGPAx1wo96FpyGa8aC/Fx9ntXalZBW1E8L233Outxh
C9V2vNdtpwzFn9KepzYKqvRPpUsM9a0hUF18QEh/hR1PeCrEl/IPUxhVK4jhb98l
KMC0u6n41AoQr//zjLLpSsXFPctp7oZDlH7l5JHEDWlNeEmJwZHIFfpqZ8JxUeeC
BVgnNxTvrchvfuNW3lUnQx9zaEptVouBqHW1hxN2W0m8NPTodU3av5xqOYkydl6q
j/b+Uhe94qVixEsItr6DLHhd/U3afUsOmNcBkr8esxmdLfRRpx0+CqSfMSgiylE4
3nuf3I4+INgnmmbAGQPr9ppvZcHE3wkd1Y1z2ZX3xwaGDXpRm+cBYDq9w0IMjv4f
aUoNk2QXGgGq6B6f1JPHbZ0dwDjICUsUCUYzTeD4fu7ouikss0yf0aI5E1fM5xCv
uOu6krpDlK680oiV5xx8M8XEnmXn0kem6W8sg9TWvsHg/YFs7TcsSXItvHQ6Tx4S
m6gnkBTjMX0IANktoklofLMVHhQ0bjJhHZE4wPQpgwcIczex1oaNtArt84+jahGs
2VbzU7K1GJeppSYFnmbnTMPZxMlsBjlCqwIAfI70mQvciMEVkTJ5Qngh3JU5jThZ
s3IA+zoIq3qtcwbFFxBNatRKysN+fLcvCm+8+CrIT+vI/prwmYvNgruBxbQFaRYh
s6MCO9ZtTAMLcyyIYQcJDFK5lfG5l87mZI41cBNfwP+nLmAnl0FxwKQDyGxu8ez+
3YjWK2UQPQVpdU9PxZSlaO0CwLpTztfS1RHAfA+6O8GCMpCeqWlVHgeYmfQo/euC
nl4KICzQbasWMgMpxMpyZhaFAqtYTZP303YxGGquSWKUXVtx6ApAmK6x3bmMYiJ5
xrPN0KugAAbnAgNk+XIyJeqIi843wJs9UhluopD/V74r7yuXEi5PLSKp0JN4vKnR
0w0Wwn7KihmzdBTlQc37iRBUhcJMCulk5fd+CQIBt8VPOs3VX88azNhRTeSk8Yuk
uFN/T1lgUS5qSRnIHYqQ5ra4B0bgZaixLVQEV34eDoSTTrxdlNmUNiFjdq/vl56J
xS12yFJjPFmlDR4/b+4GcilTRXx1CIT55on77qNsKEwVTvYFyrlKzIhlUxEyfpzf
Q9ukwkm1G8loO7kBSFOhi6Zes902+5rsisSBZb+Lt/rD9cLCfW6XHNleAu6D6k2P
P9I11lx9jPmlqBk0xERL7MD0L919czBlmGtOQVX4HqnNy4U0zbIG3D1qWzXqMy62
//h6T8yeIRxftYe4A4qABtowzktZoyVBPAPMizaHRt+JMpRj7OjP1Yrk8xhc5Uqw
ecedmIxYPCFDDOfV0dch9p0sjF+Ua74AIub5g3vh9dbfdq3SGu7DcRHcnWcQR3dd
ehriuL0N4p/pXMK0merFaRXw6IVAmFB8sTZwG+ioKQKKOnpiHcpSXv/P8cM0LZO7
yuaP7LIoKpap4x6EjDRB2gBw6Samz/SaY1XFPl2dTB+bUBocO2cw6oYbiADsKhUe
wyxoKbqfdAxnDWlHOQLOB/8HqPKKh8RN8Knk8kal26DfqhAHUKrtlCWsAQjGkyvo
CD8dN5XAahRG+4hBo/AmkaDZQ2oK34Fk3ZoeVNjanEDkV1i8jo/NHHXf5ECRmKaX
+gu/6iRG+2eNpJm/H2I9Zb4z8BTAKGeVWPvEH6jez9bJLn1VDgZOofLZHBa7TVaL
QqU/b3lLa1eSuVps+13Vv8WbzvVff+3YjoX/ylERQg52rvj471YkyKbQIbXxQJmf
Be4vh0r8MfXrx1Z+kfyXn2B36Gqt6iXheyyaPqOH2girshvkOBzrsoK//tU2Ltr6
W/TIhKR2FM/ztbLE7vDbs8URnlq2W4/Yw0LaxMjWOWQ7/O5ES7PFtt2PIjCTPiR3
q05RfqkowtB3QyemYyy5nrkuuYavRk3EImGBpONf4a+JMFAsHsFd5F7DylLYle8/
YVS0goWbaBhTnsycovDpI4MgPflgD7mkoIejwMTaTG+1rewUHNPePoOVO45rMJOS
du84isPLBsWdFh2DcBjLW4xza0z6hKHAFBlQt7ZE+hwU+PORuMp+92k7RWdyB/+i
igQbm97zztHTpR33SYfK43+MZ3Z4XiD8ZTpcvrJppBDzA+OHPrNZvQbV2USsYQTP
14Z85gBdCMTvABeOkTMM4Fz66+kMafL89NYeHrACVw0fztKklLCx8GBSENAz2zaK
Fhsq2kEjSXvdZl7kMysA5Umi2QByoVJWOijwucuf/IGYxo2j31N1Ec/w8DnMn8Ep
tA8hcPmePx4nC/EFx1q9UHUX+PxxPowTZaE8PHBZyz1tH5w+yj3qGdhPHkGHrwOs
65iCfB2eB6j6je6wQ0dGF6cRnCji4jUOZatfeV8hztdhE0oEaLd4XYo4LKPsbUYZ
doliqx1aUMjG+8Uf0gDofis19fXQIyTKYc9a7lSsILLUwBTvWuDB0Sicxqb1GXgw
V7sTsCIjs4D9IhKnJDajaKzegbiRNdyp+WMoxFBWu+g/bkFlTJnqS2Az4hynldG2
pKLlDxkm8waLxVL6AiPKXQDqEOXH6/mDVxvjvE40BYYx0t9y9dI47U/Feqrw+f3T
vQyHRVVWoIpKdWK5zHVYqOfmyyr5s7Ywm96clU/mPCVDsZRtq41yuwrNb/wW1ztS
l7qTsNlypcyVetZfDINPORiX6MJ6JLKSX9l9PcNr7w4zIv5JMy01dMjF3ifcF+3/
twguwKjkjZCEuSzMhfp/8+lMEe0ZzvQOxcUWCDdEtyztuRQfb75brWpFM/cKx7O7
o264h0peRj+1xpg1uca5x/5P2AiMyFu2S98tlAeOARhIzz/em8+4V8y3xt9EI2A1
TepY88mPbmg3Ka/+pG6Wosy2mKBb+k5a5IRzI4uC3BwkyhmDjnlgytwKEMKPC0er
Jv+mWnYM4wbRuVfzujDUa+eD0qtHzHpZqeqWGVMgb1P6Zskk8fLNnqSZxS52gW5F
RvCQZi9iibxS9Z5vFr1jCVjX+eDI3/G9Y6NANSVPyYkFdsmtyeh8e2obOuZrB2wq
tlK1qrlPH447oiCWsj4VWXdzA6jYqFBhjoO1ad9JIBRW3kHScbMy+c0w+L697c8E
Es1d2+FxhAFN0latIyprgRRKxw+pv7t1JvCwQQ+vXpf8absCbsnlre4BJUZcCkgW
2Cw4BP9G7bBeAgSbSuDzSMpf6xNWV6UvyrpYB2X8yFTjrgEUIFbfLJn38KQUxQFv
Qk3BgdJmxExYAt1gQ0rrX9xoeBInlAI0zdZPxcQo8gmmszpdDDWYPEkz0KXWL1BS
ooV82Wm22nJsIBc/HLeTw3bwAF1AOHZAlqGnIV+Aa9zzHGTIJC7qvoia+FGi0KoA
q2ddiIWVq3l9sS7NXFt9HvVJpeeDnwRDtLNsU7JIIXuIOVEZo1Vh+2ywuu9uCSHJ
x9k0+IiMUjpohqJyTEjNrHrcY3JGZm90PCvvHo+pturJ4h+PLWAGxkHed0XpAXh1
yusK0Qkz4ruhF0vEWiBNELqkJRiogI+EkaRqHRPTzQ9yBo9g9VYcJmc+qDxMdyp6
iH0rB6RIOnKGDIZf1ARY6yC+0Su422r1lb149QFLM30mqqbQk1oGSDf4UvFQ0zPG
uwBLwPrwVisjgTmKnHLD+GOR9SnEtNB47AiLTaTcDSPGJZ0zQknv0YEFCjNdjkGL
rWZcet73mxsbTXJ60tDrIWvckIiMCdkWxxZ9y9KyocRW/qwmBcKWMtAmlo/FDQD8
mzLlK5xPmGDTzw5kMa1dy2Dh3iknqKwZBJ9y8nj/i3TaRi2XbPyazuB03jowXkXX
7WGw026Hp95dYuSnGzTZrW4XD/h2DCC9fLujYXDAJlg3U15zVzRHFtg9uEIruizo
6ERcS+7EU8PFq32sqTzPxSKSpXAd6abQNdet8k/pj5w/Q4g5C6u3WN0OMZ79N0Mh
zlExqJMXSMODlTZ1rX5pa+MBwN9esZk30DjPUWvaJ2d/dhpNsNNCOiLxnDSDvcHa
KQPWa5B5MlLQkZIQ0BQu/TbsLRV+MRkxPKSbMkddRb9w95unFUEzYGFP6vLjqZPx
EUeBjwU66YudtCQz4OM05nzGcbKNZxbIGvjcniK+22mtfWWs8sB5Muqg9flTcw7N
WE9KTds5uu3Ote7V51FQdLNZRQYIrV/agDX6Zj2SpBz8fK2e1SYDcBfgsB0aDS+0
J21iQvKtuFRt8ijwC+h/BhFKks7GUvCv8FuS4lhvmOpsCiiulUas36nCP3matxWg
bE9A6u1NqIb++uRLHv3MS+XqcKXu32UgpqVWzFAwImwLb1PX1fRLv1D4oPRb8Jg6
cUULZApqG56muwXMtACMzGPFlOxgzsoupurbeN4q+O+KyEhSlBThmp9jKdhDGtJL
qrbqJQ8sSK0eGuhC+ovricVJQykdYUj6EKQfDZqkGOHcNViIO5ussFDUhsHq16r1
zBspesKnNVdyVdJmOQn4h6Tnx2MkZ5sff+M6cvO9Ih8m9F/YUoYR+tDnzfew/5Sr
QEuJvNKKSaDme3BYhIQlY+1ykJh5DtzmEH4BANQnCqIAHxaJqRQDrsDFWbNFMVkI
jk4k8ReZGMvIL/OGw6x74Bt2V/iJ/rXf+QfFsWdQ8hTpfAkFn/uv1EXGD+iASo4b
gHE1FcewpvK7c1bwKWH/ZEFlPtbQGMIus/MJewIX1hWFGfj/TPDOwsHD88zj92Pc
LJ/38r0KumcvS3mel5kO2cY3C6yJGmY+f2DQfzwTONw+PeJBe5/KebRxxoc5zhTh
Feeboj/l4atzhe6aMdrO7z28mCpZdGe8rtsVRXVZN+OXeYWoGtgSZjwSUnrXZNqG
9DykReHPzGAhNvlIKvb8ItAJeFz8hjOMVuW38QGakKq7LDrnO8wVdr5xqGmUWUI0
+1Sem1SDPFxHibdVmNsrpUjvywlPaMtQ8dypSJzYzOwjOkC6rPBeQcBcdm8hgfp6
RBf5WhUTxZA3Zy0T1s79F1xefGdHyN1U3AyB1GV3no9YrJDYy687pIGJG/mcoBx7
uxfE3QC5X9xa9SudHpYwlupjM56NWPTVuSkHgvGZUKkfyvqzRZoQh2IlST+xAix+
4FuZOAdP9Fwi7IKLnEOS0c6fZ5As6b24JXNrvb8eoEo9GfvSGF1Sy55cxrUri6M3
dwPOieBBQwrE8BxiD41whxAUUXsBm0QxblpV1FRyeLQbryuGxPvFrrMYcIMYd9PK
o0/tglHDMGA7EUOmTDeriZ01myL9xUHpde6J4FLRgy9pREepzIByQciyaC1kBrVb
pvRbwObDewhzy3Fb/r0gEABXQ52G++ilpcHHAWabRHi3yfiSEKhcxzJSuX9HmhPU
HYsU13ei2C7Oa5iEGCYOK2D+cIksyMie/OwodMpvgM0OyoK83Is4iX/kSkBmVQgO
RCpuNd17mo1x0UrUv2aVVz6JeDIwI6MP7VH5+Y0VS3LFOY9rpfiRQcOWjqrecosw
YOIhFwXZloW+7ZZxA5WkPyXTk5iNBZdNIbbwYtYZP9lGE+EaWHLTOL/RogsYnitc
Qvp6vzr8W48APp7dfueMVKq2sRfbe1melvZuV792kbwzEpQcl8rYroZCbRiNpxAf
oVIx0FSx1lRJ2/CqOnQhjbayiE8/9wxfSFwIBCPUIC+TwZAcJglVAMZm+DPSbhlw
6USjxbRe4cXteLgCysDJxHW2PkEEBoDdi2KbFyLhe9IsMj7IWz+MnF2Y3lBdqJmF
KX8wr8ipEdpYEcwHEnTx1myZy/6f/27uAecaVhzKkGftoT9Oe7I30AN+d3sH/ZiN
pQtQbn5M+DZdSwnZSIECFibbJZ90oKhPFLJRegSWh7wq5IqxvwIqnHviHlndqyeZ
0Hw4ba+an25a9dmEvPy0dLLXnjBg4KdG5NiweV9DQLfa4TN52k1x0gTMmQfujOEt
2xzHMAEZ/NxxDH4+r9RmcWIGl3ib3VvEi8LV55r9ZltfRxJVmOPGT8GZ8huGHGTS
IxHMfidciLL3oQbryro3SkB5FxXSOwOHp8zwQ1L2kYmwwLEMAAjIehgXWb5I8wKw
GG+Rx1HtgN7ZZUYTJETm104MQkPnePzi66qfattbo64EByxkfYuafV5uAYbsVYOu
3h+aMB3fc0pChYgPNkVWnQVFrAcpgZ4GoCwmONuLYMuYIp8V81eQ223YJJey9ZMA
7Z10qPMxL2TwkIl0MRTsaDImvV5RldhojmB5kB6Qk30j6hKxh+YtXK9FkhrhmDfb
8ih/GbpcqV1DuH7JFxHH0P9Vu5aKoZAUzrlzk9I12crmyWSUbzQ0bQB4tHPsGKdk
M3HnuJNJ26+dPcKl8VaR/AaIv29mSJVYzqt5EByCwQMpHOZlvPMA4YUIKXWFj3B+
YnT2yeGD/E8YE2oSBfWyOuJd2RzBFvvYiasWuAiJT6+vPN03bFdryqXs+zsE7MJP
GCAI29GQvV65stPPWZv/4xZdn8tgLY05skAhIlKx/LB6ym42SfQdPtHU7yt2BTr/
BHN3YqrrOqoqKRMF4znyoJo/QelvOlmuyrdmaes2iO93Gt4Ic5bxb7KZHEDIJk4l
SX/4cyBFmjiSAQpeUWUut4KT8pV+qu7fLDuiqSZSlW0PKIqV2y8WBAlLwQ4E7mcs
T1bn81+4Ym3EFkfVLnspCSLYq1le9XIUrxcSr3476IX/+wk1OI+Urk/xjXuEN1IB
muAW9O6peSQkt+cvyWax91/01BLtWDPJV/tS/O1vrPPI1tuP0OUD+a/0DneQh1I+
mEFrlcOGyWpZaiqO733NcR4zxuaKI8h4vjr9rSCbicxF+MkrupabAtWcTafP8AQ2
BBSWgPy5u8otBBk6mCmAKWHmb87XpDfuOzRik5dktZwlgUAkH/qskF4AFJ3OU4nu
fZtwWpkSDut0Ro+APmqPU81zatGkWeP2funwTCkd7lHPMrdO9iX7/qxlFfh8UpNu
g+BuohbhpBMWQi2tWHEJpzGNIWRjoL8W9LA0ONKxuzrguToPYBMyvx5vcESkPwoz
NxIpA0TMV/dzX49DFpXyGnkc0o5JjzPgxONgCW4W6SPtkf9XNitM40H0Dte8EVm/
viaI6oJXuE+AAI3mi63DZhgWuiJIJ4A+ux0UXR2G/A5XNfIgCjyAhQLO5YUXw8c4
UujrkMiYJewaN6DeDTeIP114+Oy1hMJWwRkSfw7IXCXL5zYlUQvZjV+JKjej7WsR
o+uzmkpf8p+XGp2a7wm4MFpX01I6yKhaydkDfT2ZZm0qDurA5rtNdYgtKruItSOW
MK/8nnHlSnEUa7zhMdL4qLpr6grXQURwb5SEuNosxxa00raQ++ctiSSHsebb5/Vc
GSi0vEFpKfNbwXLqNYV9u/hPl7ZM6x+M6irlDZ1a+awRT18J46cZ8P3st1CRKYnI
+9lshVxnJeE4E5K8Zg4UkmbvGULNvrAvWunQrDAFsleaCwyeFFuKEN5Z+L85UhgK
bZOZ46WVRlp7J8LxZBILGt6QQqYJhdQEmP2gAGPIzsP1ahQo4QXvqIydLbEYQzXk
I8SPy+rq62TQtTx7s8jn7ahSuiAFH+Z2nF8BNBajH/+KvbQSCJw1JzHtlMCyhReR
kdcKl/M9NUnTgvFnprhA0N3I/NLkIrAiB39hwpTAkWpdSmogJvaXvRmW9gBKzghW
TXQQoEiMfVJt7ltjbCDr2iNu5Ki6fhwE2hHdzgNj9m7ZHwbsuq3cS/5brjCSRMru
8p+2TAlVqsGAYPJRKM0GUini41ZwcO4jumz40blVWu47GIQ+Hc1E8J85DGf/fA3Q
3ICEryubkC9HCz2rVq/ib4KErhHwAkOK7huJRvnfWxEuk5nWq0+AQE1w+DIJQb5C
gNCoHhrRIq2IHaDVhxIuCVfFsPOnrfhtsRWusB6jUbt08Ze3SN5gda1Ul0jT8E4h
cGYRvwYzmJUJFduLGedF8I1jWMXsPAENhs3CKQir43NT1PQaJ2hE+cXDEVq+0Ang
cBVhAMSjG8UUMqzTPEDNBfhl4I9z20xEZr8aORQfnFE+hRmRSBD9OpeDsvK+I/sB
bvEktpqhiHo6VjP7vzXP7MXArUpnVSMNMjP4KxzuO9mw3JtdmvGJY0CDW97TYVaZ
bqm+V22HCjiPAdW/SZVPL7ujSEKUnw5d90XhdLvCkG2KDj9QRd+a31Ts2LzQGZ4W
T1TB9p0l32xWnKwnoqKCd+EVbNHIKcFAuqxQzAe99f2ZgJAgUJGQKSkwXIi2bbCz
FccKkl7+Uv5Ugk0xJZwHzhaSJz5ycRWty0nzDyRTh0GkqQA+aiiIhhNEKtGSL/tD
zH58YrjzmYzqCCQpQROoriKPJ+9+COs6iRflHsLgBdeUaTUiOBhPkG80wz9NE7uS
CHt/lLeAQs17sf8zVLutEyLsiJ7OrtY8bJr6dg5x8I0pl0nGdyAidk6BV1fIf7Fy
cMgVzwGUsAZxmEDdzLiT2/vFnOarJ6f6mbo3yxb+pnzmBm9zeUUFe2p8UJZVMccT
I1kmdLZcCuwNeFKkTcD5WEnvIH/kYL3tDLx8fS/6q40gB8yN7HOVtivXTPocnoRQ
m50iRh9fRXxqtDJprrx5zQIvpfFesEz+C/R2tamnQOo+4Tgr2IQOHHvw+xJRZs/M
i+MxbPU7O7fK7ail3LvkhcQiusWfAi30gbQMsZ/kcnLWRCiH9uemI1JKgoy5rctx
FDDZ6vq4B2t77ABTfnqKClMNkmsl5K5Od1QvIVRV65JfGtzaBefRxe9GQkXcXtnA
KGjzm2n2Oi0TYeD/F6JLz+5l/mnOK+tXhBhVzRUT64JSkI3nceEwHbQjBkb7sjc7
nSenTwCPjQRytlVpzq6dMCdlPu+DCgNunoUdRXMZx8uGS+8ejPI8sNfISrEcrwBm
+1t/QTXzlVSlcoZMHmiCO0DUEpYDPq6q5V/CMEBh3Rtt+LsspewhjCRkWmHstFWF
FXF46HGPqb//DxDTad0lyG5mlNkn3YZ7yqmNe8GjZ/Yg2+fCxG7Nc1qjdqUa32JR
d6+wDIsGHYckRv4byKAmefg8mpWwIqqOYDYXtJ9bMa702Zox8zvuT3CMeZIyIlDP
Ozn7LeI10RMW678lNROHNGwjwDx6fFrSDEmmvpGMcl/wUodTA36/WfVLeF4m0OFl
hSXmoLfah1XsrI7+yOa78G1fFZ+O+bFlK4A7zhqwCPW6k5yxwfPIwmrbimrTUF7F
YqBb1LP5D+PDdqWJ0ciKER66l0gI3ICZHtyS1uZVFutf7NsJ8l2EE0jHtGg9ZO8M
jdlo4JYkKjdWtSKBfvy2gneQF7hlft3UpuJM7cRigJcR62b7MYc30IfFoIDf8UYN
S9mtv+akKx3Al06fPJo772d0lMIvUurtW5MdHt1CjhsdOkCNPBBvt1wvqLpMZyvM
rhx3cPUHAWNV2brOS+akP2M1RBAfL77PjknwxwJN6SVNpxxoOcdvIQNt8vznGROW
7rkgm6SCvgTtXYNnxxp+vsN+1TwdF4h8PXqO467P5SI0HSg+czNUf9/RFDihwtZK
k9Y9QC0ptNpJhy68mtsQUnIfwLIaGiWS+Q25kW8PZZLalOAsPoanIAsvp7CJYscK
0i4b1qOAT2AdF921YLWH7N6rqaHR1TPflAVf42hgVZCBHiUYePcT22VRoA1bJMiI
FEuurFglcMKHcLqZ13/2YZ6kjvaAXx3HYvr5E75Q3fSdJlT9KHSpC1c8CuhuHJgc
sGCIrLsmXzsVD9EMNl0Mfh6IzRdegRq60SzmhNv6nXCiRvmCPbsVFffxhYVfynLa
j1XigF0N1n+LCSjsIwQsTfHR56BGgdp6hAj3GU81rz0Bw+U4mtZJWWsC3Dgz1VcR
bSLsYM2QsQ0ER6sFagWwUh/Q/eAhGzdg4MV4TTop9aOXQlJwX5NPvl7n5+hJZzOv
2YdRngdec6GUF9ZLHAmneDeJKcC4zSsm4cs1voE3TNsKzt1Yu9d7dAYrRCkm3fKh
vdcxZZIz2CA3mJI9gS+xnhfmmQMi1pZ98P4eJLZOhNbNmtRSZUO/Zz/+8l8uoJQG
XSuywf2+okZpTGpayoELgtUNMw1++eibQKJX4SaeCfGq0xzOxzrH1CgRXr/2DLij
TljwfqGLgGcxpB48DgKEoe5eWWaWXR7H535QZeFcCXNzMnkicPsRQ/J0qSYRHR7Q
N8Z724x0LEiJlFvMV/TrOXnBKMwlKxCQcG9XDcEPu8BfaCZ+49hrYof5r9xyYGD8
UecQKRQCylRxKxzmwuQE1mCpUdnNUxCbLSlVNjR8TJCZ+dVeI7fsts/CQRCQB8AX
JHVUzMfTvMo6MWRylHfcv2sewcNQl2sUw3SWls5UCCyaARI9tOeGMwybVwSLGzUf
kbU3LMbYHDaA/eLs6eHGmxAC0UBmZ70IkG7PvO/vUzpLzxMEEYZomWf3JngXIdsc
2VJJdEVAJqX5biyqqZHOJOYBAAqQ5dDzTTaW2gypnv+MCOT5LREqp1y2L4dwSnJ8
1eVs2esbsogIjYAuUEZfGvYpUViFnHzrggPI7nr3MsfD1L+Nrnrb4cpTtpP27S3j
5o0IvH+M5B2Td7wGobNniszgIo/PW3A2LKUrFeggbVj0CQrBZcHG+bgktalqjRZo
kS4QkCTqd9KQXtY4a6Cm8RGyGW9la6j3k4tk2e3WcEh5qo8jryrQZMclDDQ1jo4+
2BuWTcyfqNjvS8i/df0rfMGfkKgI1hY7N2+UtfjbaILRaBylmqTBuG0dlZbfxYex
KIEkhHl1HM9/QoU5LN8GM/9OOGu1GTv+NLNWZXft5K4UmhxlwTe3k8x30ziYQ3Hd
0PfbOpHJAEcMr9IWtwcWnfObhklJIMJxsNX3Mrie12URrxl0CtgnI/DtaNMK7IzH
/SLxyGItCJCVfIOjuHrvk0dkQi1hwWQrxPIlAVObSMvbm8Eh001qCdzVnCUFO/yT
gEmGBQjs3nr901FuuhlLfgOvZDd4+5VFRGLIzPyXbcugyY6vJlucS9DZhBMtgmUc
4PXvP8ZoDw35nKXhwvmXdX+tEjHkCKvERR+8xT/RsEUE1AdriK+9ChPL6mT4Dl6J
hqxKxB3JQgX54jO9Z5QQhvukAZp5XcUvIQJ5lccYZGxQSQjNS9nVkn17okK+ruGk
da9TANstKk2LhaXfzoGqZcJY6NzdnJDr+o78KncYQLZ+8OwzW8wFm/Qc5ZxXvpvC
AaVr7ycyev6UOEnuyZ6p8XA4k3qW9GtFtT6tRLIVdZp20Jby4kSAzuFnawjqZPq1
utXnN4A+4exkGJF1TToaBgNDUDxjK0SZMPSFmhOyQk3ZSQNhvRRzpu+4mL2vSJIZ
KhrwoQvd/iY5v0BS5srqKswr1fPjKrEFFTujyupB3A/e71fnXq+np8nRfvQJXvVA
3eNSdUWZEcAkOOoBkLzyrcgHyqy+wIxfpXOq0ZYe4UHFOWr2Z4065FqZX+1/n9qG
Bkml/A1aLf/8EeOuwEZLy5Uk5JrGXUL5/brnJrRnY68FxkYIZgNJcvhXAFJdDAZV
2xAugytze2mIcFOsu0gM4onmi7KEW6yfzeyvPAa69zU6O4Q2vGEbVgMcfCJmMTfB
ihoVqNmlj9/0lGbZlS4TSogiwPmzRyh6GSif20VAjLyFkjDx9I8spe6tpqSpwnnb
BZOsffM6FriDheNpcDpTMtuUEZVWdWisUezkV2gHsNt2Rg7WeD7nRPWe1DjOnr/B
3ti/Q/qQupiP0vgj80AySo3R3/Q6DI8ZPW9E/PAOQhQnPXfPQ+zkdfOReQsn5pPn
i5A6Y26SIp5Qt5maLA6no6a3PeB2r8bl5SzzT6CzzOjMgs4BNWU6dKeCOu1pVcpw
2rf7ed++a8LU4ZW5zRh+WzaGl3yDuWtoz9TvPOAtYkIEbdcY31rodCq6+FObhgsG
iQ/AR7/w+n3fDbcgClvwHaMJE5f5XbgYWfG6vtHF6uJGPYEGwCYjQolEiEwA/VE+
nGOQI+DKe3sXk5KE+I6OwBPPyxzvCl4zFYU+B4z7V3VcYSE7u9FhBl/ICqLTbPaF
zcr1CRZcaUuEwWYuXwD7pU5HFR+BHRmIrq4G3bo2GflRqjJ9UXZeJNi3xs7QGtOz
+703ktxsL5Vl1bdhFL9uB/ZgFx6zut4NO9KywitWlslJtc1fxPOOBFqt1saksMso
kTPtngdtMfnsz1+2UmWhwEcvk3R3iWtsQgEFcv5x6qfSVqFdtcDoQEKyl/+75Y4t
Pj2p5ftB7eDXmQs/NVjPJ9cVhcW5uG2NA+zliOjtyjMJhOPRQohHoLz7Se+q6u77
b1oQ8V9v641qDoELi8uNx01Qla0H6/KIsszQa29tLdrTUvu9BnGNJQGslPiXxeoQ
dlaQuG9tFIkSnlpIRpVCKZiyczF8g1eYMD/AQx34mKpBxG9OXjT5C2JEiF+XKzce
d0t7czL0YtmgEcX50MGmdudhoqcP7GXRpVblOro5AIaiBzywLWUyooEHYZyeKTAP
SIOdecc3zyXjFmIx2pcuetQKB6h+kM9SdPeT2maUBUe0DZ3mXVh6YomkbR+H4oBe
igWUbPgc2BP4BMVhN3l48OFLMyqbYX1oEM4laL5JkU4mqFV3xfWHD2ztztGKeZUV
lIYceeID3tiIPqatxQwOeaJje2uHgUuDaTyoVznniQZxvZsy+CNZU7cu2qmWZ3Od
kxtT28a/01psAi1GKzJg/6u555mKAU3KtNrAotm5WoPzABlHcZOz1oYxrGBHKXeb
pjXkdIR4kMe0/kJW/YA6ebAurpkBUwfOB+ixoonrKJQni2euYlh5VChD2Qxe7n7A
VGnwcvNXgo3rZkSc463qGodOIElArUooYeSYFjIO4YITpDnUJ/a9mroY9iI3qq+N
zkK4ugBvdVrAHxkUrZ/iL7nwFhne0DlstHOLgKlHvzNDvUa7drJivoMgk7qPqP48
sRfsFauM306xAKnps72kCOTHQmKOk57+K/0/NPcul6RcteOiiHXBnyjhdJHnSlyr
UKqOT1ePL8ynv577R6V11IOzJAEH3kedm7GO8tKlfqXi60ZHWqGHWla0BQlN3Ya/
aUF+JcvVq7LkpEXOa56stO964BnbKwo8FtFLAp8XT0zUUFFziEOyRDmihGxaRiTa
LmAXMgLHRNq1T51UKPIc8Q4puTS/zHwCWz2lSYqcAiUcH0ILNdD5q8MbvnrPYvUB
AtcMyVl6/V4Dru+2SsBdNu/IEzNG9rImjTyH+dsoqpMaglhvEwppgjpThS/ocT/x
koigQIRWw5qqRqsKbmupe6hZF0F4AVWr4hlOuVwRu1uBPZa95mwMYG46Mt4MbvuM
gfh6hxqLYW8D57Jjb7l4+luTAfVAP+y9PTy/5yQ8Ep77+JLWTNVE7cUaTfMoCjTS
qZ5xtTA+upTNbky4nkLKxBie1vabSwNgMADxmgUx+Fer6X/CBwxkGG7Zt0+54BEX
/BQUNf8cMtAJ9yqzqRrOv8CipU5osnvh5EYUWoDmHB0WPPplTTLqxHmPOtMv293x
Q4FqaSaIBSacn9BfdxBasMEUPhmnQmugU68BLtjpd09+Aw5mewego+hOw3wwdERP
mMXqsCJdMYhsDhMocZWsxe+7S/0cS1tfgbtMpevePpx+5KZmO7iIV8dzSp9FpIWQ
CrPTJZPZQv1fbvgzeahWrUKwoigu4zFDoOTfbO2bA+FHaN+X174zJyVEU9hTipa9
gPatHtOPig29r4E6cz0BEhq1s7oqsfgt/WB191LycKFfVW5rwkFsRZph+E/Asmxp
o5A+Tl5grI7y2dXzFCJxctlv/OhydrDf8trzS4XNIAONC5UPYi17zHY8LTEIdkyJ
Ibv9lkt6d2PWwFxWO+xvfu6jsuEec2n7eACnmdj4cEHGduhPbHRAFG3YUNgsfD3X
2/TMQEV/BwTdSjqf1Sv+ETK6i2KNJBNcDaPI2C1KKL6nc8k+9OlKOAUSXwc0JIMQ
Nl4axdVMM66efKXP7dYK4ZLF9LHzmqTAUBdAD8rNBdXfKxCfYPukikKdlGA4XY+M
dWYnMdZ3tIMbko0bxL9HrUz9oj1Z3p0pbQTVJNcUmaO6gymKnL7bF1MHp331dD8z
Jz3yUocl1BIVsopwN0L1kX+OK5PBR7wpSxAiHpsKJcE+wSUxATLYi32PzOUbjrNv
EKzrVV11bqCq6Jwu8ridyIy3LKcq02lo8VxoKn/QQRSIfAtm8sNOg4+eACdLnItR
3vBC8vzJisDbPXc9OcfJP4hVcY9nmGdtqvMKwa8V6oIfnEuM+gjG67QYVlBwxFhz
zaFfr+AULhjM8J7jOpy8gRiBgmRV9C67W3IbwWGkBDtueUnOCZihM+F1cMLQYGNp
sDiyFD3roPqAMkhFsTLQ7EtF0TbMxZAnHn2ikXfAuum/HiLvCfIMk2RQnbO0aTWF
hKKIJNZhKjSpgAcmCBM/CVnGlRxrUc9tpkKjVVwrXH9OGbSwvjQ5SfEtrbXv93J7
jK6WkMa9nvb5OkC9n5CcwoywvvZY/92PQFp8QZur1BnF4B4sVCce5lpYl3hLLq7X
WqAb+LQ9Vns8a8zLGrpEldvL+M5LjyUqJvTPyXg5gl85PyOm1dlIWcM/3cBzGLL+
zbBBqrl64pyoXHpDn1YT88BS3S+LiuQ9SKEGMCWl2rD3UV7F8aOTIUi3pOOehHVR
jXOmfmp1ycZ8ZWJR3zb8MPO3M5KvDkAtabPsA4sqgJYwZJuN4ZBrVFBCkRIT4bBX
6qiPaRk45C932BdsneqL6U81mTlIF1rRZaqTKYxCSfErzN9/S5XrTqcO0bqEp4o1
RTytP+hj/h3Vk3MWlC62pUABMCbAShkbrr/XwFmjH9DzvxqNpwNQJyIHGQgJAA4+
u9GQPuqDcZ72mHGfRj1dtP4lY+Vg5obz6jfRxiRsBMH46NYZVaSJ806MKxwhcJge
T4cob+CNoU/QwOxh56ZQgXQyJbvz6rr3xluw2PgxtzAbqC6g2LrS64gYpqluk7oY
zy3IQZJrvpCepAunUrQejHqZu8cKa07Ajd5o95Gf0G3sAmaOHYbTyExTuIPDiFkb
TL6ZsDMig/pWZ+N2aVWGZ2cWzMowKe1ODOpOmIRCeXMiehQzfMZqdAPNunC2J9Ji
OirANu8x6ABv23VVtAPnnhzvkOn0azFXjtQ+IU6OGEe21y5IIULHqeIUekntcKch
uCZJKvLJtSVIpqJ/5h/S5tvgNaJEjXPuPxrxo5tUjcgPGaoNJbGSuAaKWxJFtblt
Z2ZN30ZuIykKdlNJ8wg18Fr0dhsVe5JNwTjz6Po9+LlugcCQC5mNEAXUrxtoNXC7
B5jZqzNirVBIFp4aYpsIX25E5o5OO2AcUSulv3d7eO1BINbp1bGrjxGWSy7jasbk
kFrcH06sxfTFW2GVfGQ/wfIIskROZqjBn4hfWxRLhsTQNp4QayVWm12XhubF+hn0
XYcOm6G7wPp8QfjrziNbOtpPEDI3ahfcE2zTVjCEubuHHIN2ocUk/DueVOR9YV7n
Ze3gxOLTBPk4f1XwShpAVULSR0TMkAu/O3PanIkaip1n7H1Xh7eWiorXNQIi6DdV
j+6MoG+SBUzXrxVoTtl0f4Cqt+6jOYVCHh4J7K5LDV6ij8h+zkMLnxKp1py9Vtnl
cgYLQoBm6p6hu9FHVVsn1564FcdNliWRKK9ZaiEKC6AerplhcLt59bBs5tqjl6HZ
CjC3peEkVadb28PL0FzG7ns11Ak61ibGi/FaX34n30O8xoEts/lWZLUurVMNJYAH
C+E3p3/AXYR8oHarEkgQbQZx+PbCdemUQs4HN1r9D9JWhwk3cz3WIW4toHzqmw92
Qths60Q9Kjz7ZshtEdcYDh4ifALZ0sdtDd5MVVlnsr6QryQt8PQTni2lKzWdb/S1
8ZR29XSG/hfzHdY+lJOgkV5ysJyb0YFlFJXVJOtUQ5GmbKtEYLdH+usQ9sfydRxS
3ueXX9+vuFyjUbQH/kbeR4fQUfjqQADz0IPrNaXuUYgq6dGbO1PyKUhTDalLfQLh
ri9p8yvFYI51edtzGZ6HzFn/OIeEEwk9HFlPFrMjUsZB4d5sPXEpRlMWkzn3ts42
ZYzzTdYWdoSjIo1XXDL9n9CpwChwkgelM/YTLVuEUnNY0q8FEk9drhFCy79UhRN2
NA1u5BO+NAzDFU4yUPGgh0Rgr1wm5xwcAPCCgj4mRzYPZryIB1xz/P/k1AywSXWy
zH9RgiDvIdlNChB/5Ri2pAOYjPLcg/Rx+SD3kszGBV0cZ4b3OAGUGlt0luLmqVD1
dV2njvPLMBkxypyw0RBP/ylIt+jSt+73pvvkB67HHUBGejBMd9ay13mxXq+88YD1
7dM/z6V+MS+Hp95PXijQ8rJ2SlVphIzpN0erwUMGylDXYJMTebWdJw0AhpX8wE6w
411JfMQl94HAxqG7QCfC5Zcs92fDOzN6H5guo1cqLKn34E3eDpi1gCenarupfdIn
aGPrTwlpH4bZKPVcQhaluH3242apThKD70CpYcKMxMLTXk5+fNo5p0xnJOMtuBr/
xnMryRSrrA4epgnPp1q7ZYRJGCrHlqHnHa7CDYjtb7HnuHHSVDQoJvEPGDdsp5IM
RnR0/gZ4TuOJRa/ziJQqv1EhXwRBfh1RhNiZKfQHJc21cCTrk5efenO4fbvel+zL
nEO/+NLPcL8Dcgq2Q1/VIsSn6iVXThBrTL0dSukxgIA4a9MBPH5lcQH22h3afXl5
m5qS3maz7sCcJlNHnxt6MndSkdMzkU06mBd9Btc0wXtTIa88RYyH6K3eS1prTymS
wDpwAxHUVt3PCgWlb8gdReotJeOX32+SRYfBxkNdkVEB/Uzg2OhqOHNuUKh0eVX4
nqIxoUF/XwQ8kOubb9bWfe33yRB09qrt/4dQufUL3ymfPMXZLhAe/VheKzpVOYx5
05YWp7fTzYy1i2z+/JJyVCameZtcKDgSjoHSutebgIy5HPtHHRQWEtuUKocnJ8Wo
ilFdGS8zzmBxrb12ciI7i7HpqZ7wJlR0t4Ykv38SKS/SGkgE7HktSl9xe+Xc61qZ
g0D2QrNbtVks1/W9nSGia/jvZE5t92s8ftnyBfRZ6FT6rd2oReoq6/RbEICMdFYg
RNqc8vUtqevIj88LvMXLaTARCeMaKIwbPjeT1MXBacU7yMVAxBXL5NL2+jCc1oAr
vuW0a8rBrup2SBHebjN1xufaNbwvJHzfaxIQwT01vlHAhE0QQF2Q3bT1WTkQD+TT
b6ttg0c2E5Qvv8NzKgmzfuAbhp2MvqFwy7dScEIWzFU=
`protect end_protected