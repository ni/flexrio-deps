`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvGvuPnXIgPfeTrv0s4IGtKEgW/yR+wOGzKhnvCFCUK0y
Ged/EnTG52dYEz2IMPo7ACMmLg6sDf2F+QlM+1fxrClccjcsScBoR1EewDsaFpC1
hlaUCWXmRJcbpA714sFQnEis+UupIA5bNOTa4Bhr+F+XtZipuSqzZncIhyIUakMf
MMU4AdU5IiMxdB3glk8B/vgBZS20s+Psj8Tgvx/NwvPqkGiDLOU2+Prga+CHPbr3
yArECPNNyTsD7BulDDGoypmgpgac6oy8eyYJ/3s5SAxGGB9Ife3D30vyAmz+HCtb
fek5S+jvD2kyfjjhsEoqg7CzrWHLc/IrMyTssA8NU4IZU9KniKpU3gliXWRFLgBi
qat5dgsk6cUFRmPllX/dlN1zIBb/OBztPWuEV0a8tsNUXoZNSMq/IVMS5E4UFJJm
UN+WUM50Vv+7l1svJQm6TwkE25g8yHkM6V6gBOFkPdGli2uNSfsgH7v2zqxkQ71e
lANJUd2Mv5Fy++rpd1jC6J64BcnLvOZyPSqWnEvY84tlPYAkUgEvzLqbF8n2Vfpv
Ov1fa/1tIS8a1ceH8Blmoe02mNmp/3VMnkXowM0SImWlzQWjLDA6nGsvNALoDxCV
fczfIyvKv0kS4fg9E63yzDOrJdJBA9C1cuSMZW9Kx6X6TqFCvxNDn/TlE/h0Sdbd
ClclD2thTCcTnnL/9+fLmcrc+7+GAzqLKOZkozxeapkwvMjHiBKfjmsPywYwR4v9
L7lCQCLOAoUg2tMYHEDvzpNvD3+k1+0qH9ATgN68O51pQ0UmMpMciTecjDnNU+nK
t5safJ9U+vCD6gBm5b/ATr5QJ0chvfnhG9lj22G/6kp5WfSNxEPfzu9TAg6YTFmd
gNGK9XnQ97xGytx9zbfRevBhM/h272V3TWOBpdmS3dHQnuBoUKpRK2kEIGvmA+sw
1G9J6ChTyqjlNN/W92HGXoDywlBNuLMy3mpJautU0HlpDCYCWDRq2icfAUT2mrnD
l5/FiRJ8j5Lys4iilskqfRk9Y87QPtddV7lqdpJaqzKP8H/U0wOM1HIE0LRmDCFA
xowgii08jPaweAOI3J3UEWCd+5iycjTAkwHtbkYU1rKqkfzKylaGFGvag4g4OL1W
gVvWVq4WKe63ve+eiSOMRPx1Qa9fjmOJQW5KutyiMo8DEji3zKgj2FrEQ/UBWAOW
EmShg+epDN20ujANghS2IbgdPefuvJz+aPrM6+YMfDf0z0v3mt9ixx2dCwK70duq
DlDNGsh9ezC1TfJFO6/xvaGue8Sg3tTJqCCYgRSqvXrus12twjYYe9iFxVVAWyXJ
1itnabHeLaRvTHmagiS0usDoaTMAo2OaUdyjDzyApUPZwmQAQMOj+Mob8+Txx6fb
d2EuvXu9zeXkF2W4uTLsXK/b5iX7/Ieh4cFvd8B8KnZBtzrU7bmMORYlm+gTUyti
v5qKOJuUUPGyQP1ppmSmD2FH6kbfEPxQeapiWygtSiBFcjhPjO93pUuvrIpKiE9y
C02DW5WzQ5x7yMia4+eGy7QNrNOVus+zuDx6bG+hWQpMPsUHQ9Dz8iseQg4QsrzC
+bRZyHEzVFZwuy61CXR2waLWrlnYY3BpApdvycflHt+g5il8VgeG0x52JIUq5eAp
TRDsO5S7vbGiawJ2WWzzvvsrZp1cDNSVI1onSuu9/AGWk0SFFvVsSd0jiABdX3UK
UJ6TZ7lNH70NQ/WMK11CecIFcV6vvMIMQT0zicvAKVpIgLzvymJkNRD/p9X2Zqlc
o9ce6URu9VCZpLD59qOkQH93FFLs6SR66urZ9Hnb2qzxKYLIvtrZPiJDT9jsLBC8
gcWpvpstNMJDk1AWRtKHPfl83lItlhYvdcvK4Zl+1h0ualYDLcB+TUqrOHFpjyKR
TPYnMZkCG/vhquYFXCToNNNto8Sj4ji4eYJ8jbQLL6mWv+EOa6JMkpMgAFm/w2Q6
8ZDV3WQqYTv4CogJexF3I40iSmEM+/AFFYTxfPhCVE8NtR7/lMHJPN+deMSrQtd6
8Cxqlr4leWxIpFDJKm9bHek+2SM7IrIVReSHkUks9DafMrNSthpLVeMLRDAxM9Ms
eWtH9XMierwQvvaHrOSq4nIH1U4cyF0U0UR7RKl35SY6wbiUwQknzgwv5gvWBpTP
4dx3SOpuZ4UDNVjUu1wOMCxjLt7fHjQNb/y0nMI/OTkJjYPSZ82MCcl3BjI9/b5V
r3eON3YeU8HwuOqbsl0TfLTtFHo/bBD0R3arXwLIh4YdMuOpcKKmzas6SM/i6CKE
rF8Y/Gn03asfORrIlt5lwoR2PtxUBBTGCCnsydPiEwgjAg/UlnfiuL+zLQbqqNVo
e6sA2jI04pdDgSkgaLPlCPN/O5StYKTRvn6K9oIExFAPyIrkx3laki7DPQqNHPMP
gAC1akQVNXNVwWiG03L7TaBculL9RS+D6JOdxVJwmS9QI2yCSNjzW6rnjjAzQega
eK9kRiMGXqPlCcTg6n8hOXGpVW1u1fHEUPtviR3EZyI4nRaQiTz4ooUe+I6pmBQn
VoVciZSZCqLnTZ+hUKmg3O1T211xMjuN7IIr0nPljsTMVw6b5XzEqGs8aEx0iT71
4yssu5JAiFBtvMXEdN4IilpXP+zSi+oealKS3UzxA2E93jrUfkpV7LbNzP4Tx9Eo
a04Ijlmgz524bdJo9qP8DAsRKHMqH0UaFG24KGNocy/X82Yj1nE1unieln3UANjd
SbC4ZMNxyF4Nk7Bbbno9z4PGsZgZKKwa6agDIcs8jieST/b/nUCRZnZuQafj40QU
r4sXK5BKPayUwmV2UoOufuFD0fsav0o2ezoZnlWbI4g48CkFdZoyRRW2uaJeknyX
ONCLxmBuDKMSOfUwMsFuw3fXXtZLYWd/gbfYHYqrIDJ6nE8nQWifmYnzXOfxs0HU
PSzszUJatxPCk5k4ln+dYZvVJkq8LOH2ig1BrOsCavALjNnoQBMizHwr3wcvrDa2
cH4Jrm0T03AmWUw1DjuznE2e69j/lRlQ7d2NU5pPQ1lxh4aG0JPRUKGNTs7OuodA
c3ALhPfGTw+NjtnUN9NvTnTOVvt1zNwTiGaC7iEuxOPt8SNyOzQ3JfOCZioJmMRn
XCGBVjlsutQvViGhSj2/sdYOS6su1Hu0eKiZ85YQQRK3xcJtSv5ER9mHNCAG0/fr
845VikkbqIiHa1LdVO26yUhsHxxB2+LUHQwXD80GQXGJetlOxlMxZwgUBRXyhnug
7xTAHZLeiOoRQVpT9K+s5zrMRmFZ9VSP3XeaPMAuH+txx94QAnZx7pPCQvZ+SFGP
XtCA/YFTMYVVXLpsthYPk5OIzGFUtO/vAmrkh3Pvhob59G4Z59w04shNk6xXukkJ
kUZt+gCd8Ey1o25lR6MbwLoX02WUO0R/AD5Hkt1yyV+rqBEIpwu9TZu3GVfl/0PI
C3Pgf8pz2OAWcctUPsRdLoS9rYv+XJLY73TKW4PyrkJW4QxThXbbAn8BOTAl1JZW
6sTj9Io+qvpluSjbxia+IqqZwq/sQDDUjyBmoxpdy3rnUR4vfqigJ5PDqVzPCDVB
T+vjrcHnCZfvVZMVt8Uv+x36/hgRXCDdMeGRxbAr4kWFpu++xDdv4TfLhcUEcIZE
RwQne/pXoz/XDgAbHvJq83xDQQxzFTug1L8RKctfOP+C6x9bvsRX8Rn17jcUlfir
cHI9ql6LZSrrx9p+iXmoP1cEkAgtmm48lrZsLdptSVGDQDPdcl9fC2dEVSBKwhnE
/laOVv09L20ScgamDRCPnLPJV8RzDnOrJ5t62PIUP5uldEJRrSNct3OlUmUqYtUK
VbfbNKc92PVB9f6gYMoy1wYy6lO8sAtRc4FwAUrbtAuFumYXh6fV3OV3EooWCtKE
3zIt2I7SLYqH9rXS88rBOBIxzth8y9gQ5X7KYKaS0WbQUVPRtUbnLfra2G15WTFE
3wZavsJneFEsoODW0RPktpyWDUUKBrMrAlPx3dpvBs9w+PzcXAa69ElWQoLo0LDW
bVFxguEfY3pSsdceZ6rm4AqKtrlU8zCvJAKqgPRlCNz0KNVa7f6huv34EPHSzI5r
1pnCd5goUlKBxI97npV8fgF6wVGj2KFdG252U5jZOm5nsrSJvK/TdGXmBHt2M8k4
lAGBamXa3iScn8WjbUPogEOR7pdcqdaq2no4a8Xra4drTP4W8Pzu5+NgeOeFJ4ml
08YHpqXrFEWRCXdkrR7R3s8m8pkJ5Ih7mFhTsJktirvqE8cwAMm5lKgnsMubFIoc
dbkPi2Etxx/+OdiPDd9hEg4DtRwyTtbMKNgNYeg+uoQvFwDvKGN5Eo5aUJLDJcP1
o9UsJjJ/mbxb/aX3dJ4MNBvqja+AVIdx4uGbQpTygH5qlD0RP8lghyrhLAFj8sVB
9lXiwdi99778HI81qgXDjRaZEHB6CkaQKnQMlvmrw7CE83j1EgoXjMC9jIL9rjSS
CMZxjrpcsOEIXkFqL9IY7D1q09U7qKr1+LAF5IxDvSddHviCKzRzSQqAtktafzLX
zg3jWyJbgjIqQ/BTeHbrIqs4N7PFJCYYqCRGzE7qsTb9Km095nKe+gB6PZpzKzq7
uLW5hUZXDmxEK5bp0MDIKZM0JkCsdB8yb+73PLwiIntGvXJ9gbW1Fqx7Dm+SkdaW
Fl6XTEEMX2qvL9Cap1V/S4bhUy+ev1ezSXe1wtsD68x9bfiyVkVry7VlVRZcKUOI
5KxMAvTpx0VdC0jabv7rCeweuUntwn/wvit+BdZaOKpNZlsAOZ10ve5PTYVaUif8
TNfXGyikc5VU9KmmExdkb/3EHU8oSgoIqhRRdDQPJCBmxw1M8VQzo2yRr1JQ4oai
feb452Y+UcjOK5RKe1+UlkBfc9vRJysiq3j0Y/DnXUUs0cLRYJJIChq5DWpl3/Yl
RZJzUKV+DI/sMo1ZDYs/rJ8/dgvgNlvZju6RwMfz0tL8XvgvG74wYfR8B1vd4ymE
m4hXOkPoNiedmUKpTYYnQlS4WFOP3+qaizH+XDo7l3pMgo7pMTcBYBYP9ptMoFNJ
p8L47l4n1Ogl2v2K2xFOI14rmNDrDJvQkRRmFsUVfVOxPPOSE0tH7Zp08M2UnyTW
BL/10yHxhzQCO38YH7mvADDwQOwflmucdQGJgpWhNj34LwDpv1abl9bpad9jidBt
WNgT4Ys+1RzOlJ94CkYsb0sKuQe+SEsrKKzBQzuayDyqAjmLU5gYZwR8aUx226vD
35ICjJUsWoKa4UptXPGl7+aDKNI612/PAZBXEk3WosujIsPMaVwoq02J6gEzI7n2
5Sv372H6NpDZ6vMteFYNs19Sci2iIWxipimCNKM7p3hHG7QqSzN7aoVePr0NqMa7
jjP2HxYlIzPemb4SWyZ67ii/VtRqUsq7DuIqcb2M0aJu7VRp17AoC6oc9nh41LK2
qnW8B7WF0H8QYYuXxGVyVAkM7QxC/57D4+fiAKuHNdfGxPTcYz+8X0Zw+SUJv0vc
pUei/gX7cCNQdV+GlY/mOQvyMcgSmxGcxwSC6QikDsI07bpIRpr8Q7DfNM/jeRiR
Wf1e6P4tHM2gY+MhcpuzsaRwb2Dk7+SbAr1NA9bLTSB+4O4Tz4JA6O6XTdCi+7uW
b10hVY+vCdqmEmcg8Ib77M8zdQOAQvx0xOTvB1Pi/qRhtc0Kt+fH5yqM6cdwUucw
qYMss4ZBele70rmRG02VFxg1gdNt2StDm5WjOwJPcCp0DJ2AVuJaECzaZritSvxH
p4pEIPk4RPyhjcNSOvzwpi71YDSc6QJk6pAqW4akwQvLI+6FTh8cq7DwZqSy5yVO
v8EY1Hht1Mh2pA2cR9kOZnLy4Qx2MHZY6ChQ0y+C4QYuso3+tPVjl0qC736icFPx
xfe76ANuTzTpz7rL7E8ONvyBvJmHbjkLbEL+mNK3e78Y7SHyA8s3aQU2cwPQ8+i+
OmQVuDYJ6mxKlH46lIhVfIonvx3GnhDOBUIB99T90klF9bDI5KXIJ00c5ZBY2124
f4w0C8M0ywPJjrkw2Wciaji+BFH3G8bLreK9AwpFZrgajeL3+d2vQi4i8E2iOidd
rGr2oS4EVPumwT0gFOtsjMqMaYXpX4YGdGzUMbpLNwOKkhzPckhjaIvXQkyagfnO
DYHY0fsnG/D+JxtT3K2nuip155dQkWYYKvzjhC6lHQcgU2WTVjWWA8KgNttsw9cB
0lImCyNFB/7tUjgoA3dQ9eCMQI/WCwnODSiA7e4Y21Lb6AValRyTB5nhXZ2Xnqs5
zxz4JN1jDBwpLUV5M0BJFgD52Au6CGfL4sNE6IPQUhQfrCz5UJhJ0kE7/tSJgoQq
2J+uzaLkf+Dv9kYqdZv5i5IS9j9budcPQ/wyQQ/r/jFCWdkTGs52VIbbh27Kqpor
QhXNWeDRicc29A3e7h+ummxltuDhp1olxqfvA32BuiIbrc2pYKGY1tVpcf5Cz/s7
ZbBdGa3iGrTT/FB2HJcUirl9Rc+etCeieXaXYD0QVBJF4iYuhfv3Jz8J/7LgQ9ok
Hxa9UctH7BZu07vzRhplJ5j32scKdc2bkx+bJXM2Cbtt3STY4DURfz1PwP5TDz+N
BJOeshR0zt5/wkUHtZb9IyQisNgwR7pAYHbAD/zxz9Q7MXWvQRd+pagaOAoUtSme
mU5LB3WgKsFXEKNCa9mMRddzbvrdBK5VQxnMOl64tsbTACN2XXPOvEPQtImOQmBi
lPUW06+ARQ0eeslW3C7FQp5tnKOBFoNnvFxSXmap9MvSv6GhYfAG23n/2KbJmjLk
NPvgMn51BDzY4VXGnQMBIGttWn95SwE24xHxZVCL6yY7iyTYQ4PIgHPiSHrevYjY
/s3QQGVCw/VA7jpnGT6PAFWErZJQhYaBXnXwPyUUAPduxFWQZO+FewT1/Vqs7L6x
jds5dT17AFH8FNGTH/Fd/IExQQPP0EFXRRcNw7L+qYkr/5jlTB09dSJc7Zh+53Of
XtXUHUsDxTRJ7Pht+XrNeBItO4J8fbgUB8rgwuYscD7BtYYpf2q+d2CFj/117LjV
ODgMnPo7OOU65Ss708SBw7MXToPdpmlg0P/q1oze3Wph2nwVsb2wkK26IfUrEqG/
IJWgnzDSdzmZTc+qiaH50pHXB+UphuOA7yoOWKV/+md2NkpXvEWj+P0JDEbaJq0O
vzcLEgbN6HwcanrhfgfmvJ1W5+tRNxfKsZ3A/4CVrqQTytUyc9HyfvGrdvV8e3CE
RL73AZKatzBLVYM0wyj9ZHhd7HhGe2QYd6+ilhrNYdvfu8B/9k/1Xotdgb5zCrhj
RVIE5BeZSYRr0EGVALZB1arjXKH+alGCEl+IdPfH4tR7QBk7oe4kQruzt2LR7gTZ
ZGCqg1tGsAW8hl40PukGtScKeM/5vpd85az6lcHCXJLe4d72/R0xEnTlL5OR+h4v
zANMRf9J2kR6aoXxwL/CqgBw1A7mIz9ad0W5CCbDVcjvltXb/BsJBC3iIMOpwCgX
ExM+TJCJU4DmON2rp2r4GuN7dm+xYiOvfUbstaXO1X3Pqv00rOaGTQk1tvSIY1Ng
0at4StbuR/mwr+NauIolU7rQzOA0ZS3cSe/EyaTeiFnP2wmpfiKcewLmqYd9bsMF
lDpSlyF8u118M9aPwyVPsBcD+7c5hE72c8RQYXIfxGSpC8/DAbEhV6smTmdZoW/N
p8Wevj4lWFeXZqSMQ26GqNKM7qo1qiInd5PRYNtxyQ74tnDKsPJD4SaXXsWdFT4a
wHh2eGY5HrXyBAZUxohOaWfITt478d1fPgKpqTCUJsiX0cCZaR7rUNamgRZHYNTJ
eq8VVjmhYoNrnaej7tNsl77o8dSTcPTeyHJnwjKU4b3nobTsjvMiKEiBfvqzdFEg
yKQO02/hCIScgqZXd4QTE8k16NlUoNA7qB8s04ILQYzdZpxrNoQcdI2Y7jopqCAg
iOEuFAtV1vGZD4l3h7C5JjlyEJETmNPPabdFjAMtAhTom/w+7e4sTWi+sUEUDUF1
62C+ULuW2mN3+0Xs9kOXd6N8vg2YO77frcZlhXGMvUOPgwuT7N1zmDEdQ4rRHCgF
TOqmyTxJwubxvuFSHT2xZjzqkoZ5wP2udt9wRN38d6ELy5ZgCeX7FTDVUskt/pm2
ECWMsnUrgW8xOAqEr/AcbfHXVRAAhYqrbho1CHPisbRtcq+PPPY4JL+fiK33Wrfx
oog45g6Spt/+XC4aQw863YOnpLpkjevx8uMne4YZ16gsBF3aW6ilUuvghjdD5ji7
Pbp3fa8o0SnCLRUbNrxdmgiLUr4x1NsrjgnOkVjoBIF05o9HtxDlFE3vDxC2J0+I
gTt72rdREQDDWXIdo9qsuhFJfywnZoDwvzmzI7c7NhcNTs7yjeCAZdvtArxkPThT
8NuTFrjXNf2Z2oH61UVoUMRFSTUDCDK+30ohRnqtEZGKJuQnJdHMrBbziY2t1l9v
2cWGBxi89eiTywECE6cRMf/vT0iBJEzjzdZusz4NSTSq6pGRUMSFqWBPFoTBkldT
bdCy6RPuXXhLfcA28CjReZbtty9Q9zNRRJkHfs7/DgZ4m7Q8b5QeJT7N13RTycbE
lyUOEcg9FqR0qD1KToxGGo01IhpXAA0TKdKTURlopCkVV+BQ+U+CsxG/bWeMADBJ
W8Dq6IKemY/sxCGhWgaOZp84ubCbSmvYZHc5nxOcu+/Z3bBbnJLrN4cKM3G+nqx5
J4ViDd6ZCsQE6/f+ImffuRmQaBH+scNbOaIogSlzXaMOmy7vEE1rZxsRkxEETkYU
r8MzI5uq9inohRER0x7PHzaGajh2b6cGUk7Uml8ZTOmGLXab47OuhVsprLqAd9ac
E/zk1H0KhqPGLDQS2oz9VaXuaDyvhUY3snC7XYcPM8bJJcvYRadpAI/PxTc8KJhi
rDLmzXmHW8H62zWj6aIUbQFKiXOTKbynRokFNBDDxmjRDX4SqsinEcwKgJLBCiUO
cg6kpzBb7H0yU7pUO6O2NJxcsVkC3/blSrcwXy/RWYrZlg+cr0mVhMNc0GH9XY+x
14IuxfK/Y50m0CfXGkByHIJ86/hlb8JJw6Xf1q2KyCvUzGDqbkhKcfyt7J+ORwha
G77JNFGev26yCsirW0qxSW8Ks0DAmxSatn1K4lIhIQhOGNZrB20UbbnBVa3e7xb6
/Txcdpemh684PC9XWwtw1Lb4MP3s317CzMefG8Qmy/SUxlP7AZ461sg9C6EH/8LY
y0iVE8USFWDjuHIiTKIyemQ5gV5A5cTDDlN868lrj0dmnA18irYrmoU996cMWItf
lFt88xaAYwNS3FH7wxUBA/8gFjU8yXq/oxI2CcDHeR09MndxY9oRM2bHBp5k494B
4RpNoFrs1Z53A+HVq88sQKOC8ztovd78rSkv5MAysMrAZPT0IbPzTcX1Y3PcJ0E9
vrKIGFUKh3X9Z3RfYx3iCg+bw41/EMoEjmvlcRvx32ky4rX8AcpZTc834ferweub
TrhIrxPhmSUO3iyJRkI391jdxnX4WyICOcFBwK+nsQLuak/xKEaQQEt92tRdzoEL
QY4n0AiuZX+2fItpl0ZZif4YbCed6nAE9Erg+TrUBWUfwRzc3fkIntSvO+O4XC5h
JjlIA5tGunuqq77TIl1vs2nySeQC9RcVtTUSgnFBIMsG9XQkuoMEg+FikXX8U/bg
/zz/0Z/Vzo6k11VGxZpNi79XxK8n1+buiQ83dpse2OdTplXKUE5kPoJ44OokiRz1
EwjR3S5hZExk7oYhEAEove54Yw7saWa9G9svn7dm12LcJgB76dybZcMdBLbEd1G1
trCWEDxj33OK25IcpkkP9+l3fX9T5Rjb/NgMsazlk6TMIzO8rdt87gB16kE6Cn/t
CrjGXFiBKj0gVsBFB/f6AToFkY4Y8sjyLmxSmUnH6eKpxMY9s1YzJaXdtTm+Z60T
NciY2HoyVYhbz4eMq0f62jXeZpm5EnazqGeqwpipH8Hjv2DkLvypH+XNcXCBLZUw
+Fa1wUi8K2bBCGddL8Qki3bNdmSNm3VC6W66PdwjbCfanxMg2XHZPhBgTXuuEWgd
2cOMbo8g6Fp7TYTwF8ESQQ9IxE42w5blTG1qnjHN6j2te/AUzkMGmXowCaenR7dA
nUfM8Ngs3/WEEoLvwRQ1XuH+NsaSsuf/FDkV07c5mWnYPlm16gZnPjUO7RIT/o9P
XtOOz7vYpuFSBjS0Ptd7ne15lsbGUSCCOMLbsDZfwwn9Tat+R10uJbDCdLOCga5V
WUm5v6m/JCABkXYuQp/oCMJG5kjMM2jT/+rKsfiac8vCoCu1/KmRA4YOKY30lTlX
GdmghQPqlA08POeNK0u9val2E4c2m2I8XXDAIEtJGCGcRqkqfGe2YkztUWZvrWHh
JXkyE1tDsZxm6rLAsujV5rSJbSauycFoF8UCs4D1etKXc0u6tK4L4qkWQk+HZRDd
8f7Bk6FjH++yBvcEyBpLPnhwwWH6cQYeJDIx8rBu/2Lc6c0ZHKEvVPikCOeDh1PB
tBMlDmfgW+0TiiRS6+3OOp1r+9oYKMIAH9cHF3FkPmxoh4VrSUuxSg7bduM2Q3Gb
LfpU5ge/dh+RH/EOw3BsUsVpxwFa+vsXHDyg38U/+ESQxl4+9v0kQNr3V24zUM8P
FxmSACiHmehch+gXmiH/L5AVBqfkWyCFQHZkvDFUnuz9ZnHB/DEEoi3M/Z5bJJHq
7e99p5UTj9bVLVZx5FcwJUOKkHP7Wz/U7WF41fQCyYKpr8n5LZY95WfdgJRo5GfR
18UPmhC2euueLOKYxl33mW/WwRV21c8w9KlCRXZzebUkwBaiDUwqNzKqnBVnyHWZ
BJXj254POpzTP7S7857Fj0PmGQM66cAAkWRAi1OmonTEdhe+UqzknEp9mrfFSIXn
u0Ghftshn2gDy9qyUnP6aJWLcjywwJhpt0iwOkqiYI3u33/jjIJo/bn6Tey5uPGD
79Vv6lZrr+YYYXlIyxicYwC8baqQBIAEG9EzYtz4aB1iieqdRqb5pRjTUIUFoiTV
R/oNfYgrat9txQON/0Jj5UX/pb2DosityQ+oWkdArbAUYMOF83G5SEnQdK/CpoaG
FIrHZXIzhhu1hYZOSJEz65D1R5/Jtb+gLMAalPMMcBMS/uhs1OubR4DPkcFenKXO
1UwBvxfWz4Cse6nyz30HRU/Cp/mh9/ePSpenbcH5P5AvYxHG7/CKNgrxz/42YsOH
+My234wwagTA+OQG/kK16Wpbhp8ariroSIZ2kEsJ8jJ5LU0s6OC8S9qNKoovihXg
V3l7kKXIqHptMXeaTmPbNnY6dY7ZArmfrnW/dkr8wgqomH5hnEgrLbLtPQgDG77+
iB8TfBj+lb9YVVJZn2NpwXMJ31v9OrG52wchu7LuwhjXSnBsx34UDCN1cPhSFdmu
IfJpuSvGtHO8WQlaB0mdhfvAVq++C60+Wp4nOBayvSPGNnf2mbS1E73/1cjYxPLv
xxZuSd8D3gDZKu+AxGv0zBnDmKWtJAVRTtSV7ShBSfs7zUP4IRK3nDex6k3kBJH4
fxG4uxnWxpVKKxXIKcw6pCOTVgzaysGRqw+yt/ZMlHcCnruldfBtKoDp+lk/qDl/
CEgWN4i7rthWfeGhaErEcUqzRkxMQvIgaboMc2VPwVxJeDwbiCQ26J7bN8QW34pe
6tqBobdBh8GRYTJFKZXr6a7zpdNT/qjZUK6WkzhbFNM+phg2YA0P0jlRlhxpH7hi
Tj4whyi5X/fmAC//9/JNWyztCDiFG9fgwMIOKhKW+hzLJJ4Q4EBcb5Mqz7rhWVTY
w3aK/RCeNKMXG4XV2lf7kRFubh/1ftJwMtef3f5tEiRKU3yyvQ04EEXVxww7ZJoW
8Knh+oLU4BcFr6sHCotdJo9K2CtFEW6wDU0NQtvunq/H3yIIyvRqhh/FprNTnSh5
UhRVr51e+WKnkt097eK/qIqUf7OMTRZsZ9+6vYPIyI0C5ynO7X449t3+V4OG5sXW
C4SNufepW4kuS7GQ95vvqVbEWDmxaxigCOc4nWkcIQ9l/Lwrn5iRmkBQIkCbxz1L
O5FLZxLQgnQ5zSNSXCTHt7hdVKhRCtsbHY7myFjBj1mKYzPv+OvP/jvE/28mDn9c
024ClhM6C0vqClSBgimtktqMAdWWdL+ztSIm4Xf/b64g3n1L/z5EAG+jwA/GQr4b
qGw/wZGtQ/9J4pR6RH0J5wFtIrIdBNEgVPO27n+pUffq8WTHubemxiy9t2lNFkG1
geeKIw3qNHjYjScJzRjs6GPUCb3lEXx3TSnTMG2VhJqkXdA9MSI1xWxOuDpemvyr
Uk4rlPC0tcgq8aRjh3bvju9cEFjOe20LTA0Nhn/uwGYWlsvgY4jT9m7NcYvCYPe0
WmjIBZREvhE0PMS85dvIEpCd76AL5IVwZLDxCFA8HuZkKAISEp1XEwHMRGcKXXiM
YYQXSjLbmw+AXKNFr+kSgOqj+Z0dFmt7e3+fnUgv5UE5oxt6WSwGx/5PkWfhhjYW
IBecGjlkPFUcqyml5pIwoc6uG+jdWquR9rmSoPzKnQoOB9pfwH1dxoQMyvESAsvJ
b+ziZMYcvqSMO4OX0HBgLklGynaroMqEo/tmMuEhR7x3AyWJKR/dXfaB/coXMlR6
x7ToHTSHaz0fJ+4xhPIJFSrdRms+PATH3eQiZUrvS5QEm5ThN34ScyxBMMYTOMth
SBeeVJTXxqkcSIYuohf3goz4WScAywp0iTs7SZKdTBIdl9Z67IFDa2MXbfPLTW3A
qOU0HD/ifd89Yy3TLzMHfHMAoHM4r6LbKVB5Y7Ci4R/jhh7OmRzUgio67TlkPdTr
ix+61RIvVBuSiMBW+z5Cz6ePsqwQCXwIGWdQkIYTEq+fzC+lYiM8q4025Z1R8bq9
3SPPs0cbz7FkE+m4+SLOF8Vg0vQHUK7fUA3PKRTJjekNjOgaAutNVyeEaIgsnY5p
5nVwEGZWdTO0ivHCHtFXYxODw3ZaNUnUSs1wf8VQj/mk/ngS9MXOB4D2IR+9HFqi
/Iqtjw983h6IfIAdTEy4w2qkhqlB/8yV3yK9sZ3hJ+WlK5PYIdMbqqnQM7vTxuxm
7wMIAy8IhsFQk4cmvA6BK/61CaLWDV1ZT+7bBmOExYkNDBIH2YdK+oONXcE64zlA
Zqo1AIjc9j8DyCXtdxlnmVCYGKFijSCt/1GszWCzkq4fbs4G+mEocK5qV99Kekk4
av9e43QYYPCN12ozFa5FiiZwf2+AA3epx1SLJe8WHhiG9MKJKcMJr+vBx/BBe0z2
yaVaZXUy2NZXhSS+ITpCL518Em8p/poYtYuV+mGu4degfNajUY/O7l16Jm0UN4F6
fc0o9w0CuT9R7b6VkMXWHKx4JLtHP0uojG+QAvhjSj+97MOb3pH3z/2DyoAJmwhD
YUCNzi7qzZkj86NNuWLPmdfPsP1rnoqYDZMZXFqlGKVETeIf6BDuUa+Zjd0Y68KE
SwUpbvN2dSCjpSfwZathuDh1MwUDfKj0E9bt1d71LwwJeq12I1qZ6RfPYnKLN6xS
gBUNtAjNQOAzgoH7sG0E0goDinc9CQmmSGHzjEdhwDtC3WrXsrEz5d/UXdq6WDrB
d8DLml/CY+LnIzx8KvN+Afda8KvCrc4LAealVq6BWSESlrlygbl+4EVJY9qoYYWB
GA4fXeFhnHG+9FeD3GlxSKnglbKyxXxUPYdeVXP54OnbXzxTu9E0tH/gpZGDqTh1
5+jlfEY35QCeOM2eU7R8S/mpNS6jb0i/q3palVzeisS4724nLRkt3mnx0hAhb5l/
i+9D8tk/QSJ5xL0C/P08nQK5fy8dOzEFfLNV5rlaapgZIgQm4dsh9Jbu12kh58Ft
Dya022Uu91mknefU52ZFxF+kBnPQIEnTc+daCuhOQzgqt+t7fNqOiv9cNFFeH3cb
HH3Nj+QTvsiievaLaXRSzVn+LZdFNGH1g1QFQJe/VBhEy09gYKh2xMiIvtMpih7a
dRfKdL29rKudtugppbEcfX36O3whK9ZqTvNr3nX80xWht7ovqeSMn1jL0iUpd60S
uVvCGSsPKtrIp1DqMFJ7KUQ9g8hqCcOQWTw4B+nXhxWxffzI08ZqXeZpHor8ZnTs
odzi/NShcUDbp+QnMW0WsncA0WtSyMzABMBCG/m1WzrGjehfWY0MAPAvoOQYlqx0
dGnca6rnAz5qFTtdVbCRZDG/E/sreKRt/mv28OfrSuWu/Aw+UH52lhK0yZYXqDFM
izQF7oURAG0I7TQ9C/YfYuc7OAlEROsxJl0bgkUe8jXvAdPLwgR30cDC/EkiFaWy
Oj2B9GAJlXDWhORNltXVMSK3KEi6oor4pBhQcD1ocu+9TSdl6IHy9vGaGvBmbQ+Q
OksgPwXwvDReJrWyf2Jsj7+HR4uL9Q+NtWR43Hr5kLIJNerIv54dD1PJVx9LGE7v
Yulit9Rqj48CpH159HMuiNxP0ecsRQhBIlyYwxb6eiVkFeLa0vdoNhr8CA/cgEnO
O4SrrWO8tp7n16OylEK2F6Z4AIRfUahDtq4Z1tFUMHqvndpJuMGlBST6UscB9ZB2
2mwobgif6DdXm6cbY+MVmO1Y5+9cI9d14yKkVB+ph8e2S7Ho90BWZtXfd6oJ+Kct
5101SMep51q8HpkGDuqjQDZpjDmGRv3WXvu7EsdqpRLYGstUnew4p+f5CAWI4kCT
vImS/mTawgOKJpMRzjYuX5DKHbLP3GKafuoLAwVKir7e62b7udSM1AYWcWMbbaaz
JoMaepHaPzyctnfKk+10XxG0BgSWlgfcmKYf+2TFDirZYUE3CAzwBEw7cseMgDZo
Bd3pjTzsnxAM0LI7szSHw3UtFQkugVsxkvKHhoYSBFeml8EHs9IFYqFc3dcizEgP
zb1Fs3EvEWQi9wnUy66SXqcaUoHtYGqv9DG6BHqUAE56CQwNRZ6DunFMDpl3A4ZN
TBYr7CCNXuLt9L9A91uYxaK/fkoOIQi1EEb3p3ekYM7i23AvPDK/CMKsGDILbUd9
l1bUJb5eWnV57H1HwjZ5Nji+Ol8D3ce+o9F8B2nsD78KcluVByaR9ME6IIzicWEm
NeO3EQmA0SWX6Ud/dSrn0Et5j+SRTjxwEfQYNyg5OyjXpumNEuAGsBv8l5ZkPh1A
tX6CaBp9C2hbl5C/rEiTCya276lHGj9JEo93Jn2lv9BdF8mK6RFiqIx6jtWIZyQR
EHh8oGokZ9ojHtkS09eKerAs6tnwLTCWGU3O6PbzSoG/cZgtwv4pQA0Ert+zGqEj
3HncRbPECsf9dqpPq/9Y2f+xhl5+CGPznZ5VTRtMfK7HLaCOuYDvYYJP17pSxIgv
R8TXOmn9/PljAUVLsU92djMG0Ae0iRaUJcfhIPqOigdLzTEXyO9QQ6uuskIWKS+a
QaF60FFhITaGUPgFplltGbQJDo3uzxFtNgHXNEnGlz8kjbBOLjFWdu6rjiZxd4MK
oN8vYoOHmWsNDro0hOgQxPrJyzUPgu/5xwLZYtOm+vEkDktgOzYFAnIP7JsDzhEw
h9hH1RNQ9WoC8ZyTUdsOAVzWFouLGB6evoAro3wMxptbX609g2z9qY8CXamFa/qr
r3x7GEkopFa2UWdM1YHXofniPQtnZvi+x/D1paaSb1I5AN03zV22zb1UJSpr/tYv
/Y3N2XOflJOhPRx44rytpZL2xX9tEzn3/L0gQt+talHNQruZWREzcfS0djpafApr
b4LrxbOQUkKmuyFQaRUXOo7DiYoC65FHHxcMCijbrlymuBd2MGmrCWMrY5dgHPCO
xtTjA1lngRnk1o88HdhqLM9nbx97c+3/CmuVDDktc+sRB/luY1THhYkSL/L1IUSp
eevQDfDwRMsv/Mce4QScU4LeWEtEECDlLNpalNvEaIajJH9rrmCQLyr/D32DRvoX
SQlgqCF83yOLD03jF6be6QnUrjX0iYAlwyQfNRWUgbVnlxUBLfNrvllfn+4YLskp
fU3OmVsFKpskBgDexmwYSx6fC1P44ehdKgztCJ/60Uu8+Y+bjlJ+/cTOS9PG63r1
LpCFIqfQztzEGXVihktxU+cDMJ+praqyx8T9QoaiwSKhlHn5Ikv51VxYjQBArjsA
c6DWR6r8ho8dEoy3aGCr+sOUS06fg0bs1IeZJqCBrhw/3rCUxVCoOag/RDcpgp+D
liQqEQSnETpKZeYFeFtkvvjJJ0kSG8SsGZs246po3UTKYWIsieu+x/+WX89BPlej
IJPhg1zCQduAKH4x3WGkW1ATMFlZGxXXPr723n27vlgobgXTYKkMMsDIxRsuo4lO
nU3ZCe9PJn0KhG1zcadZ02tmRQJtT7402myh/d/3dGmRjmpppd3HWgk80w3fb/eS
b7Y1R8QCm1/BFAzxNAfrY8PM6752LDXOYh/W2DSH1Tlq4bx66VxiuJqthR1uOxZk
65qCmzncsWT5qSgYutWum9bZ6hKwhvbXaeDGEn6fwfqWkt/G9wPfISwL6NW85UBB
hrEEOaFrI6YNiDfJMcojgnOxRx45mgyh50mDD0Fyj0p71xcHDF62ZZzGCow14Vy+
/gcC9xSlYEwEb2JYqfJEfbhKVpEVPXQ5qWERCoV6Sj2O3HTw153c/IC7V5D+/xwx
yyWaWro9J7NQB/peMVO6oLOsOAD9TPBBxI818GtA3GClEunB+UzfPkz9/0JtITnN
z1+n5OuCmzBAH4LcUsYwI2B708+gC9cCWbVSiJC3iQExx37J4WrnbWCoxVZxpkN6
MMj0Z6Unm7IcKVHjO39+VxOQlj6PiMqOQBzgBS1BP0X991bG6BnPolbOy9Swj2au
N8/IiuY0tk6kTCUPbCrVcPIICctJA/rnx3GU7iT2dsm1NscjUIDYCczUnttt4d/t
4h6z0cVMuces1owRpbJ/JZY30H/uByXQt0u9Y2gfh2LL9GHtVgdeLvX125P+aCm/
CtPB2QYhKGT+/OQYHxPkaiuztoCO5MYXNqAq/WVPRuLDJoJdAnVoalxzLWFT2SHS
ti8/nkWgcRORKcZD6qziFfaI/2Q1zewsnM5xAalpWNkl8JgfQGzoYN6Ia/I2NvIa
r4Mwq6TMBdfX2QuEnZ/xuMKI7PEzJaaqdu631T0dQLT7NyOEyOiGxLXNtg3GXZWI
/TUhh2i7KyhFcwYC9fvda9sYXJG61uz21DKtQB9tgigqtWtRwqXsWZ29tLB+4B10
7Gp/xHnCjChkQn2U3h7L+jE3l9r/KZmY/WdpPwsEEEYdljxmR7PMBcUbb3b8RUB0
JLlZhDfpUV0HlqATMaLVq+W/BJnOLheRD6e52F6LI43c309+g/ykCRtDSlWK8R/Y
zQbciQcvXnSNr7FH2sVwCPxggUrHF2VB+z7TKsKfnRdsHcL6bsacmh6ziqUTuoiP
JeK0y2cTxDTu45yTUXw0LiP51BUq1HrJDNVTwYIjhgmfXiRROVCJ/o0W5e1kqMzt
jEmK0PNjXohryAB8I6I20d1Lr9aFkzwyNiBYrxv0O8IGcu8P8H27gT7dr0D/+mCn
A2ad8ucQm6onCM0XilxWYETiWrNg+zHlF21piWoFrcqk8/9nO1qzimDZI3gn2hTL
/aagabKZnOrsLW94w84bSHc0lhVk4qDwSPUZWlRHqtlk2CiG4pVnBVqS3dWAHYDM
uWw/pF9J1KfOtuu/qK4S7ZY84REV5Qa9Z9CulXq5dRZ0rW/qy9bFzPZo/HfAZude
YXDi694RyCGzNnTqfHmTcFUfATNlEpsf576vDX+PZy+m6L7FAfW9WsbeDYB9ICYi
GUxi7W5murtT1NwXv6xfbiuoh2/zt7ldH2HZz0LpGhPmRBhJ+pRdv6u4eiXGdVJy
VUhzq32xgZpkhDSRqAJLg2XmIfAN41V9GjGuhT14QN4dBkcNKoF18IkGQ0S8D7Vv
gH0twFEUMsRwqfJNNDWgCEv1jrllL8DdzAv4PPO41Sb2DBjyPzEaiAbqFSPmh5og
GtSLDgGyzbD3dIArLMEJDcTQjDQevLFVSh7WptdTPmjOLGUpIe3+MBsunz8a9M8L
J7k7onHeYs0FZH2wgLwHHlno22TCWxL+mhhOKXqCpFqjYbEW2+Cn1URRaUVAjbrf
lX0D5Lv87VMtXVOCacrILWSra1LiiFtFTx24A6mIQBv+Ma6icP2KdAkTsas6in/W
30b4odWOP1hl/43fhMdrAHt/Kd/c9tMI8ilRFJzYk6DkxA0mIiZ2MpsPGEzWJG5U
IOa0XbqztXp6BsIVpuDKFE3TxQiKruTxykfvvUGNgZTyd3O067Ys+nOoGGu6VfiY
r0OuScRbIAeiU4lYxvs2PRmBZEsxuNqRctjTYOubvZPUtQZWe0uG3JT3oqixeyKK
R6SujuisgdDuIACf3ZLAOdGuzDfbOIBHD7+PMMzRuKK5Vqp5LCDyhrQyLlrL1m2z
FZTLvTToe1FT5g63AjRVm834pHTE3NGUuu0wt/awz56V+UJoTG4lMMsWv6jyyC5d
vqdVoMm9yK83pO+mc/lwoiqqlDM/Wbsc1rCy7hVtzjhp0QlWSCzxdpawt521Rvdm
ajDASM9opL5NgkEOlQ7Zf/+4t01Msk5Z/d/lJ2+n/OnWHvXz/2iJ1NjvlxQIAjiR
xti49TP9YeBpJsycqx7cOtcgOsxqNpretSup9biZ7DO/C/fJGsjOcYFUerheevlF
6CM3n3pHELabPgjDVVmbho5fR0yN6AEhd1iLONaN/o/cDaA5ct9Ey/suB++aAVZE
l5e2SDYYQCP20T3wYFqXiq6wqj856Lap+RGAmFi2j3BXJTERQcMATbMYckN12l8/
+lLlEore3yAFlTycoyadKfgdEZEcBwzT1KIU/+KpGD4fXW7C1okitNxcoaM+kYQM
cVtFZyDU3McbJqAZFrKZy1Ok+8Ko/Ds4mSYqd/QVy3LGYGB8MXtG/paKx35CEMki
+YqSs5pn3tcrrF34VIWCXhcj798br2PTTP/DerO48+Bmj1QY8ySSSPy2iF7iDvZ2
MDrF44rucUfT93qsomrii74jCSZxRiaK51Xd9rxW43kf+sndqDv/Ryl2bxyt8QCL
IUGZOV8PTpYosc2H9/TM3PkPJCQNOTx73Ni4MiV6W9BsFJpXK8FGY9dwV8EiObyi
aVCVhLMYK6kNfLvvBMNeUMY0agzxjx3oOHcFvkf87HywCjd4YfwvhAO6a87pm+FA
+44ZulXMHBE7YwAyIdGHi2z/nqKdFJk9skYtc+Eajxj0QXrmRvCqeu72qNq0arGi
PiCv8p6wyt4zru1bYQmZnwx1NzFAhc+Ciaj0PoDoSFM+olSsau22AS36axHkXs7v
ekRbLkzeUpwEg9jEh7Nxsy+zstG1+w/ovS0h53sDh5LwEN9qaeGFoU/Ijx+QsT99
jqP9eu8mSFY1/E/taDo8mW08cv57oAF89UIQ5UmKIu8RG7FAVSnKOpWAMB44dy5U
VDhAOGgS36U9kYOJEq6YckqfiknE6yIuPgy9hJwuFF51tL9RoLGoE/tQEZF2Bh6O
qgo1OidvkP75zINmui35E785w/9tBMYJcXlCFpzZiojCnj+xA0BVAr0g5n8wcUVL
ocNpdb91YZB2GA2FZfYKye74laXx61pdc8fdx9CjAI4PGwpmRifPW0WVkqFniadE
nxns+dE+Bt/1D+WPBMpeLHeQR5Dun8Fiy0fYrusDORKaO1kaIaLxWWLItSS/qKVg
Qw5//aFBAYtwG5w44xQVLvXfN1/ntVzxDi1tjRWi/Y9eLzUeFTHYqurEVG/zEZd4
CiNv/UBNnnheBr0ddhn5enGzjyC9WAsg1RErHL84KRGT1xyEa6hTsAcLl4uQA2WZ
Vj3M/q1/MXqg+CIbNGti3gjgQ61pjZ37Uhk6Ic5sP56MZ8U+8Ucz7ppUOOh0l6Sc
3IjZZZj72D14U8cemDwislPaC1/3hZtu8xPehXb8zAzoXXMLWhM1pm2z7WE0U83N
M4UcMRvAsvxLh1AxWFoCnc8uj2fzdBvjSAM8JIc+041VOgHf/xh3+aG3SjweBx0l
M6Z9tKZKrZsRXkZmkvFyypxBIKTn3Vj6E4ATVKmKDLVsCP/RNEGnhEWiF/7hJmEk
84yP1FUY22yevh4m9PsGDQzVti83hvvs6w3V6ZXXhHGn29MmAid56UbE7+2/0Vlv
dpzvpYq+0fLq1OXwR0dRdO0qxkJVhbgQKot/AnqVb/7vHmGMXWXJxg8RmYDtF/Lu
mHFQ4ZvhqW0gpunsdTRpHDjI7q1MCsypAXNaYN0O4SqRXlhw6nTInSWshcV3DrjY
+cTVipaDaT3kryl2MzSCreezSnEpw7EOsnT8jxsUIIz0pHTzlTKbSSp6PuZ7tAc2
DxwTAOmGVkH+P2VFZe6u3q7NEz5M3fyEbTS3y5T+AVI7JtyLf1eZdDT4dM4GLs7V
qOZNh1h3kLi8lHSZ9KVcJdyG2FYdfSkuO/4+91VeXB6Z+THQvR0bolS8RtRHZyKA
6a1h9t2JMPzpt1UK9aEGYLi9OHX+322Mi5gdamv4JR4bCvpn/HsPpKYC2+pMFi2I
jp+Ie4O5ZIqr9TjIPJgzHr0l/OKRQkOKiA6KYPenQBtwBaJ9FOPUEuLRZav2ICBs
pQA+S1c3Ir78544bf2wjxVHuXP3JVrNU38k9UCUMEYLiiaKtLB9xlMrL0LT/XAyi
kR25wAS9G2Stp66eLQypv3YegOjRzhrI8wjMee0QPlNVhii4bd0HW/0SLVf9FSXm
7vfbQIz8eugE0BTqthQKxcCionP1Bgw/6XGpr7HcI0cqYOMsQGGkyVjr+b9f1r0J
UbUsmfGb1zHeeVIPyXC3p0vUArkU7iNf40p2tmAl83cof/K05sc13p4qSTFtV2dn
lZBrs47RkiEmXxFCptuPICUWoXNcMxZ87ZVXazEij3PYaD32/o9uVJyp4SB9lvjM
gUR2I5Ko8aZ6F/tMhnfjgsApf+BGelse5RjURRn0nXnAEaF5mvVeXI4120Ekz7Cm
7yqWpX306orbxpdIbit1jOYWWggDOBDLYyjpN78lOkcssELXyOXVhFc1T/JIyvKw
w3ArvdlvkLYiM4D2GtzUMiS5BOEiCPjVnmlyYhbw97n7tAleuE5/rzr5yKOJtztz
l0LNSLBPew8ZCNBeA36ZKbTBl7wHKtYmhwJShZfsX5swc1UyP4voHjp4v1N2Z1Qo
n7ix14f2Kdd2eb0M4LQJyzLW0ix1GBwHKhywXHvRX2njmD9CXLK+QWYDTO3Il2js
LkedIUYfY2PogAAwNGspe+5BCvonk57hfJb6W953qC33K/PXPKb4prQYuh4bBJk5
1s+33F58OpHw4S3W6O0Gzmc9hpX4hkHS2MysCgtmucDP33EeDg7BFw39INMGICJi
7tLLJaBNNWP34E8Y0qQtCqifJ9Fqhd5ULJrI0YJAS3yIexd5e0hLoKlIlnMqv7zK
Kd19JyKZFnLGfMwNKHTuNbbAX+Dug7KLKaWltWf6JULK0Kl/a6XYmQQRfqGSGpji
6vubYuSVZdK3Pgn5wX9hXaRQ45DB9HeLgA+xqVTZR9/x0CwmX2eXJEp+ZLF6ytgq
QwD5s1yFULFmHZJ8Omeqrf935tBvp0KMD8/DHuIYgJEUr98HmuTi93X09hYWpZPL
PAWOk+QQRjXIMXDCA/lz/QW2JzBWsCzz/1CkHubjumXktJI+0Uzumpnovvsp9sMW
bqPio77CiHfJm4hLNq/u11T/kF93AIR8R0+GPBIaQnemsk+6+pDS4e9XlKR+VDVs
v7kzYKm5LEXoHYYosajyJ99xfd56smZ0e+7sX205wH5ELb30EOZBqAlwRPolwAh4
iGLdQbWpSceo9eODRje0Q5kSD/btUrMJtAV7BOxEAYBkCUPlLizX/R7J8I9FnLum
zj9qRhzQJtBfBwsroA+igz+TJSE6ZClSQ5qAjKA1/+8wj8Cn2JsoIpFKdYvpeFyf
UsIZWB/H9hsneN4FzilM4m1OOKllCfLKCqhuW+s2bBoVfxOwPx+g1+8PQfjgp+f1
aDQQN8E9gXScMsDhx29H0SDwe7M5syxKaOi4Y/qchpF6kLJjvVrrO/oXZcNatdlB
Y7SzbyhWxV/lrUcU+eI2QwvV4gDMHDQ6B/8/hmMeIlvC3A1b3y2PeACw4Z65nppf
i85v4GPSsnDgq1u8eBdmqnjunc9Rm0UBxuvJCtIrVSAqYZlMnzMS40Ltq4RDx+Av
GItmDby4v4KpDSKu8qUrBAJkgPcLnYDY5buRbvbenHTYFDCNE2n5OFSua16J/225
c+iIJOvu12Bk0Abf1fwIRzLFH60Ka87Jp7VkA6DMM5U63pcQbhnpDVgHpgoEvmGF
s3skELS1qLoIq1d8bGOLaZBmRVirbjyWWTh3mlmiJDhepDn75VZi8IbUFs1njRfN
L8RuHLQEoo00omJjGgBUv9QZk/j0HgCKW5soDvtMuzgNMC2o4Tjk6g/Sog7IT7XM
hksi5Un6WTSrdSYljXCSwxLTLQ4bsrvA1XJCKQb9hHCJ0mx/BzL1RZN+Ulj850xK
Lq114riS9ukxCAe+u89/NnG+VDvz2BcRi8ChIH8qlTQgazCVWf9rSvZQ5nu610Sr
w4Ff+Uap6iLsl1rzOQ6J/wPU8k46kMmLBe9CqlFZqzd4AaTTmsMpgjj27B1a3xm2
l5vIeMY0tEm20y7VIv+Gdd2YJtM6bzSabEW7pLM7k5hqoh8Dm/VKT2q2a3dUmnTJ
37TQx+jHblig3kVemrPkhKRmH2MHjFsayvKgiTKFhYqKP8mTVfi4tLSDsuLyHQql
n1wqMav7DnLdGxiGFkM+fug1AhrbKZ3DKa3tOsoRcaNepmNdpkkB4fu4XTIr8DVD
/GT2kK3lfSFngHtjUqOX3CGBLB7mfPHoxssPOdoSqXvLahSUkSywkAtgJFydVExL
iyXs7kislsz2y4LpC60y6YWIgPAhGSF9eDjtEnToqxVxKnTSLn/HX4joDHRUBSxU
8qOAUPJh1mYHVwW39t2WEKEParnblR68uOuXzY3AVx2YyWdGkX4y5MkRl/rU+H5c
rWC0LxS0TYFiKpE1bRgBBv+080OGij27H/GIYPIMW748vEaCqbitR9TSsS9B0gmY
qp6dbn2gxOKMP602+SI7l4dRs3s/Biel9DfDMLMYDktwRzfzFiB1559ScMWBDkOL
T6tHOj9q5XM/s7OEMgefH519lTzpAZ95j+dqWCNp2bGtydHWj8BG4GFdSX4DF8z3
2AmMEMr/Agk2n9tyNDaIc69oXxlRNLfy3DmkiPB+RaZePZkA0HB5lAdvZDFPcH0u
2KaWEzgzav6lSo0W3MITrHObzS217/zJLG2wSCdaSBFalVWVWOAsRU0Xbt5RhVN1
hjee00BssRqGw8PUdJW46NDLc0HxeQTMnB65lstyPX6NwEAX7KHo/jX3UNbeoDpQ
ysCdZKPtTIYfkiGBGmmfpVR4VJV/Pn1pP6jy9oA70h5iIX3+1Obf//0szxzK0reV
JtXzrkYtgzerwR6yaXTN+Fmz6SpuGoz8KMzMtxIJoWtlMLcV73XeMwL9zSiAT6JI
G3Z9XQHohz6i2fR/rzpEr7aCsFPAqqd+WzUqn3fk3nmso6Z5+2b53+8iugyarDBd
Wtqjb6P+yNJ75Otud0bv4DO4ZcAiaL4MasTzQo9gx1yPVmLabdf3kcwMORDLeF2d
Fbu9RvLFQ1sg4KollZHXuIiKvA9UeqZzZbFNXU//HWmqb3q0i0LIi7EjaVCx4qqv
ylqjmtBePdnKXD2WgBUJ7ACPNmvLcLA+Kvk+V1jJKv6Kf+S3zkgSzzA/EWOFx7IE
KwZUDmin39RaxaVu+b/hCpg/+MnH62fkv+HCbzDpyRKj7Kk9NdkX9mIELFPRGkpB
xt/Rg+zAlWKe8X3MH8cULPHq765w2OYgsKV8D9KeJFs9M9QP5Ur7TbcqcR6GrcuN
a5Y35o+uCYo2ablFQ5/vDQ08GKAQaTo6c0ccAZzj8ZvnnLZmcRdAHYqLvZ1e2RJ7
D2hxzfP701ZqNXZpUROop4LX5/Qp/cajYQLPC32C7PdNUsZCO5nKjhEwiND95v5C
H3GPei4fUwLzxgk3sw6EsGjfkOVGGNfeu/DpPAvXvZa6N7Kn/pyYrYCvaImK5DFd
GSJA9nV2Kb2KovBk5LWr6Vb9qEhSQ5h1M0D21xuUhqDbyq744F5JqkIEO2/uc+hY
GCRZ2Zka8vWqYdmLvNvLO2gFn6D2bx5kJXjCAjKrlQxzKEVMxQvd83SCBXLUNgDS
ufbNapjg2UzsU5/Y0ErNpmHDQcfduTeQmBmWIdTy4PPc6rkdZGwOTEiiAo5j1Yve
Chu54bvx+EW8STn7BZjJYpZLMVv7J87Fhwi5VQxItcsAo+KvIdpnh1uR3u8trRuH
M2d9wPkbMSoj1CM0c/EPJbU56RRCGlVVZj3TNkeFEfFGctNcJZAxszRWTvyqjMR4
CndQ4eOMui0MVJqOSLyGfATvNZvcGEFMFFGYQM8qqIaRWrQEeatQv8Do6AaDEFhY
Qfkhixg/e1iFHqplKtbgh2gEP5bdIaHxSvkAsEAvBg3wVKQLlfN6hNkbpmAQwoM4
DOXL87D0vOOuEoeGNNlxZzDWHbYD1or6ynNSYgZJ5+INeiQwHYG+GYgcVJbzLKg4
xbzc7ecmGGHxvUwRkz/u/F3OhcJlXiupcOiGhvGQPdXvhIzDfGNC9pZqNBPJ84YF
LH/0RZkFqpwZYwWVdeVYxRgfuyiZX/WpxKYTHFW51PyVKd69MNveC5S4SzqgRWHy
RYhwiUIMxPfg84/+Ath9dI6j/TenjYIcuRBiOK5YBis7u7FIQq/snsUnGspZBWVd
6ch9qsk2VXcgWfzW2ju+A4elxp5VKkDC+W5Edk0912BJrLTQkEpbys4RRyMspAVI
oiiTBln35j+MWkzH73X+tXA9NqDyyV0BIYN5Gc6g7MOJ4sdG5qsO0j/6xYvBBk+Q
iUwnBXORV9qlFUpjEo0Lez9C5MSfEa0F54wOHA+fFlzeQo3SOl4ZjY7KUynge1o2
844tejds+lJ2ngXNpkcWHMtsQ1kClhFarjM+oMRgeijtPdHA3wMluYuGC6HvsNXp
0KbSScWkq0lW6+0Gw70SUy9+cDzwHZURmCBny8UK6URXHwzi699Dq1AH+r5BJR/d
XDNs7H+R9o9egsb2jqSw5HA3PQeiDTTMxGGrvyl1u6HsU9qsk6BVQky8peOBx1Oc
2CRwyNvFtlW34UZ7L1fCu/S/8PAQ3bYyvIn4cB+hUTOkdmH1KJeEZTxxLc7XjjMz
qL1iLOZBd8Jt6eDkljQr5m3pcEGLM4uRA0ASk2q0JXmPASyaqxlfBrmfSNv7+XCp
REKYNXcZoJtCVGJNDaRRBbZ5hMY+jJRpWBq34SH4Ow6y7BCrw2vFXd6xLTmURsV4
WzPTRMPUyF1n2j8jNTQHsiz2PrXzebq+9lgV7yI5rUhJQvrJGQdlP4JeiRuwxjz0
Yuj4CVq+nbg3DVp76MDt7NxFqEDrTKZ4UBEkeBTjDGMbdqtYomPO4XVosSRSzugG
2mwcwH34nP9KRHXz3YuwLyK3TwsUJB4OD2Y6glatcIEmtZYKZxf7NK4z09HkPcRc
d/N+vUoB2dzJJCt42+/Clpr9tIbWEK+EIK1hNB0fioib4Z4obJ+ORTzCoIv5iRiD
PCziUjC4FYPdyEWNENzbHql/83eo9fUs+ihZWdQyIo7c1mtqNHasQnof6yA9Ohr8
cIT8QzqE5vRSzzZS9x0JtXtwj7LHvhLtqfEXSday+c/pGouRgmvTEQQkdFIHTCSp
q6WUaABb/6d5+TeWYQBWAy1Nfxfn5Hv+CL4ixaCYa6Dlt5pIpkL9mdKFOMcXT3JJ
IYk4o8TLo3B86+ANs+D+5yXaIfWfcdoy36vvvWwMj6YycIBCH9VOYC9wNbzUChso
Cp4AvQ9Bh7plZz+1Hp8shlpaVg2Bz4/+85aTyoaw3vc29TEPTuHB7Q5lpZIN7Kei
oVOpjDmsFfoyQAJ6D71G2yOZ6u0P/b6dPBgMmSv6ntSYxDZMZRjQ2aj5DUqJKLEv
t6EmZtWKdPbF0zWU5ClOX1K2FTidhBVh2WYZlair2kRTjhX62ffNp0Py9qU9DqOP
vrhOU20bIt/XM4JAs9bEe37/x1RpqjYUj77ELpeyTk8tUlWZyTrjwfqXz83brgYU
bRfRfUjeKHwTL/p9/CM/pJ0j6UfypLUTbnujsuvhMdPfnYAtW0/2Xz0Ymi90yC/s
JPvkrMVFSAyzlyer6x+27i4UFTjP1f0GIT+I/9dCscH8MmdSNSYXN8SoA6AnC9GW
vSXRLddYVz4MLdl97yKBC25X2iEiUyAUuUIb1mTZjrnkQkRW7RZWZJRJYaZuz9y7
7FZlNxaN6dolNnZFvX2NdZeRXuYecjNUCwrFHlbCbpxUbYwPw/tuyt7cXHpPL5IC
rm+OUulceY8OrQ/YAxyJ/B56daVZIo0qBOQohodxlzsnOOTULfFN+FtZainjM0oo
DBr3V8fPkt9OOg0ira38wOJCO25k+KuCGN103oopuAlALprwGA58+3g3gli2abrH
m7vJtCyC4QoEnPjNLrCeVzdkbT1TOeg6AsfKy2/MQBqOPQE9O9OPcxvw1pjDKPX7
v1AJAu4Fo/C6tMNj8zNe3k3OHhaqhXFeFg99MifD4rOuf8FptG1UFbk9xemdiHY1
mDaZMcCk2nwsVXEfNm5KTXbe+99hQP6s3q4/8WOteZ+a/RFZxkLxBYBo+vkQs8Mk
S0DxwTfTC2gKUbElNL7PHVA/yfHHsQhsLYng+wXjjIfzfJVA7LiFp7NH34dR0ED/
10R03+LlFjaCU3gr1waH5YZWCBuPRIGfpa85UCLAbIL8ernjSUllqeUeF0HH9kYX
u7wtpdCa8+J3fV07TlfgjbIiYC8YQqzZeObXf5P01+imUxWqFm9i8J+z3mS9d9FF
T0Ljz04UHf+qFCpvR+25vYQHUYI958FOT2XpwI5cHax6TTVrwiSKi3Ct61AJRQ5a
NDoZFhKQ++O4yMDeBRY6Nepwj9v8ZjvHa/QI1GVum5QUltg/jC4b/xFSekOolhli
1rI5wd+nry8gC6SPQIMqzy1gePPWO99OIOQDHCT+VjrCgNxI1aDdOJAGEx1rjLXk
Y8MMkOA6fvyeEykUXTd4LMjnLbgvD5d0R9//PT2qTugRLu4IrlDXFgVV9b5NyBGE
AxOwqhTz2v12c4JG13blgNcBAEpA/tMQqmJYUoXSe0kQMVI9CV68h/FbXx9DZ8Rs
MOdrYuI8foEM8l2cshu1tdrfWn38tiehHUbUAK9TKSKezTHyTrsbtRhYT5wJo+Dk
a/YiqmCb4DycKLInrzFecuIJTuAO7LyiDW5n7ihIHKAJI0dLMGRYVYlurKOyFxEo
mV9vu20iJYKUaKeJs/bYdIuVPxzSuBdTD18+aEBjQ5Vd84cekrriBuV/jl+NoiIM
dxnCFS2+LiEMwJG7gLoLJ2NDovGdG/E/bFarRs2oqWefLdM8jwNyD8wV3X5j1ao1
Gz/KqSxtYPR7px27Wy/DRSHlXoPmplDFSS/B4p0/4QswcG9hObtfbaMgNRe+X/0J
Sj4mnlDwAQQgbQ0ENtePg5lVB0mpRq8Mep8UFHKidOvU/EnupQ7aByZSPbl0/qX/
U71Tq5/JW32GG4S2E3W1U3v/aznuE3qCbf8mxg1sI/OjqkHvqX5UkiDpq/maWuYq
WfDN8jidtC8P6+gviO1xgWZ2wHg0Zu1etlSAc32CWF3a8MgRrQsbhlcVzghpOfm/
n2GZIuP/NbesWYclYOkFARUin/VRRXhhyLwMU6Zptv9H+CW7rj3XJnXKBHiQNeT8
PqWKWU+lGk/mlMJ7uWzzlu/yLYHvLtGs4gdrsCg+Fadvo1c70KhaAu8afVu7fGZA
CAu5UV4umi0AM+/0oum1l3d0xKWlsLSuDyFU6d7SxoCeoBBgSh6dfPlzJ3y16Vfp
v5Piu3S04hJl5+A3v8WEvTdn7C8fpPQAkC999P/2BvrB827Uk/KwsrYK5/C3ZcnV
AW+ADxks0T4yhUoYenIKYqQ5IJZxroEoaEzigtic6ajvogRkvUPp9+UDk+COGMhN
ccFkSro856ff3Mnq9jw3eRuvHoR1Kcm3PSOHpAX2jJ8uIMql2GTxyGHIG8nKdg9O
v8rqiXsE3WowHjQTHgMHj4vyiwHY9OweT4SuiBPaB+5184ZTxq6+Jve7Zn1lPF08
ofvrxzEdWMD9gYF6PZuafy/Ig5aLaxWHiw/J68O1BqscLIRncVcJOZPs7EOVD9+q
fVJtxOeJMRJph1a87vRTRsy/mCjcvl3dxvrH26KzwzBNfYE4n3nFMAa3+N1tEi9b
y0ZMtG59zSTWUMfMhEvFLp3QujnTYL9nKnyISmgpEJefb804bFsBNjJXjLNwgxe5
1as6M6PBj3Vt9HQnf06u0YTLz4kuMeWjW9B7bT5zfJ9UukJhfgYwpKgRx6Hxl/Eb
8ZueeScL+a3Fhubd1xTN8A9OuRipuRJ2Z426Z0v0EdyzeLl+AbIqc1v5e/5ZUTnd
R8NOFsZYT3xx4c2M/Hn9wNrgienW1X/KNQxGyfw+Fu4TFrgovGbRk2b6ewxtM97h
9UpQOeh4FQ559f67WoFOrwDg+4MJrvCMNQJVJG2OvO9PZBK/VZvZwE7vAKdxsmzr
rOPVX7TvpMnAGHY/edubXERV22b/9iRf4gxsu9LFBN7N+wA5vqmng0w8ty35GRyP
wWVemCMwY9EA3G0YRgn8AXI0op5IHplbE69VnoUQRQf76ez/Zqzb6NBq9xDleXnf
x7SmkaG+kTEz24ToBoI/1iBw4g/4RXFDBURlFa7XHpDjPffhjVn0H8HTMPDxdpzh
mECgpE9jCXcXxWcpaRB2Mi6jKv7OE7OGNnl7yk4EUE2RNMTfbAdm2b+gmMz/vdkW
y8gcyKP2kBSKdGkrZFnJwk3GaHm3UfYDpMTI0VNG46yYxG/uapW2zM8Yt3fxA6Zx
DC+m1EMi/SrhnEk0RCKr+ibNTyrmVEpK6RdlmzwhNPURuCWDgzAYP0zYKvDaRE0X
sxVG1z544YKAwSBq2TiDzWSQDO5dv2630uWG6FIJJyOt/YXo6AKGSaUqBUAMnclP
Oqc63GzEpvrWRfle3JsbyHso6wkeGXZHsVJdFB/r9Rxk2bVNhONh1FB1dZMNmeAz
WnIdwPXuaRldsQH6MPbEFQmen58CurYISdIyvB5jLlJMhUI35+WH9ljXhsvpu4S2
hq3Zp2PL99QFDVKOmSZxsMSqVJxusyahOrN6XKR6lxunrxWfsi3l2WFhZqQLSdXF
kZnMSWNpb7tX2wFtH307UXSjRBB4l0J0fi0+YqXWLTAh+/iYfax5rSWv1t0ItmH4
E9UOcap24TWSXH17vdcvw2dScH9zLLeJOVmz81INduxeN+ysTnj8t/vOMGYb3E3+
mO56RvHVDuNb6z6rUwJJP8inIQ+b4yRKPEEz+BQ7MFT5ZZTvjEZpe40ugyDunAYf
fMX14ZWgaKlB0s9MvmMusecS1VS8+yfDCRYZ6JUQC8iRv4eokF7AaCkAYWOhoTeh
A5Ar2zFD1B8EizhFwMEDg40iZhrsEhGmZ26GxHcmiUcxj1gIt5zFJIUPHvL0Zlfd
Irx+TrablbqD7ZXO5xNuheu/Ls829rhHEGBjmVRyzwo7iZXF8hhO17kxhD0BluEl
fgmtsIJ7kE+mDdXKUHVlULeizx109Ebm+FuOsBg6n37HF8dB1HwyffGSBUHwCUrH
Z70J7T9IroR3YaisDO0O3BtjWEQTk9gMnHkan0DbkGhhnI3ag960+fKbFVsuDfrC
jiGz4+7L6glpajzt5hT5UXw2CzAdx7SuiN8ALc2ZsdGGwfqPKrbD3YXU9bUh4Ba/
PS0TWwiqHmR6jJ9Y0+g7AK/JcYL/503Z18zIyfKe6DB3W9mum7WC5+f+YjutePRL
A2E2VUgQWbs1DxKKpmcqcuB3g8599GulIHlOnjHxmS6/jmlI3e8uZbZcaJXxFqdD
5OkopSYEmxhYQzZLm2SBOYYQ7a2SRJYwaWh/OVhJF6HGFg0KB8zS2V2OUm4LlmRs
y4AvTpbH0OP8hI/BJq6N0/9VA/aVGm00UqUlQdWj6At73wXIJYs+FnUStkmCWOk0
t4caHmhwBAALLPLURUsVEDt6GInO5XTRuSCMi4Fp4Fpc7FTWEwfbufBDIYR+iMj9
ZYkE9EarUjrTKoXBoP0SwEbpxdyEx/BiGd4h/23e2StoWbR5cEknwjf3kY5Uphc+
3Fbwf/0k2VV9FPBjYiBTUkQT+HhhwECyxKXL6ohTrcvWqLabW/8KAmZifkbyPepG
Rh6Z6gac32/v5G2C6hdhK+/mKUPY7kX/dM8xARGP0OkJaaaLGd8aGTkdnTD9gu0h
Sf48qYf6U2mYgEgAN18/1K/DA0PodOyViv7EnQAmuq3AvlpmVPj1ivrm5/EHGG5/
AN3DKa/cUzJlVvrXYC4Pq9rL62kaAKYM6pCEcECTQ4m/xr6PX6vSYJuG5p1hVTUf
YEyncOAGErjA+hpZ40f2zbwQ8Oct/JxA6sMIVWSd5ThUE3rVHmDn+jRV/FGp7wuC
+m2aP/oCLb/tVFXzDl6H//epBgjLlYmTzUyPQf5OnUA8nZhL0NxB33AW2ALwJosI
ZoI1YUXxnyL4lX2GagMuy6XQJ9igv85QvNzZ5x4rnEdq41KhEQvIcizj/eyBZTeF
voncVYXxXvWX2Tn138bigfy1gjrDMSn7QczVNrtqHfAb+fwZlzRiH75WhppiP400
gvJpvJjnT2dRW/eC/1WaTTZ87qELTCEay8uSJWzWpMaeHZoP+ryFHcXXEJLJA8Uh
OS4Ysjs/wDefPAckOtAr9tIlq5pRcIjJ2j+rhrs4YOoXqfEOh8AE4RZtPhTJfR9r
/cTrhacd0GxCea4YLxKOYthL+ZYS+qkC1wW7kp5TTZM+fUYkw4ksw540pa+ZNjOO
rs+sS70pd82rinpcemJmkT94GPVujnQDEIfgV9lheXvspBKt6APSngPawrLhmaEh
Ero8iFSHrES9rSp/PJ0rpTjWLggfXhV3vBqBjEZx8c0RRQdLddYgGb737rSe+16P
0SjgQcWGpCd/t39jfT9Kmh4jAVsDRYhwaamAUrxcIrSMq9wOCSs5vr7wr6mN2Acf
hqmtjYe/TAw2g2rGGhOJS4axSjf3jUL9nZxi8QHbIMcHy/YKDN/oSlafZ0iZcxnu
2sfsQAs27PmoSKHmWZensVT/nkTXGxKAZ2gqYCM0gXA31Y3m7fYrkpg9o+nyWDYp
UHwN7Roclv2W0t4xirxknVFCXMIRrXKkU8HlrjeRQgIqwQ4FnvtG4309FFOp7UnC
JzNjD03W0YK27t/nZiZS68DIHY8H6LDCPhCsZpmENyKKnNXd+NzDL1Ht6ZA/TS+z
UpKWja7UcRhHFOGOLzeVhXATsc/ixY2RrHpFWA2epd046QjwfLWtmVBu3tb1zCdG
PvFcBwgCVUwwBpMZnSQY/D6clXrazojpQzEY1FkseVUga8cgFFKskiRIbkhkP+ll
B4Va2k+ms9oCpKgitFROpBnD+SHZwYOQFSO5R27ejdSJut/mvOpajhdiplIo+S8z
qTZ6UGQ0TSgngePxt2lkQsVSdMuCcsRBXXSG8y89pVsL5k5Qcu+AeTEWHocOazG9
ail5UllaZhuvZGtNxPapa2lOar58mvArujhdS1jKzS7n8SIwtq4n6zgfT5GZdfxx
oh6iTH0jfj9AUcF8I6W44vVVKZdFvmhbHko5QgaWSvAYOnpJMskT/JBhzvnNJQYn
EVmTfk0lKVeRj0cKhlMJLL1tQKVuu538XZKIlu41HTI0HTXVDHGyyywNvzle/5ut
zm1xs8v+OcNr0Yv/Hb4bZ4tCvbTmsF+QipsJhS2PfdY0lwmQgFyYungxIvQgQ4ju
Dt6m8F3Au7dljI/zySLxAh70WqzrlLr3QNJpyYJGZzvulb8AZKSi+opS8JSmEdea
hfsrgDJybfbbFrWk0bN7eVig72+6Rd5fCZn4pgogHDw360+9u7/iJgkELzSJbO/W
n7wdTxrX4Lj1NyS0CfjY6eIYLSJdtzeZza+h1R+HdETQrclqyJfYjKYeDKqmzBDz
Dy/wqHuvyEUzdcM6OfcR8o9tah/SFe+DF7tkuSO8zaIhdjRba95VdkUc872oFDjw
0YgNXj1o4I+MUR/CO8o/3joIxInvgZfw4dSn2wTRRdc=
`protect end_protected