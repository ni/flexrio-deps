`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTLkTmGIPhou9gzYhuquNWHaQglcJPF2HHF8re6T0msPw
MLd+HKnk/7Xr5auvEzc/g0LZylnVdAJldUhqGEOUWN9/KTPq+OtPqgkLGKUOmG7S
Z7t9j0sv2PEXSTyHpUXoQenBOjhxPr0dcAASNwVYShNQdeefFBDP4K9+/VEbwhs2
lk76mUyf0ZydvgoGwVhCkOuu+jHOx9e1O+DV9GMOjsOOnuHo4+3VjfZNKUZFRBuK
dlbMh+w8+od5v1CFf/pANJa/PivcvvChf9fnTt6z66MhbtAaxx1pM4652wii4hPR
+aHtTORU9B+5oqTkLprl0R7pEDELOlxmRzXz4+63QS11ttvu286RTSQc+MYkX2HE
V1cuI3chXSpDQJIXtX5C3GfHB6gPZgDxi4pLeiTME3nPWMkxA4SiaDAJjDfAOV6K
iZo2wP3dr1gPED67xmDSYnRgDDG6Z2q6LJyVfppl1jqJ1M0SQcyqfCW7iXmhj7aW
tlOOUkhx6wp4sUpaNMy9sxO0CirpG1Xt/jkOSAcnd+FK4TUnaNKt+UMXrVNIBj1A
1ERW/LpzgDQypSYLO56tsBKPYyQ0Jvl8Ht8Xik5xF7oYWIJcbMmTiq0ncQmRUSCh
hJNaVqIySZmuNQG4evPlKpm+OfnROjCIwDlMId+hxKBxg4/ihpVR9o+xk6IJzYAW
7C8Nb70nlAziTEKB1utcDV/iWp8IRqQomwJWO1wWH8pE0d2yC/DhvYX0l0d0JEg/
07tGvJam/wzhmA45lPUzyPFCnblfwizqiqtQh/nSGHySGn/2wpb3N+qn7843Janj
dIpZEPdmsw2dwZN7AutPLnpDq41EJ696J893NrqNu0rXIiTwhNfvJmz4DY0V+MIh
WlttVd8JSvQ9BAFZzHHwMGX+1o+UMJMvvPuM549Y+/OtTjFN3r/8BHx8Zon80pBw
nRqKdABDyE+tefP6MTHdx/xTkougDj0t+gvxE20usJevu4iqqlrNl+ev3fVS/MNv
8giYK+FEjZp9B6wgXOZ26gDVgooVQDSU5irHLEmoT39ESHsjTprWTsEBK+OYE5Ws
4tNycC4wPfbCHpUdHumGfFVpzXVhxYkrBtUMpzsbTGibAVLwSXoYzND2rJ8XoSjW
oZGYNVfvWDLSTAA0nNkLy+iHbb9YVbwYzFasHbnU9fVWhRQkieAq3ArhOIFM/Rpa
StzX/1OvZ3NlHgEmn8C6PZPc3Zoj1YHsOdf77zSnlbjBdX1SRaRQqn/FAXO2JyYN
zziQM0FBEUvCj4yTo0NvZeffz3BTpFC70hhYlRiYS/hfqe2LRcyyXhQwTTFRd1j8
jCmxss2k7foMPg63OrZdfVQAJs47hQhNqaEkmNspZiBT5H9CgaTEf34KvQV7x5Bq
/rnN7UwXTIRDH7yYGu8EovDvEuiYfNKkfAVomcmXxP83kka8FAKLe4Zo+8XNlrG0
O0XHvs9LstXUHGLAQYtpe9zmmGcRHWK+mY4mzO4WwAijUrQpZmCRT99yVOjAEV2i
0z084H7LicQUtz0jj3w1r633sNLReSKb9/20EyCiBl56VlpVmlmsyAWFd4trzjwq
fC+n8czqRixMuVUSyp/OG/EZpu0JmsPWP47wSTxMEXgUbmCBeRRM0C5qqZO+A3Zi
yPZNhhbh0/Vha9hP8NJyz9eqHYZSO13jB8RAck8XbH24Ox+mafRXHg2TTbHw1s7F
tss8wYn0Xbqnu3BESXXDGxvJxDuKxLDECr0Z2v2OoknBhFu7j630F6eDIe4I8rPW
l3PbyDf6yga0GBnrKi7o9WQr/mFZcDCJfO150C8xomo8UPTvNdytmQyRdlpuuT0k
L5oyFuCBP+W2tJvncw+0kO1txG8c2EBOKDaImRNZo/+SLgsmkQ9BWE319S9c1jTm
MaouRRtVkUzgz/ZTx/1Y4rgpie91lQuJhBU5iPH+I9ASq8MHLciIjthycLDeseON
/Mnfmm59TRIn93NuJzRQ+FPrJEEO0ywxIc2wcO3pOjT4wZX238KPNqIdgjUV2ygD
Mb4Db47mWNKK8k7lC7VWZDLZQJqXQY4AblKCLW0mdX/7XGXz6L7deXOZVtvAmeqA
4iTGRn0IyYhodJnmk2PLgUdls65cyCrJMTc6Lh2zucrlHmoIWeBZwP0s2bPSTsZq
2COa79Rr27CHpLrQAiTO6CtceYABGtmK+gBtlxNRzMo0HTPOw8lLbprW7k3jC3uC
rNBayLRSmzjasIW7rBmgJSy5og+M0IzuxZ4K0HSXND+cj9of15LdSEpXic7OxSJ1
5/nydFOrd/sU7ackDEtJ+fvPZIJFLhSSnuOcT/Tu1dTJaJ6H2/9sQnBvv7siV068
0jdHYMTLLNEZRq2Q3D3zXoth7Wg11fc+QEg0sJBxTAi7c3e8T6qYRolbcWnmLbLS
hVJEY+KIviQVFFFp9FJPtwOqw5pgV4Jz89ndXle1NtBk5yAp+hw18pcIz3+IZiv5
dwGo02PLcX1BG5IGyjm227iYZsr5PoXavYiA0bbbMU8Fv5Ys/rOjDl/PLiE8agzP
1qeFC8+s4lBu2/LjWie9wl4Ny93QxLxbw/KdOC5/q4QDtI/d0ITU9HQG+z+2eujx
wn5rnwGfTB2BZoU36kuIqncNNGH20AfePnaDpgtBNFEr1gqjRi98mdFRzOHYjILy
aWWMs6IIXCpJt1wz/bFdZSbeflvagCBqO2QGhToU+ZJtrEQffQHwCSAg5stTagFq
0TL7qnbCVlk1CLFyNsA3y2rcKcmVnPC8+qzeAXpXI5LhtKO+4WH7EI8eztVPlWHs
mMnKUyCTBF2tl0/wBuC2iceedpfA8KVNsuWRX7SPyoD9mp3U7RMjC9+LYszrwGFR
95o8ZpxeSfIum17lAczEDDVI3MVkeos/frKqVIqOrvDcMgHAG8ObzhPDIElHBbT9
QXj4Ww7J/sgSKeyTz9pfIBOfLOdKFpZXu4IThbw69HdPLBrhxjPhCo5Gu0OL8Ahx
iF9F8wDSuPwYt6IOuMEbsObjmAHwtHLIgkXgNN+voy8agaykn9auRjnqsd1Z5qT4
U7k/gNkWyvhURChS5Ddbym5tF9mHOtThRpmj5nxoPcbm6W5/fLnTlt1TISQWs5EJ
0ublR356pKjJpCI4pg3WCJAX7Nf9Ki0maKgf+mt72GRJ4ry4xvC/d9AUFhOQ9A0y
Y0TPvw6Up/Xik/yS34BZVEkOJBTB/JpEdXpSEguEQPOGDUeo23NGGvPCRZTLz2xo
W85sCVrrmgf4lIwvqztg+e3vFMAJD1+3eTggVnx7hPJDOpX26gPxnKxuGNGDqGcH
9GAY117qOtj69uVO88u9wn6AItx5M4f1+A5xPBrBCTkSGrKnpnz41YbmjtmxZ0Kk
My9s8Z+5q+C8RadJRZS9og+4TYry9efrpS2NWosLq/DYdt6zPI9k7lBND+IzuYD+
iTuVXQeDtEm8LZgahaaK7TPeIFQGRzmRaSgWY5PtVAXfurc1APXFwoFqA7AwRE7/
84roF7We9F7jwtrYGD7VqR2GqG+Jh3CiwHNNvk+isMeXXs79y3syX2mFl+yt0vKa
xH2HC97OShSZUfs2iYqfC+jbYP4rpI7UueOj0FZQ3e21nC8cR1VhnvHQy1XLywgN
gHvd+zPL/5EP0RsPt4RNj9fXQ/sU9WDVYa1Zvzypw5QE0qLmgx9chadmuhAXUz+s
HTlH/iHLcTLqfw+ztUte0YII04BcuEWbV3D9SQg83yPmnLNjsNPnG9mjRySOJmg5
1aEWU1tEVCS6ADMlfh7OumGtYYMUmCUsHQIVrYfefiv5hULl+bdAORtMh7Cizotc
fYWlgJ4bJwMQj7kyGqmfrsWBCmRfH1OTibCz5F3oN0MvBTWHOH0Ipvi0KWQaqtVa
KSo3HlqjqLjUrH3Dem7AoJYyJw8gCGqr/H8Xt5fqLAoKp/+6XoWHX/QAbE3gPfNv
MBKzFGGHe8by1+LeQQumF3jk4LenLv4hQOkyNf9XC5eSKjN9PTYlDzGuFN0s7WUt
T0y99HBCrUKn3ICxW3m7NWAusTNlMbtHjor5rUUU6KZXVyERcTol5SPRDfY5EjF9
uNr2luExeEWJ6Qx838qM3CIR8D+j08xlEldgmWzDdq2H7soTBttRlwAYkNOBIadW
gA2/yKX9FRxmqbInj3ByPl9eM46GUhEmY5EaJod0TtBHckf6Ka+ZsM2NGi+2jrhp
ya1PZ1w3PlPaDKjff8F+ZRj5CE1d6HVssVAPY27+BdcH/OPFlSZCFqAxUbR4MFN/
pb69sCx3V8nRjXNPmkgC8vX3YCya5tkZrEOU7qvmaNvtDdi0KB5TytTvjVrt8Lgz
KU5j+2+KcaLv4gDB1rO+ZZGZ6J+LyLy7IHpQ0nq4QKTIqTZh2xHzaPZ0EaRUk8iN
WxZ1tbFnFQ0FkdvwlePFhtBFMic5NzhACcLNgchkbNbBvgl5xni6IjCtgEbr78Ii
6Xt/FZDLbkp/byvpU2sQZnuLvg+wcnwLbOCAdxAfKhA3hxX30snkZRtMoJXYrQwo
5IBTHfKW+Kk3VVi61WicGVRbxTYg7XxP7SPyDgcKNenP+eFA3/GdxCz1BQFnpfKD
jKiv/M5tdnpke73YGrR+WlOv8AMDzDxCcw6BUP8abcGxT0qywlhtu4JXEB43PQBh
dMf2AGL+C0bpZxN8CMl83PdYTXFc1No8ueCbvOjXn4vI6IJaHtER3OmNquM+EgdP
oeFMEBMInvJcm/aL27U5DsYmLbc0QHYjVTpZtauKhJGrgg0ZJb+qJKzIEfFvXca3
WDi8gYttNAkfdRn7Ki3mbXpGtQ4+NZWgkzvXbfMgd7yNKiOgZtgzLN2b+y1tDvLM
8QgXYumg1ItdsXQfrXRRsbxaYKhs1gU5CXsMyqdwVqgLaP12Viuk2lJr94Qlmq7n
sP9XaOkzXDg+erl79rsT7WjogDY6+LeF74pjeiD408KwFcbUUIgFKfow2jgoWqoq
+PtOSvGKBJFtujXDOSAQbO+4/+AJ1dWQM5tQBhr1aUx5nk+lSyNIGwdQ/3sL+a09
24LKAASHXExage7MZXhoYaObTr/3Ypu4T8hiRVViRkEayutWtKd4MdMxUhPP9wGG
yG4sp25P6ghWAGH9RNhCWELB2RwNkXWgaJg4Dt4Hcs5Q2sqLviN93qgPH5v/jk02
EfaHjBYnv6lxQSBP/K0upf6xjORs1QtDRP01vYUQJ81NEovzrrPhVAOvX2UXczmM
QlMeGslFLp/04kNs1S+m++s1tpfrkLSbsjt+9byu81QRajidTzqu828u1Pljihvi
58q4j1SJHm9zVGc9rmX+/85yWa0QEtI/iW11JmZLSoISYV22JyqA9pAEEafTqub0
Rr7JcW4cnPRMQaAvl8AdwGJIzKagiWOGUbdWlDz4I3TuFY7/M5u6CODoqip6qNmn
UN3usv2icuvEiiUE7urbGa7QbHm49NsSUota4X/Qfuiz2QKUu9Va2idFe1kUnlOD
O02iGMAjyPGk0tS31CD8r6DEdZCF2BHRJA99BE20qH6qp2qaSvBqC11wzCEG+dvA
QJcvwCXF9936N5sVYJ3ACY50iXKu4lS5TNvNt8y2gJcvWoDytNg/hVMiJecH7fQG
FkW++Lzz7Da3bHoTt1890FQ0zm+ytMhgB4WeJ7tWivAVoKUWsKemdp0BxMYELgOO
mvPwzU2UmfCyWSp7qHoZZG6BuRyKt2tn/VBkwfcehp0sXShoBChc/mJqczhpDZkz
kk8b8owAvchhfaPtOd/5XrKe0Bs69TqdKcUCWtA3QxKgyucyENwAlaD+cG/Cyvfa
is2DNTE7Fs/otgw/TkK5aXLNQQDEpp91BC9/mkOrEnPfy9i/49LNHvpQWaErKml8
kZBmLbcLxBTAPCpv0Zcez4X2f1zFPgsSS51qiSNmkVJPCt5hh12vHVaHQkSH9+Ra
ryj8pMALx0tuORfHqZuSyR0vtHC0dO7b9GjhNxuCcaMs5UIXPANKtqdcQgXLpLB1
o6YrLsV5MjInmbDVm590SXRWDSWi8EgGyyrQpigZ95DsPMOuqgsULKFQDscZOsGq
LgPS1sqHXdykTbYbuv+ZIZyHPMMsmqQwD3XXVmlYIWcZOEY497OKk5Qz+mxZ3PP7
ssgqSSqTyU60h3otT8RuiqEjwLLbpv2KYAoKup2i9mWY8eAQU3K9J7wumW05EvKb
S/gpFB5q3BuZgRVJ94hDaIVxgRAGcSophCtrLIaxXG/dIkUJ27ow6otx8yk5zg35
ub9tAWfrsWMi2qQG9znuu/pFP7vr17q8WfxMyILWqOISSB0qmdzKnTb4YfsFcE5A
C18vLgbMY6xphU3W1iyH8u6qj5UYyDPt0CmaLng+4f9CeWe4znrNzsDvoGm8isz+
aX4qOu9LfGPjhm6lkj6BL9oV9Bk4aZohVG+zuWzB253u26o7Kp0y3cGhRu2DbaI5
9sTa2lvM2/u67wT9qZ/baARB9u+Q/jceQOETecRy819Fref0+mQu5YUq5uf6km5l
Nj2b/FEZyQ3QU61u2DClpBg/BzRGUU1NReOgTdpDixwSfFzEICfxDQSkQ/tLoCDn
V4Tstd2Tg2fg2395J7FOkrOKWhC/BMWtCiDNpf5S8DHxjrth3jQrzrW/P0ShssUd
Hg5QHDXEwx4rRzoQjp4bSGmmNuYOvb1U5i9UPdRLBUenlKcOeuIBmYJkX79uyCP8
sXAdaD8SdKfWhe8qtHSpOlDcOB14V7nuT7XAyavIy78f6NvYUEVbjDq7Jr6PUVTM
UP2wslxCbUVC8ycOgmZWypou1+xQa9s6gRep3p4uawVPTV+2lnECHKxv6K9V86jI
XGYzJ1LimlXBsCuTsy2YVuspb40eMznaj8E19jI97ciMCXowFHmk3XlbpIEoRJfj
Uw50MdV3MpCGZoWuDdGwdeWCCrL2mmwMdghE9PboR2Rq4zCj4AqJMTn//OkTc9D0
8UimWs+kPMlXgKUJg3ZBoLwmDb+2oGEcxtVlKno+TN5IJbZwY457qujA1dRbNSnP
IBZ7VlVqaZZhCvLA4KIqUb3/Q+4xcTjXmIUrR3sRV6bdWEW3w/D98uL943t/RtvU
A+qeEtD7xxtX2w+NtmCXjlz1Y/oObjeP/pScEo2uYZFDAxEPq1QOiZ3rsM+yBZ7v
vXF6PS0qQafCI4gHgXSJmHG3IHuocYfFX+FrT2UH2rNWX1pH2U8EV8EyZ8S5jAE0
cRhOv8cs4HfH7OUUTiqrMLuF3E8FKcdrwtxLNPDiQZWM12DXKm8w1C1/ACMUoJpK
Vox1nos42mfWKV/jHMYWwvr5vC4Xy2eaiXc5sTd9/G7U3wxElAFRMxGVlyKifOBI
cG60z8sM6egtFouXtg56JfnzyZ1n51N3AXpgKKGwIsPoRh/cDjT6L555iGvDJSnA
r7dL2/tHAAAT16/SBrpU6/OpArWD/xyLiSPdKQJ6oKXWT1xPjf2lPYU4ULhnL7vS
fbCej9k8deCOGTalIc4YPWUCvv1BJOLgE8o370VdbA9VMRhlJI9QwUIJFb/n52tF
fFvGRyAkRYWdxAO3snjmxdIj7qTBsMpugMzTfgJhv2QluIsy2gocmoIvbKzc3ECf
NqNOUZauQyoFmyZVFbJ0fZ3KS9M7N4cF5bNuiM6H7UR4vqvOhN+9W00Ti0JpeOQe
CuqXjbTMMPR48VNQv29+Yj8d/BpR/7c4gbqOqF/yuKHkfVI+AAo7qs8f/FDuTR7Q
xbXgadK6d4UPicGQ3IuxRMdr74LIj3vHIeJWCARqyKuDjqKYta2eAPFVAoNZi/bb
cHlekx6rObEq5sGQHqlYafJr1ZLGn+IsT3OZMn0suEqrZsNlATqjhY0B0GcCyR6h
rGjK/gmur2PeUJKzBXK3dsn0GATRXJC02kmxnmx7XFYVd0QvqdOHHEwN/8F70ZYl
q17Lm5haUJBXsPhdvVAQRx0OW9pmbDhrMs8UwCb2Hj1emgZ8+F9OjAmuCk1DbQBC
vbfvlE5nKkBCPN56aX+qOq7C4ZQ3Vs540VCqVDnX6xPNzrIIM86r5X2SCfAePgPQ
hjYRHCZVwPQGyO2Tnlar0XPoZ15TNupivZ7cY4cOHxAEn+Wg2bx76bnS/tdK667W
hQSB+KS6ICDjGPdAWsFr/sUtA5omroYQrG40/A/l+A7pta8dGBK5AVXYW7UDJSH+
VoFvfwA/GghNV0BTXKHiL82Q0/I64NkoBkzEUdKChtoaW65tKHsrr2xTo1fqT+Ph
c/sMG9Bp7JmM5jLgTjsok6UO61X6Uz4KnCQv5cUbnl9/JJbNmAQEzQD46QYgu4du
T3aotRuFT72X9bx9nHbypBpE3JIwabIYNTAcroCpf7bwHT8Sdfc3nye7fXOmyra/
YcD8AbjsWWP6E8U4NQBbcs32m/qmiAiMrz9Ncfd10uMdP+ZCr2rBQRuFqubegxBU
O1BKNVAjMFuPBHKScp2DUy26cQaJFOV8luHX/4xUqJhqSdKcSdkowR5IMcJZ/P8M
nohS11YPe7H546cTZgA5O2S0xPMNNs4VohpSgprstwUP+M0/V6lvXEDo5rx9a8Za
dE9EpePvsi041Tc12YKsZGcdJYDuAB0ii99myxZjIP9NVfbQyL+s3ncWNsygeBAA
oBmExwmA0qHuSRtyByKboUL42LrO7tVernU+P9D0UfDOvJCyJt60PKhMHiFIPUNj
uBQ0ZsR4QOiWoH+pLOUuY/J1iIZNvC1z+ZevYg6d1hyoJDzAVJ2+xUX6/US8qDB4
Xd3j1DP7eRh3daaMgEOnU/OY9WHMUOnn9cngigrDgYUVxgx3vgB8R+E19h0rrV5H
dqJuULyIxf5gIzrX23A7hDOWitmNzuXF5r9CldWUQx1+Oiu+a9iqZuiuttbh87kC
gPdowkN/FhccMopVfK4cq77+XfUKCnesO3eCMyJzQ6LKAV1YIUBD0cWFQUDOnL28
7bjcPYhKzwxAzqIx+76+UWcBQDJ6fQFFYu3/gvjDIKdCdpcAnoQPjMTdtLWSmezd
3ksRfYxn0MoqQzfOrrS9eAqQZC9wvDWEN3ig1qTj6nYlJH90l3mwVza9d483D3Ol
XgVAlSnUQTmJzTn41fvjt/jTWOqHWZ2o4zeH2RkQ16tjq7dxkDk6iBSAeY2eReP6
ABd0XmXKxy683VVcbsqLnroOts5V8iM5Sz7PqPWzbE5eiJF1VRJfu+QzKQBpfHBH
OD4vz7oRcSqUUhansSMajxxRqkB3ZP0eU4V0GfU31dRuXbGmNCRFMNEt4ZRomDcs
mRIBJL7CqPoRtjrQWHOex1nfEUXD6/AJonxi3z/eMnxS3uhU2Uj2nKtb9DIQ/NBr
sgESlX93nxF0XRkLPlrty3pDutHOOyNoQtSmviXBwQOmnbwmmhc73IN83jYcusHQ
JsJdSGqlC9+4AX/HA+04Qup1I7oH4ocgH8nvZ0+HdLcJG/11uW+Iz/ZVy+w3/HKB
444r4ZNd/iXyg3GU2rnhbuA0moLQaIUizJYxjRPu+zXwLo25k67348Mq2rORrPeH
iEoGwIvUdPk4N7NN9W2ntAqDAkmNuSNx/OtG28mC2ufvQXAAOGy4kS3mWQj8BAtE
kcbPeVrOi8ZVeyPLidnTccW3QASoP3Wg+5D8cbb19FkJM1br5WQV2ydf0v89RZnJ
fZkC6mJxJoH3WlfC1ERNfOHD0QkxOvQ95nzVlIjemYjwArfJ/v9EZ5FMLf90C7vK
1/EWyfAlahpXf7Ir5rpNi1Fi0bHfpwQCXB6kMbXjHi2BAO6Om4Ot7qUEuoNAzoEn
uwswagchuL3/6FBFa18hTVlxHGKWECA6PzXkPHrwES2xoWKnZ7Wv9MqPWZB5zR6J
9b4rTIlNHEK9jQLyBCeGvAHvILt7U7vXR4S7sbF/vnuR4zW+5FQuWXX5sb4gdzLk
rNt+xnfv4xqqff+aoF2B6ufQ1pH6UNhqpQRlhHpfd5MkP312eF1dpmPNzBW0nPu8
i19rZ/qxSMCufWpecTo9k4nOGmPhHnFp5TJeV8T/n7Evk6W5g4tShE1RUj4rMR3S
Bb5XGN6AqBiCBdSVTMqf+PNGXqMTkkgOK0WK1EQA4+ZzZyTfMY/pv8ZQT53579KU
jAhCFvHrVuM+BqrTOGdpWf6RC7a3gKauscbBxET+PBHPHSSYYUIa0+W6SLY6ABDq
WJtV/kIazlKb8+NXqVow98uoxfxdzexuinamp5d9XLBC91iXdXAWS0jZSO8FCbVF
1kyPVNpXnmMbzsz5cEDS5/uFxaDRyqITSZRfl35tTHt+Z6P2339+3uKNupZtRpyK
v4zeWpvWC0hWPpmuNG500ekesCsa741spMptZDCMeQChutwvn0mRICojpfipwi+v
Np4q4rsyjRjdFl0aJJky1SQSRineJ1kyK6o2qQfSHUCJn+0wJ6GcQDGjJtY8ajMU
wh6r7I5VFjUnf0juwoMDFqj1yahZuSGm5zR9IdPvtsgFdRIwnG1W0VdbUDaSzEPj
R+J8DOpPCQDLBJxlwyd7yaDow6MYtQZ4rS7iIAhcDGLJtLnfVksPnYqOfCuJ0SUK
LfSH0V2dglZWKkprCHZ3bx6rQJ83XC2cz3fTx268ZJuxoHjSgQchN6z/8bW0+Gh3
TwQx2r+zHaU/kD8PFWEhB0vmZ649pOgwUlgG4TVn++S5xDbtGYgFBYsweB9iN2vn
/BXrogFMrufwIsrU50bGjiH02JFFRQGY5K7xeynu9hoin75TAgLbvu1zG1dRB275
11S3Pn0CkuNksStbOnftXCI/xPg2GeWWVymgOAx/+OVb6XVh4FBLwOwoAfmJH0vp
j7KLpjk9Ezw7xrAIwZITUoOe5cMqctWqdBqlH0H0AfzbZbSiIL+qwjHtHYOB2jvd
wLZ0a5+4qOijLELUfC3an3qSj770+lXveR3R5f/YFigYk0/ajba6ph8MBYkCH869
zvx6R4E5ulDVNVcE7J0fxZcGFVFpr+LSSVXhczVGLZdOjPnlqQYddcSBStKWGm6u
RG49+qRByl3gcM7143aLwNwWo9E8OCF59Fpx1It3j40eUOsOjHGbl8y0ocG3Owky
+jW/0w/2RhFTrrFrsPmp3b1k02UvAHAx4O8lhqNSUjqNXxY2vESmsYvUn/UvDbxs
npjaMfzRqt4PsmjKKPhpPqKasT56CtDxV2/78xbtJAR2uCnxNWI4ucqZel4JdZiI
CHbF8/u9wHjLTLewjmhbSCnsxlbi3jDHs/OiYd/EMB/9zOHiIeH6/U2wSpEOH8pQ
ResoKKuL0QTuE2PmOxXZ4PsZxS/0HHL9j7zcwMwiy6GR0f0i42RbTNCcAcIvsz83
lfEct0ejquUx+6UnXmbnWaGes1tGLJabYFcmNLo486okLv4Gyr6BWVDKo7IAA2RG
Vi14DchR94dd+di+bDAmOCVFCyD78wIKj+yOM8Ul0k0j+jy/84Qzq/u7hlDDLbFZ
LLw2V3lHvODIpDM1uh2LMWT0s+6Z9lc8Kr2FQ+24YbwOB/QqDyYvzcbXbBTWlgVU
RpXvy8bw0T4cX05n+Dw5F/a37QqL4l9duJvYTQzp/+OMfMphmeeYbuvCmGla0Gyk
rUEKHKR5nWuZQLHHkitV7XsTErfkmoERd90epQ7bFWyBXKLZ2wKe8tsUnkMVGYAG
8lZoDyDGitwudoh9d0Fm0v/128B5Eq7Gkicq/14WlqgEupG/DRT0hiU8UpEcEul9
sur/kuvc9I09+JEGTCacdUdng+b+xzGct6gy9biuL9gtPosovybSpHxvB6pY0J8w
w3dpKL3M1FK5ejAccI8+7l0U006839VMrP72REroZG2XhPVGbjI0HQvvFXqphbP2
s7wPXS0LfMMMa4P9LRQpY4dih+/Nkejo64gu0U95cL0e55xSxLxopwW1Go2Xb/1k
N4M2XVr04q3La9h47j+O3xMBfJu9vwzcMvcrhdTrbX41p/H9ik0vuPngXs1uAJoT
gnhBBrZgYFaA4pDy3ans6YjDBiK4Zf7IlfEfPZOtEONLrNs+wcfDdhXbIfAUKMK1
VmxOBNiX1B78ijh27QKXA/RJj4r3310FhtTH80kOX7aaI+nZNy0QApT7z8oh2Yey
OPqi3ByphEIoi6YjdvzPJ0i2eBGbg4S9UihKsvSwzPB37g7JJu1mT735LD06gUm/
qddq/8X/RjouxSVWAL4vzRLXCkP1U6xmaIodOTEAFqAY+sVr6U7qpvcOHPCkQhbU
FBIPg+d8yTOsEvwSD3N9Wxip6u34iyvEmJwGT0QIogGLVysg1Ft1xHML3qZC6QOh
jFjuYhUgj57+UtVFLoOTgnlFzy/ZwwqMgGHPsHlY5MeDBMc6flwgbHhQx2mZf6cw
F4x03aUvNyKn9XL65bQrH8HIFYyEcmkv7Ukb7KOTytjvm05S2kFFrYHoZtDYU/L5
u4/FngrJVy7EpbYvmZmkNLAeMqqdYAY0nkhBdkHPw5QJxSDGM2cLSDt3NyN0wn5e
fDegiOyLSzzQzAgoNa9s+s0QCipEM0CzSNaJNvL0H0OO79cL03RuSZFbiV+x1hW1
Q/M7hd7apD2Afxoo+t+ysxd/tu60O9+/rAvvoVO7/iKCe2l4Iq+CA4J2we76lOXO
2UrtszyW5cDEJ72eqqZrFf9bhMxUQg3MkQNCMuGGzf3D+sNrbqshKh71Z9XWOv5s
9/OnbUtBEt+zb20S7deJlzMeIMPcQILEZZX9v5edkCj3Dw7Qn4d05vBeUIvI2uTr
NGyPBzecyCE+HGzXSMbC5sWYeZJ/lC/eMNXMKVgBvJ1NQpYdxK5GMEm30nEeYb1V
M6RatOG8j6zts78S/x9QkFbaFNGPX/+gg2CFhcGKXjC4DioPPMyELCv25xOznCaw
hCYbvLqmzHIi9MSaFJKlFANmOYuF4WGR1KTsZsQc9xIcxIrxY2wEq2B2Y+Qs7jGr
JkoYra8OHcAtolE7w7alz8ltEFAPU4ElMytBEge94VGmiQOZsiTjFpnDi8692n21
+T5RH9HjAZI1siRkIp0aDPkeeGTcStAXHgAByinpLX9rKqvLJXK+y2IUcVSUWwt8
/lTqwOe/SaDHVFVzw8ypVMPbnTvScstXcnHyfxMcG8PYwRVQuso0rL0Bkxq61QVK
YX90Stu3Hcio0AwUvP6/YF8+GaL+ArM3CqmkzjvhZxzpyYEdaVDFHl/PfYu3jnKv
hb5HWthmNoBvLUXadTCDrBPt1yPav8a2FAn3CN1WzH18C1o0IqI92ESfQ/fOvMvu
MLF82Fns7087IAgL9yCTpEYo3KAvZFKwaQToYFp4qe+ZAtYyje2odvJpfSXMRnkK
Lgk2WTpmgQsacy0hZtI1gfgS/pULci7ZaHGsaw/Z2OdGpTC3aDHinGpU7xr3m/Jd
2kJiem/si49+q79zkFHpPHe5NJaRUm+nesp+I5WjNAN36/uhjTQkMEqO5f9u/Lgx
AdtMgrJCRtbC4bGVwfLwFCBG8o3WnE2lzQfllnIS7hUqQNJQ7Kwkty98OoIvfcJ6
nhWJU2WmmnDRE/8hd8ayWx63BjhDHn6rW56n3RCHqeit+X8iUaa6yF6pxs/Gq14g
hYJvtdw5WvlltWswqsaBuxlNayGo/WZ4V+q3046By38qeB4f3VjHGDFUMtwtIj2S
V/VSrA/3s0k9S81aN20bd8LA4HEa4K0M3d+LNHEUmB/leLThyGj/6Kv6WsTSm22Q
HzjMG+i1ZXqLP+X/JxE1prf84suyMM9Zf3GqG2XfrZg/bmJqTcaIMp+1CTLxX0xG
BGkdqtTPn3WhMvN5FHAh3sMDuAWNLoHdZTvxXd3zEofiVlz6i2d6hoSuJe73+mpE
byRl+PRFl1F8WjFXXzw3+nHnoTInmE7/RbCOA6g9SsKugbSOPTSuXgGhzpeRNEuM
NM8Txoww90VuSS31y3khvT2NmxGkMn+ApH3vVapSta+yWUOreJbMGmYxAthi6y8i
Cpq/6G/w+Oze5ZIc2ce+IuM+PE13a+LN3gMajI6IV3LoJZgcfjlhDjmSYwZSQotw
yY3KXlAYiqvswJCRF3vhYooJmk6rrv2d2QMXO5fEdTXofCbPVZ1FqXH8NmSGGt79
K7D++mPQvyJGQBp0fTIfUF58D3/79MGFX41UF2Yx+Vn8YJPPGwFNw/jqhBHZLhAP
NGy9qydeQ07gZ9+WtgDkIHTCr3JI7t67OBZmnJQj9wtpfREb6pknwLtd/TIy6jcY
0Tz+QdB4VZw6+xuJ6cflAwDndT3JTeFLrpunDAFqjTBNooEZLZq7fcxy2Swhz346
Rlpo4OrwBg1SWY8TEOwhimWbvYj2EXzJbJGHVpVfoYVaaOratBdD9sp0IPkKlN4f
UbdZwuRRzsDgkIBszm0iPWVSmNTxxNJLTqISKetguDvM90uJ6k/wVoPsg1S5YwNv
fQkgEo4Z+0WdyyjKBBB0qB61mBoKFCa/WovrjmRld/1ysYNHfmSBXiWg4//Hu1d2
XeA1POXIxtJpg0OfGGVc1EZvqTtJ05wz+baDDk0B0GOnwdf55LA1OOmXvG7gFEAv
e8F+bYztldq6z5YuqkVDaLaGe+z35i9EjbmpsIim+27YNWn4xGmqK+FFM22692K6
xKYys4fYNV8uDH6bKrJdLOI5bYTWrtN/Ii3CzVreEeg9LCFWL/C5Nkl68JcgjK9y
W9Tb4GkXnlo6CIthFXkJenosALZbQgSQMYCSf9385jJaIKUJnRas5ldzis2R6Fyg
93MRT87dM0GkE/NAmETof3EQ2yoj59Zepp36zY7XKNOdozQSiKDgsV3LwPM5VG/3
CKSbraqNWZ+PBSYE0bjy4ygdI/6VH+MDKWKH3ME64DAb7yYHO2Dxl54ZxT1x5Vmw
5PiNmAvYH1kwp3rVFYv0Tf/i4nBxvL/Yv71eqGV/WTIi76JFhf7djsLrYoNZRlXw
FVr2g8+zo5Kl7AGLWz0fK+a8ANcrtevuKH12yrLzEZely1fH9u59GIizXKSopyY5
HPqxbzJvjXJd2kYlrWFXCyUmnwlBqotc3ivwEyEDNt7+/ASt3+eMyfuo4PqHApeI
/MBJPPIBhmwic27/SAeOczGkcZ4HILPKlv4JdiTfNWMJYtk6gaQ9ga4kP/ceOFKU
TFv5GnFFBaocOcVZ/QMZF5B+19lCUB0qdgKDqBEmTj0/zpbv3OoU8WZtbJPToJm8
nWAZIzWRvAuQ6a1MSuA6uaqelAruPtf2ZLd/UyOdMtlIZd1I/wxcJq5eoenSsp9B
jquxKdamz32riiqEi8MK3zrNhfItSV9ELBu7zyQ+D4egCGxO2LYL+GOZELdMCsX5
zqpC7RDHbMLj9EsqKxVSsJob6VnDdc5tcwuehThbc/bodbG9NtFsZHDADBrq019H
Nyv/1sTMIPQ8TM1DANka5NxZPhOWlze263alBIFaDtb8lEHoiewk44LXlpjzPz4s
5FDMHFiFtpTGvO1A54W4mLKHyk76futdQ+8jUajQR2KLq2nQjzI9CXXgcOeATVne
dCj1SWUgxGSBYBOM5VotPENR+W15yFvlslJdGH+uKIw4CRNyREVil33gGZoT1nq/
D4GFPgb81C9xe4L6HU+1beq//ohx9L42tEJrk5rzbksvmha6JnBIRgA5L0sO94d5
R9qkUVKUGGUpDC2+SbWQMxf9sDCKzjQ5+Xe+W63M0ccE2nBrGbHRyePKv0m+qLx0
QxJUYKL5/8/0c9kxnuhgDtg/YNNffHjXhNdeVYak5G8wg0/zGT1ng0AiPQUNR0Hj
P4VRmxqhP+CEKqu899uXPMrdnMBJAOySH4+fgAJfm/HxM3r4zXavjQT+deprgZU/
NUslU0N88qkkIILPRx3L08K3dSiwdLpe83ZiG2WV6eGsS5XwsTWRvP2HOYb4z+Q6
iZX32RhfDFqJGZnaQZSGnA38P7AGQ7u0qg9cseF8yApsAcpqNUEu5mpFolD7/IPg
6/kFUEQ5+ImQC0+iod9gPmExNchCrO3q/yhQlBEJZee9GMVYkVdihEeEBmOqOh9o
vV1N/Ky2eWVbiTOu8QIfaFQBzSKsSbEFEVXiCqh1iLrBq+6RMzpVyVo/Ghkpt3Fb
viTf4jAy+HnMf9XUD+6eckFYJ1R9jDMIijkKjZS98UyhGfFQoQBl0YPuAebN7G/R
U0V8GeALImCcY9S7ErZB0aJi5mMKqHc/hYCLmIwrFEZ890jriWy9juckjiL5jbF8
TDPA6P+BGVF7d6trhT/s7+UFnLOyaZwfcyCxwo63mf0bnFW84jyA/dtlkTdKVSZi
bxbNiIgcSc6Io0bfQnijtge5+Co46hTuld3XsPI7Kd5Ontop46y1ou3xVOpt0x6C
s6eUe+Igv058Fowoo3A0Tclra0Vogi+paUeonvPWtdkR9bQMnV21ej9lu+x4MMcr
/g9nZ0K2GXxPAskk1ry61KYzt3ztAodfW4fdDuCZ5eKMiYpmgETB9xtwaD/eYDCS
h1IYaLdzeaSmiqgMfJv/j+0YyiUp088BPJ931R7gRjFxoOEw6EOfAmJ4ZQvpc3wC
a8M9d+nZHsDRI6UCnkljz6HwEdM+Y56DtjNK0/wIe0TZYgzZjrGW5zSBvxaJz/WB
/8s3q7ah7i9Cgqt4hWDjFS8mT0Lq9pLM5Q4fGkI0y508WYKMCyLWHbS3S77h7YLW
q8NS+/1idkMVneOvym2roqVtr5BNamJgGGLrlyI9j6St0b0DvWJYCbWv4XXcZyxR
7HsCUmotMQywCF0FnIJe/tsafdjD9HVN31shoET+PuKbarCw6JvPOgFV/qYdo9f6
/VyLEW2S361erctCJj/jbDFultJndHWG6Ipj80ju3soA3YprDm3dtmRIZF59r1n8
WvqlUGTYnSFm0hz2lGOkxMziql5VH6k5T0JSnMKA87Apwu+YW9jvIKeQ4/3oz1YP
w17N+ewHqpMvHBas9gR1ai2ajkCxrIgwX9YA7X1gfIIoq8OJA45zYfbv+QTAhmko
rfmw+HsP3Y+zPM+ObEcYSRZWbHd+l4PaCNGmCI/XaNxq6asHUwS7DBSaZMpfSt0O
Y1Ks2sjonGrdQAOJJyc1mb8YUtfV+KovLl1gCOX48ff67BOWiWjje2fxYOGXAbKU
wpn5ek32gLJYrKMklkBRyqtR3sVNA8ccSnQLrukCOIoqiqx32NlOcuh/GdJxyk/K
sOlsZpsS24NIBvKbMKIF4hiYV6pGRlfv/sJYsRWMO/bRZmD9c8/Pnh53XUuDsom5
HXSO0hyPUInYzHGVNQ4hTZilycx5+/0o2JO973O3HU4J2PdefLRZOoxFgkmDuJNa
TF/AlG7iPj8CzRMdQ498B2/GPpna+wi34VOLg8YhJxXDRZAQQwGgxcMzmW+hfzL4
HhseAhJZI+/mkjbEBCvVd9ZuIm/b6zZkgB/VVmYS5jLeHMih7Ke/6uKhygOJnCCU
sSPPCn9DFmQm3fdSHtuGXEwFUIDcjDAz3+2KGYwve9ZgcSaJljw/BcXONCEatbwF
b1L9sj428HQJVIo9D+C5+ZxKXmYbCqhl28Pb3nPVatgZcHFQE+LUKSuZSenzxDRv
CBzo9EGeUrsXxtWht/xVx9XnZWsZeqpasDRHjY8TP6iltYCqABfGkYG0HqFvQVdZ
Aiipi05cpiHPnNfsRKPP3C6BMVqlXndfAPAGIO9nzur53shNrHLEs3hKXb9XWZ0c
ac73/tfK0TO58+lTI8ujW7l6VYNj1YuIwEYEtHHq3n4sfH0UL2CGA3AZ1gRSfoyZ
60iwhCSGSr5D6YY7VXh/iKOXrisQTnUzGIm66G9lqZ3ZyhCgVqHnj487XjLxwn+O
shunU8WSI5IRT2ykXsQT5gu1fcjNpNgd06AwLqhfRdbV8B/dlbMaecSiOLW3kNGK
o4jC/8i57tbmBbFdZ3xzMeU/B3S6SGWhpChEDB/l0ti/4POExhlPrABP3uNbG4mb
iyk6r0hTJPGRFNVcSRgPgJjzABKmwdGNnyvNOMEJ87D6ADgmMnehajnf6BRQeCLn
7I6QOm5agp4nLPM9LWKtT9tigwjav36xzleE0RomNn5z0sYoBQi50a3MnR6kJPQI
TNXtYDAD494+Pu9gXggMBbEnSQM3HA6Et0sS8xSrgh0CNiWXjaubgwqEBED7y6qy
5Y8f9uYs3JVwmJZnuimTgaUsBS1VIg9yGLeMMMsxrpElBJZchGUg0hcupV0y9pqx
9IwZOBEtQ+OecZMl2HVe8xMIE7PKSR7tpeIvPEdgEwJ/gXGu/RLK6KXaFmj99VQE
3GZ60qI9h4U/8F17KPTnfQ5fRDkyLWKSx3RvdhdMvw9UlA7Bi0qR0yXI3iNoiMc1
NgQomEotrk+rtHYmG7PAu3whoTzAosB/colpI0/OeUgLFsw9yU75722JRRfbLW3j
Brfm1qqWvsfVZRu3lmpW7FTnvcauiuZR0PE6MmBFs+htcUskWDEfCcEcPOPXYwVA
b5vJiWNQMguCXGurLqTKaWpxyHq/1uUN6wlTwmqFMDnyj7N7ry+bQnOM6G19cl15
FGKIDxEW6kWd2eHzpa5Gq7I5ydM6Jd+0tUwf6O00hsIZVMiL+0+ouHe7BsLx0d3x
fKYwoJDRDVC2PmhVqkZoJi2ivvLHZ2yIU7USDhJPWRADYOfQ1JP+fZBqT8/6E5wW
ICeJELTQot7ofS79VtibiPXXEv3mb8tGpHD7+ZTNhIAIiX7dQKRO69Kpule4rnAh
InwOcTPo2dQ4T7sSbNQ6HDDR0tAMBJmCI1FiG5JXBhi/XaxT532/TD7f2jGPj4b8
u/EvGUqRg13mlgAQKK0Jgz0qrd6lNmyG/L4+6GKzYkVQwPRkIK4ShL0XwKHITVGR
kISOlyEcShLn7QaXznZrQvRnKz2l/9sdkVYJUHZpwIXgcDIfdmfaeODHXb9TlGfB
C240qdIV2C2N4TtXcas+94UCVOieBUFtxxOp9fJs585APs2dQuMc/HTXYnjAsafz
e6TcGcKq8QkAZpc2NSDdo52magRUHaYwh669kkSTShlG/pVLVi03cYG3rEZNqg/i
fP6I4CgYdTzA5JjJQ4eK/Aq671UsZE3QcMFMIiLxEoALR1F3B2GoOqalNuGkw5zo
NZj7UJ8soyOabp95ICKB2CTDB0QDE/YCfQPOAVVW+opapLU7kRzrXm3991vntKk0
dWDaAr+LY4sU0rCY10t3eDOVcUzG0UVyTUKDfwKmCmeuPO3p8b/sY8d/ygU4Yzlu
1fsrR5bqsSBYTsW68PzkIarND6F0JIp1uZCMU/Q9gtQZmXFRY5CodS2PhRiMJCXh
fjsCQAcwQDVWiHmqqBkdOtjG8kXDKk75jMeeRBnbROXgaj9kh8CIkl8yUwvxWDh0
qPrbh4OibQf2r05T3E6t3Ti44ZpmyIu0HvR+N9SyHeYp+kNyipHcQ2EfFm1GF634
fvI/d9F5IK4bN/qRpmvmfT3gJXC9+W/SVrUxCf4KAKi1+OqJFP2nvuRoczxlvQA1
BODPtt6xkodKMQcAh69zI2Qon1GFcEF+cjU8VQiAKnFNmb7CziwyLYtRk56US5b4
kurfRbpVau/ge89IYd/Rz7v6AezOBBul/iqZZdCtx9A0LkDxPYq3qSwwByNls5gc
p4NsOsYCyi/B+i1P/n0B3BbvB3QtlmZX6ZRcCfGUUG7wk+6RNIb0g/CFQYcCd4eJ
naraMG2oCMfZq6hfc/XQTUxtdDdflhQUJ5BMJVzKRijrXCbDeI16zDAVtw1+wdNT
6W++CDqIjnGVpDzPt09DsmmKwTQryYfC8uuflU4cpx55XKNZlgzDaQeKUoXmQ2V7
4Ke3gw6Hxi/WclYQecQOFhyyftHBlA2MN+zVcIisCMiC4ValoG/91ggohdCXWrDJ
f50La8pYydyJ7dSTS1G4SJEEWWbgMrQURJpLrjo9TP6U3D4Y1nKhFOIZUTZ3Z4BF
8PBCKz4BbycRpwSMsnEsmcKDFGPnqcbQhAdsQoOJljSwxzhGsQZxP7HIRClMjCQv
mOwdhlRF0aNVWilOXEtjJPZ/kJRCt1B3RkjVpUP1Mkd1FKkAah22hvvlZCFtcm80
y1CRKW11eszOjQfoIwOGn6/IatKJRckHPLQfbwAHZQYPr/bhx4x4s1DoSBLwmqi6
Jrwn4oM+EzXwrRLAr5xb+wQ8MaspCJI8qMrhILh6PEpbXrPFkXP85jziJQZr3NGH
weFKpJIQ0McmkkWZbpkM9qzwa7v1b9WHbCUN+KOVRbhGS35JKOclmf/7rUwbaygN
RZ4Uk6De6OlqJYUvbcKwtikkeaGQXbwcs1Ahj8tfZCAiwmjvTWb0FhDbYuls7LcY
7g204HEnZsJnIMrL9Qa1J3LmVvcCSJtFwgeKVsViGd3DhMDq2kZPUHraXns4vhmD
J4kzS517hgNrUt+sPxrmMyLGy+pa/SDSdMyUn19UTtMSJcwJv5WYPB7IGqlVvnLr
oOVIKVLmu61RPn9//wcnASJiVV14EZIOsmcYCgTCbL7c2+CIi54B1SP2qOmHNHLx
PDSJTw+WGldIWM0T9KCWivmlzwmdEDx6ultWN6PlaadcPA/IaRHHGKH4+1jn1PfA
cWR4daExtA6RmUqD7IK+a7U1Y49/SGuM86qxyHZKwpEvF5zAHq8by1bCdykQ+AAw
Vg3oHYK6LlFQlChiElDO8nMeq2ePVZH3ny3Bq7szxvv+wIONM4sK4VzC6h50T3WM
rLLodN2m8axdQUdf9gn9+Om+e73ikXqbkuPCxh1PnZAt9shYs/vbvbI1v7u+oHka
mpTfViEGQ3ysutpCoicpNKCxbiwa5eL9Bgj4627i12Ow59tNXKf0HS/6LRCKiEhm
O3ibVAb3xDagfwXQAxOT+ZrtPPDeJB8f5MaL2jFHscEfZKJbVOYgXjv4L18d0b8d
gDzouRw6sSCtjhsuSJfxBGqPSN4OwCz/vWUn9hp5RC7pAEiluH2H9X6WKuvW6fOc
0bskPRkAfKRwfVkUjMoCE+M0ggOrLVl3HVNnYoGRS+UZkMo/DMiOvpUmjG139Jt/
nK7DwNdRjq/iq2uetkT+eFRjcLKuUwkJs2TZhjhzTTaL7wgv3plCucipqrYu3G8v
syKI7Sgc1C66gKrb8Xit+rv6VFcjbySKfR3tD8+1VXV/ipoNjwN0LsVncoSO8Ktb
b0LKK+f8PFUDFVWku7rwQwJhHdwnCgJJ/aMH6ClgSo7zSr3x0bb+L3DWl7k/j0/2
qXPa3yen0Simvec5BE4NWX7rt0e8yMZjAx3FbnfQcew8VRKAXAiw2Q1lZV0yWcG3
PJvi5jgDLSVlFkoqcJFm9cr1uwpBCjXVYTpY1sqXll3cWOkz5PFocQCgbnJ5gjq6
Mmazwjlu2mMDEDhG3JtHvulO1UUsEN86goYn3znsBMP5DIVFc9F3Z9h4Nry4wSLZ
hWuwwY5BvTVTt8waRwowm1xTv9ApV6Z7MbwTHfsxIrJsfGm3xB4Z8Cro9NW+VvL/
xzlhEtnEXYJsyfVoIMBljrrAuaHnRtb0tJiVDgcdEvTWj4QoyC508ewd544zDbI5
5bkzwu5e0MOsH32dREDA2PTvswP8kU/4HsfvD7vbZBK4Vc/9XPVvSeLMydVuvhgr
fIlb830CUHFCCzhNWhjsP6TNDwkLLejaVsRAcMqlLsfCqTOGdTbXSqzv0lmbwHG/
d29gYMborPJecKl6nyJVgOm+qI1djBnmCMV32yb2K9TFv6LV9Ipb1b+hzu3ELQPN
GpzgVU1m8Y5leyiXyZRuAKKnN3OdU4TvosYHZ6meC1glpad1p+t43FA1elmy4vK6
DHYV0DRazB7RZV+3xRmk98KPiP15evy6MMBGiLjM9GGL88iOQbTdsG2a6KDMHUzt
4wasBwOLBmRjd21W9utuvt/rfluq7Mip1app7wBu3PShji0CmX75zfCT42JQ2MBi
ft/s6j41ERQtuRC3Wg3nlelA+iNF/UdoZRoYM2SyIh36iJZKQq0tSHkWlwJV9P2D
extQfjRsousuh8ERxsUk0kSRr9RFNCkFDrQ4o7h6/psYHnuqbh8DdYvvzXUalg6u
/f4xIuHIxhBhyLea2ZavP8EPfrGKiICAq5QkIIoQunFJHDTk4KXZmVxnLDYDK6K3
gsKxRNKpalT1IaNe6EH591yiO1QKFaV35nY0h92ADcVaC0pyTTw2jagJNk1tuc54
IguHhX+q+Gasy73ljBny5uOgi/ECdrheLn5AkYWULHme8PZtASewA6qiNq2l8JE5
nyHydj8xOAw04m+AbAINeGTJcjzWZhi0bSZYC/IsPAs9e1bsIOZXBxA0Cno9hdyq
oUiVgCu+YTeQDrq28/dKjfPASbcejZgweDDDOjdPBFAVF6XgJZ44PVbHAtEau46u
4VIF5wbEF4ubq8ruhHrRkWTfmDW/RGwuVPOhSnaaj+bXGLONpriNqjfw1mNbwmK+
AyeG4a8+5Z5hNjHgZLMbicIZx8GuZvhFOUuzB6UxIVbc0j0NLiZTP+/lNsmB2Lnd
QUhU2qIBFjgJYML45orkRYlWAs9BHEbNX1euIH5hxY05OpPOL20lRxWrGUH8PJG1
ouo9pzGjgF7j+2QKvSz/iz549cjXoZB8p21fRAT0oPlZKqqXHqfaoIUvEzmT/Se7
4pK91qRqjicKjjM88zqp5kx+oA/SqGz2U+BCQMKIbWPyxXDjoZe89ZR/H2IQv2Zg
hdqLFKuMPk6hWdYx22qGWL+ze+xjaaPy1fzCRIfFp8XqZ+MEBnfJuaA2DM9CsdWO
cV+C9sa7rZ4VP9M69UeJanGPgfJ2/xDeSq527hKOFPZjFGrJf4b95cv0HJ0fP0Wy
Qn6lxTWxRSu9vl2RpQDTn4fcVo5K4+fEUo/zfMrI+nni0PWOwM1MvFtUn8FNEOq3
1bSMEdVvK+wAK40uETLHfi8h7vI8SU497tkOp6vFog72lVh14moLYfP6OzutA7G2
prSxUmJCbbN5iw4qTg1ai6x2EOKBWOBAjFb/dxMm9MHiT0AT268nBmu/KBWD5Aaf
Ntzdf1cOK4cEhDBM7N8LGy+XYITwvhlyTON/Gsew7RfhPa7eDFAK+7dvUzwGtsV6
kSFOAv+MWsrthgRJCIhMuC74Y+Iwo3+n0fsdAHvXbBdVlG7JNafrCTtbGd14mcEs
ex0hGGFd9ZzQ7seLdWz9c278e+sgX+n/akZ1nDv5/EdHnRSJ7/keR2lCSENKkJA6
gh8bzLvK7dIpwTu3+4IoC0cLCT+LDH2892OI7QBOM+YjjCJdhUu2zLW6nFGRGASN
/jyXIs8/qram4bsZ5Fs2W6E/a2bljLLo0IHatmt536TlynAahFBr4AmIJDmpvRfz
m719c2Epc74ls3ccdhgRcB27jHF3X3A0fM8wr7SgTl4MFDL+KGlQfcLIJaB+dHoI
Ny2v153zBzWCQRKroy0tFqlFZT3ROpymHeQNTSqfPOYKW5O/mSwU059AwTTyxhSq
VCS2v7E6fMkbLGTLcVOV03Vdl3kMoOCbdXEZaT9dZ9rQGkf17ExET+n7owlguWbJ
Mz09VATyhEKo72le/B45Lq/QewNykEiDUoHfR4bzEyrZupG2k54VqhGHlafRc+Pl
nhO3t2FvYXOM0sxDMHaDZmusxb/bJSuz2xQ9iJKirwXcPufBM4i4Qvy51J3wDRC8
G5HVoGb/YvW2TMR6ou/B2Y/l9un59v7FdDin1IhCfe30/gMca3KJc+/uIJaa932C
uTjefY0IQtscm+t9vqx2s1Wi8bRaXwjGBXsjdfeBl78YBWfhDmswFgwdXfn/8hIx
0fRhjQLmJbrmpXG6BCUqRfWIUwfFG0/Mw4NeAkjXf29mnVyk0rfaezcwgNVAbCFC
WV4pQ5JaTGps+QRX6YU3CIptrP1k2YMNXsWCaosTjMaQ9IUMfQBQFCHeW2+Q71nV
FW0BSPKIPUsZHu0L4FCJ8+YaaZfmg15otHOWinwVuBelHbHvb4j3xGFxgheec1/i
utL6/CZIgJ86vMcPuOnJcTE62eAei4sDfXHSnpmFlMAJ7ksy72WGb8DV1opIJhfU
9l7dNf7nSIxoRn1pIXcup3rydYBPAdut5lkhQYei49NGeH//QjLaBjVMASL4d5lO
er9tVdbFMVYKpiFLnXU4CG1zg2pQs4nXWFa9DugLvZcLpw9rHw7SCltKw+OaRTQh
Ek54RnRhPsLPnmxrYgUAkshilNBIEqYSaA1ZTMXqmIzTLBWtkRAcuBmcyQXp6tZT
jA+hpRxD3/U8pVjwznF9rBiLJ3Yz7OrKWiWys/BBNwybKNPRTdHQdBRqVIeg7+vl
H1upA/IBYjy3rmEGcg0D/YJg0sEfW9x7ELaKZs/62pqZ9VERvm5rfubNv+NwlBuV
Or+yJKSX9HKtBZoNPMzt90uTWNqghtOCxlq/9OUwlDOuyjpF6Lnp0DDBVuixAVls
yI1qW9XWZGkT8e3/XLRcHxvSIg94VwcayJZGXrBmAu68jHUxxJ7CZhVO5avO7sHx
d2vAEck8gcdcsPzHry6XS21U04jiUO1KX4pA4EaSaCExCfBGT1XVywi1u13Wbl67
2AlYaiWZwDMc7ouWUZY7LtR+pFzePYr/s1U/zTJgcoCDQ1ghXoEWNCaTeiELnUpS
KzEHn6SRYkg8Qese0gytJKMKg4JtUimW9zD0jp2EDXbtKosvRV/z6jJfqQf882CW
AS7cDhiDJ7nwuHvxzd+b3Vtk+OoWgu71P+O7SP9nBivtWBQrq9Q9YtzAfgdu9S36
6L7U7H2LlI7uLsYVIAA3BAf+X36JRf2MyYaKEM1TEiVDkw3v5lWLbfdgQ2cBPkPR
HJO0+eqLFvPJn6o+XopsA2MoogwdUCWuOMmfhuCUfSSIuXJF2CLOVUTzYxhCWVgE
L9npQZAqbzSVmg52+CQatFMNE26p9aKUhGu5hdvrMO6P8BBTWWczJwh86Yb145oP
dEX6kzt2t10hv8685S9yxli+FHBsChR23Lw0pq9+1hVthITtbacp6yqPW66rwG3P
TXJJlNLRo+q9uYcRy74F3a5JnVZDMGt1sZVdI9h+265vuQLSq8yhCBQ6H9iTrBmv
FtVq7yzpiaH+XgfE5lGc5nfyyoClNw0xJb5J24oPtwNQ+9UM5iIIvjOxHiomBKEr
WuHM9JVOYQOHHvZlxqbu+o2pmxk0ScZU2pKBOZ+Qh+ifLLnRmrCMwEAA2U4RtNvf
duac20OfcbqP54OojvKpSAeQL9c9y63u0UgarbIAJz1rAoAixvjDIhujJ1aE98bY
AyKKxq95V9Yi3Hz8gqgUZZfleRcSHqJObfWOCzXUwHtg49GaQSlsYkE3y5b9oSbm
fmJqGPOaJxajvQiC+BEUvP5gNhLEg6GK7dImbyItD0KECJcgvjRVtYPFFXcLfjZH
97CX23f9KffBelgtlTsRgZDUW4UG8IIYEp/vMmTVlIn1Vpg1HCRLFmGDXen0RRVg
0llzuQjHN+m4kIuZUm86iITmgEfVCZUSBOgdQ+i1FDxrJ0XwHrgyThlT9q8W/p8+
6E1iYPB5dIPRe2Q7jVkbyPA+P2w+G7wzoJKfI1wnnpX7ZpDR5ZDR23WeHsaVNzzu
AuW5LOBUcv1T0icAni9GJ2tmfslg2LeJcljZdJEh4z3RT1LFZH2DKxAZEg1xU8tw
bi2HrB/BeWVXcSDFdsf3vw8y5KJXH9y2w5IAzYgCwYFVMKgYq9ZcK+TRHrb25XnM
+bHdMHrVvVz6tZUcP4JeUSIRmQC99YuPz4UiM5FG0UhX7WVTa9RsFw++YTY7BDnI
YvqYrxh14FU/pNbbv3Wqw/FXPLiHe55pEP1JixeL2PSdqimDCQNksRPzvjCzFcn4
XQfu1MZiC+SGCLCWM+4eMO/TH/I2O2sUuGLiafO5Jc0DI+SotelJlJXnJ80Akfbn
+m/k5C68WUccpirTgKxGIRdg6ysxn/PEdWUzCOiqMjy7Xhr1VuEBMleZdM/gwZEP
/AFPcexYAmOpo///JUupdIZmGpfuQzkg7Og0ImBq+dmjKoMCYPthH75ugt2ZRCw1
GsGo/B0V06SIfOuhgWieIUGNLse0yoXU4Ua7ieFdy6NKv32L7NX85GbzubKVxXT9
QDIsAD2UqmnKvbSG0l8hVx+BmpcB/IssJl/EHpopgI3dtIHGXvPB4sygF1kD2lLD
bgfNKIPTReJl4LKLxVFHV+DOs+XNBOdfD9jC4POIdtb3ax+RvrfL1M9pbYAIPHHH
MdoSQ1F1bjAwPPY3xQtO4ksBKD/w6NaeLnRmzr3pmD1oJphxRxDjywfWIuQjVyWB
tkdeWqpY5sFpPdJZ6/jz2qDyzwsEP0GYSxPqbD6hPYMJJeo8VDyZ8lGL3gdL4Udn
XsvOTLgRolFTGMAoHIP77KJ8ggV/WgEALPDijREM82FtL54SKkrlIjJs7tQ+GCNV
G37EXUNBshOQm76FAjF1AeHUGN48qojXy1sPpwLfQHJ4DbBqqKrJRatyMaRU75FR
tRfH114TP1odO0aAGp3jGscG3FFQEneTN3ISkSERQhL8gwCwijCwZ1gQEQk/Gr/r
NH4ib1bm/fxRLp+BiK1Z2TApOfNF6paI0adoOjTdBhTocW7V5xos8buV0/ymalMU
jsRXQudACGKcwjeHQNFjHG6lptGMHP/r280RtoZt1wM1Z7kkEhtBQCrbaia8nH4o
9rj5wdMfbQU24FxC0SYz9YJ6gLxZRJcU4L0dscuwhCWR6duPHK2pGWirVgE+hJ19
B2yn40oNsj/F+BDndQ/1L5mxHewtOHn8vTalsJz1xsynWB3UQLWsubk0mwSaaVjK
Ox/sSuWSDi6X08vfHsftg8yADNN8eh+sdw/WXSgH8dBViG1Ge43ISX8WkeGRHzfg
wuk+LsGbQi0POKlHY0U3fTKph9MRCJBM5nOyuwY8d4IUBrFEmvh+75/TbITA0tCm
Ymr8hxEeNUziTLEROblOLow3EcYehWTD91brpmxrh4Abdwc5W9CdnaNf+Q7kAt6p
P62H2XTnZd8nEMZ0P8/RvQ==
`protect end_protected