`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
Qrmw3cMzxQM1gA1lJQe4wVSGrYf0d54jFJ22FbCWUJif+ckm6nlPGOV7jO+cbAd4
R3OQO+MCJOgPkSEofXZXlpt1cnpEM0X6vEuZCZA5kOVBEf8bfg4QE2PxS8GDJGVi
pglCLfk2fS2CrImbtVu1acfcZ8R9qLhFWYTodNbQeFDy2L8Pi9hXenmAMDhpD+E5
8NElmoejMg7Ptie8waN0ZPuWr7jnzdx3LvcD3q6nZtPXa4fu2WS8MJgZM3+3srMH
lGJQ9KlieElTfKfUoZ9PJFm0eDyMfWbD5SYNcBhl2GOW/jW50cixET1X2lct3jfM
6Y5Vg15OmlItTlYJgwZ+eoHxo2viUJA0CsOusLqfkUObmjKAQpTjZROlokktY5CY
SbltmVUysG4TVz9vqMVWMkSzHM//jtvrfGrg9RyYJKaTWpPI4eanvlDKPDQHYSAJ
RMdJ/wMApPI3Qv2skwBJQY94HKtyFs7cfTZYe6P6WO8Ji5CmQoR+vJ6ze8o+AIoJ
JLYxl4LcjnlCOxwoUDXhGFaW7FoGAPrCuaE5+yxWc9iKhixPyfjzZalN+ewO7cni
LyVAVfT+z579NXQg+awzHYdqeGYQu4s7dSIcyZA5CSSbaoxhBH5fJe0/YilNWq9a
9hDdfGM147SIA3K9DX/kF1Na+NiAmzFN5wsNXkbsbkpQWgiSCBHzRj+IzkXSZABj
0QDsu0f270Dn8nQEAlnOWeTIgYJcslde7JrmZkfoLdsr8/YagE/XP3st0IbQG7bu
pCYTuUGAqNoqTRK5/4KCyQRaXZyhj3reW4D14YnPjRA+FfTrtQ02j6qhSri62HWO
JkHx8MPlyHzl8FsEtq5ZIzhDlMVLhPBBGEO35SG1HhyqT00UmMnzL1OJ5R9JDzBW
nruDWU5H5Ef0EEaKa/vq/vozKI87DBHDusNLicf0oBMinahE5iboD4l8GPl1FaQn
Pzs7lzePiooYu6T+8fMV3wf475FjNAV6x18FwJazuw5GRqKNrnTogoC0q/EWJW+O
2RP3bTstLE6KqPiO+uvP8c35i4cnKeLhjFtUTf4G2xu3iTT/Hm/IE6+XOt+33pwW
l44+atJPYdf+RIMFCPY15QGdPrkSCtKKFeyV9fJN8+kjcA8EZTPtMlqu1LRQhQqE
pfPcu1YdjquWWDiu1Las+O5w8MPxYRM0eHmS1QijTOseAHP6RNDRQtTzJOmJvLHX
p/fyyFfJKxve3XA0EK3GGbios8nQM/rPUJrCujv1SwtUwkf7PP7URTrij0GVfS5t
t/brKa2hxGrYLMdnxZMbvnurHifpSK19kTz8bGiFVv5eZ5eOp2kKuVFlpJJHhvjt
hTNMiol6q9Xj5spBNYCvG/HgJLSAzID5xGmy1B5zUOnlWDB1t1KolRi187xjzdil
qgO3Z91O4HkoCesB6o9LMNIq8v+J0uJy6moV33dUuO2NdQum110JxWf36kfRcrTD
q+bjhwltRYlUhx/1AdO5v65PscoxX7GKc7mZgeYTpv/8ioVhqiuFE3+Z3O1UBE6P
DJb5JxWswsGFsL7M6qbEkGorCZfhpgJIChfgmGiqss1+ygZZv1ygFK/yEjUulsq6
kK3ABVkYHs0hJ8bY2L85BbyCoxbiYfjHRKcp/PIP1bZnZgHu8fL97Za7wdUIMeR3
34PjKRNFM+A+mvr/GrkPDCsLiECj1ScI52euIsTgWhKxm9ghxrz8Bno2JxnFSZJ9
s5RcYyab6vq3SBzhK8orlB3CD8tsd2i73sJq2XWUJZuUcD4OtHnlnCDHtQx0ZZzu
OqeJ+to/qsHKVWO66cA3NdFM+kb/msCb2PjCAwqwqfEQwqiEY9j+z5ym3KGUOFuZ
i6tJeqdOS5L6DADdNILH8xpCEDwp+wyOVKMgE9nXlXIqcXVxesTEU7h3WF3rRnNf
aQeYWJ36XyUIdiAJNQ+5eMu4sTirGVu67fLM1bQKwRwVNWGBZloiDfm9HGC8JyJO
DSX5PPSGzDE0FpU9Inim8Xz9AHOgiyviLiGdnMHkTbVtK83DIegTT5Nzh8foZFgz
yJ0UNoXfW7HF0E0EEhu3itOu9rJaVZ5Bi8Ru8jGWJ8A5NqCsXHlCHKMJPziV21V6
edj7Y2X9grqomIpCrbbTteqCN72w0vaKKRHh5lSi2bfLV/8UUfCZOKzTpGWn3XDr
YXFLi267trCpv1b2SdLsMUctjIhQI+hvDtPk6zV2PzS10v/oldayEXw7VP6AUdXe
BSFHZveIHHXUavjBjWsfqssRY7nPPSD0G4kI6SzpYYrd69BNZRWgqluH4kHvqKkr
4a4+fDTrdta/E5aXPQdQWuxEjTMpd6c22BQGHpF8V8BuXMvTSnnTxU2Ejjh5jKn+
FEfxteesNRMnQ5ZuH7pXJrRywAZcMOPEcf66UOdhSI9epxTGYQPiCR+EjavssrPG
CFZ8EiQTeYJQnqZKpNVMQVWx/hHwPY+LeByC6kdTFj5nOmHVqke661qj5Y+vEzH8
gT1NSAYlem6CD7v1L/Aa3KEJaqtc1HJGijxq3Y8U9m/gw/iT/lCv5+d0gvwGF4Tq
n+Dz4Vqpi2pRkkZ9vYGm8SQwJ1rxmXsBkNFHGzDfeVXNduZA7wWYDRjiHeQpapSB
JAGQQLPiZr7XtaXXoHUcFsczHOynRGNqah655phYBCUurh2ih/JfzZK0FOPs1VMq
u6nVE9vTyO4+I6aOYm5WN08yUy2Wh/BjVXq3lnLaFlcJ0hdWLWmAcq0dNE5SaM2o
Gb4GuFmMwmZWqxfdr9HWROzZWsxuvHDSeroqi0x7OkqKAS06oD5uLrf6xgG0ofWg
Ie8IxB2/Broz9bVo9x5QB6XGDw9A2qmeIQwFo92V354cLUjUwqT7AVv6WgGvbzmD
xzqyRIwoU69+UWQH9HROemINFHEH5r5j+s8r/YiNCuploSaavYPKPCatw1F33Ay0
4IJ7MvSSbaBwkF6Qq5MbvIyos6b+iKF1D0B1awlyzp7MO8K7S8eZSASasMm4CzoL
TdzMYPIoBZWWs5I5uqsglqXMYOi7YVgttzVhQiJpEFqOHHm3l/BW0ShvOZD3WtnQ
4E34DrGKZGzyjiWwm5JGO6ejxm8gDAx8h4PD8Vo4+UzKN7vvlIBVePJFBlrOJhH4
93RGIwUkHDPUp49qebCUkJDkYd1vBpqzG+K5hwJk1UewQNwTxPXlchgogEveIGhv
jj8hMQCQc1MSlaORws1kjoLShMmoe1rEYqOR707F3z0Hrkm48gSCwQi9unKDsZCC
DJnNIin21gujGafVPP2ITpf1aXHtYJX2eIYTVyOauDDPqw4VopYxn6gc3hDJ+1Nd
I6xOFdnmJInlHjpxGwqJt1q6WU198W0BUKXnfjpaHHraAIJPojkXKoOALZ/1Y5GB
fUFibvkkrHGd69xFjhdaPTpUGXi4CV8mlSmqFbVqebxmetDqlSgCPKsN9kyFtJPr
WuJSF5/fqLr4LsIBMXTIz/Er2XWExWTN176vKWqXvBTpbxhG13d6X7SJQvGigJjs
d8h2+TN0Is5jax/2kuO4UxQw5FZgSRcXarQM4fNxW2x8MoFI8+dYZovq7qN0PwLv
DH+McpYanz9BKe2KOyIX0KLNe3y2SW+BHre0nNkeP0eiQgTeBi8p21xipZ/e1cgZ
19JaM5xS4YALQes1/pFV8rXs+MUEa3nvkBNsqX3/ZPdGI3ooODi7KueVXEpY2Xp3
9TnUbtl9OUX6pUg0UHitT7qoXGh6/a0+9C8KtJPv1BFPnYV7Hg8CABpjsKqeRvCR
vSU1oDvsGarL+U07X8geZN9598fNQkcjfbx5znFnJbHYtTXkLVZmnSC9c0k2vCn7
6w6tixqmwLBt6pfXvMht6BSnmyM3YInfatrsoogB5j1mOB5GKSwCCUCcUAawFbV0
duJevKD6jbMT9D1HFfH7wU9O7YV7UGTnIrU+L+u5FHzOeQ7WFZTVYNDq2d8HpIl5
7W+bNQ4yUB9uf57wI1yku3cdU78IO2rOzAz+u9Hutg56WMeE7UX2cTAhyzba+HoW
NBKXTc3AamV2P8W+L0w76cb60B79wZBPPCXjHxXZo4/+EnghcS7b1iQNwsO0yKCj
azmLF9Dtt3oU49eEeUgB3R3nuRJfcyn2+xepGYwiKC8BU1KZzYVh5RSCElDyjqH3
NU0rHa0JyXOo/zKXkgGAu8mZuHjFs0eJgyb+Po/uucpAXrstXWtbvY+tWejwD8oW
cPd2DWp9Jp7rqJ5z6QiVdH1+3J3+b6ndtc/wL/RNHUEHD2xX3+q7KoMqobhREWQH
lY/KIQsFngTgKyZSQKd2HFvXuGg6lbdd3QH/p0eOShQyk/UnZVD/l9PFJiUN3HDy
lEajYJtwVjteUChG/GKZKGtUPvVfKYRFSvnMrRmsoYMWDOEowpuktJ9gtulEf2c7
16p6hBBCNIeGp7DjNe3LgAL+j6Uh3fPnvaf5huGJ/KclgLgx4K6Doo1eaRUjRiM8
u6XERbvMOETfyApZnerbY1uiinHhBURdxxho9VPbXtVGTE8rDnmnDJ9u93Ex7UDK
Z7D/7AIzA27o2O/4WAsqOK2oIjsV8VYjbSvBo1+SLj4yPCBPct6Qxaszmkolg8X4
G/tg8gbAxpKrAcSsksp4kVD6PywVuCNL8otxQs+MVhyXym0VQCxX3zoPjAznZViL
ETabLbUvH8B9nm6s8A4hKrgu5HxgQw9ylnWkSwWX4n/Y9YW0hH7lkXL8SKwTsX4H
14G2NFuOBKuZqLov/imLlU/P99JHq7KaOArBgO3FtusqcUHFwAudPpRh7W2agkgX
6GSws+pqxZuXrdWcvexMTevjzMrUGPw0O2DIqQJyPd64oerxT/NtKuLCljywPxiE
eg2B9i0LNWNiIzHWa68VfEaxabu2yuo0ZjaYk4g0FzMFE/HgKL2+N1haD4aer7jE
ApgYJIdaX25qU3JvX2XHPTDjR3g1jBD5VdYQCRFqMlirkj40l0f5H5HbedfYetVP
155VonUsDPqQn41efVRMRNtcjqrUkPmfBN8BMxTL2s1zFi35THyL9Y/CI3xGguOv
iYFgCFWsZvW8zcE3bkH34/oWzI1Kltj+0qQ/h1rTDsUylZoyJFhNN3Rh1Qv0O3vj
Z1p6P18eePIydQ+hs7NnxjtT9C7M9Rh03msphZ+JQsTkeeVPc8hNlYRU1kf+arPV
j9tk5alapKppD9Qggw5U00TjDuIBmsARPYfVpKmF1k6FjpC4bdZC4w7fjlzoUNCj
Iobeg3SS0NrHZe8y/cS+5K/9T68XO1C9H72zyTkpJPa+ozBGaOe1pZSJmxgqd40V
j9q4DA04I1G03yKgXnKhDBsgQdm/zAHltPvUB7j6igHOvy84D5Pg2R5C4wWJNoX5
1s3t9/EiMJ/9TBAZLRIsk/Bvze83hV3qBfkMCNIJB56rECvYSoxE/AObXnwTym0R
4+r8IhhyfF2033gK+0Phrg6ntwnnaduO4kKE74Z/0r4Mf5vh39/zKbJ/j298zw/9
ohgzv4MKeSdrJRKm6Hvr24oaA5GULZuq7AHkmDlMfE8Wrj6asHbTNm8BbGE/ICeV
m6yxKCTVImFwBm1oJQ5flzD71tfGYTlzQg63gCTCL8rp8Mk7ka4wJl/ZjB75Fk7Z
U+JrjZ2rkammp9UokoJzf3ekqgiPwuiyK3SCKFMpOw+OfgebQTIZ9uBjXBBwDGUo
nTRTEBGtNzHF/yyaLCIROSiX6VhaQu/Fb6bjRseh9RKD9aCwE+756y0hf5G7pkFK
HudAkg04Od5V8IYE2bfIZ6iq+yeUtr17Af9ZiJg1KKcga0IOVZe5+P1HVzPQcDCa
+F8oq6FLyfdA2My4Bm66T/JGWgYwGp9YgwKRxg4i3X2iy/bkFiYvpIFOkvyLIfZV
85cflWC0LM7e/IGoU6WstHWLRGsZymiXohtp2pLIYal34k8NQV5wTCl3r5hze3AX
Nq1OgV7EVecflg9uIu08lF2tV0nIE1oo1pDWnlaVNDWvZ4amWv6g02V5rLOt82I9
oj0kFviwShd6w21hEtt9XbNyLgTUbgGZTc1lA2I/Zql6CnM05deJ/18Z7+Ts3c1H
+8v/ny3rXPjth/MZGGrn+V9MVVcQLt8FsfiG3UFxFr+N4npc5OTZTKnZix7c13BY
TfcdJMmmEt5kJ478IERQbOdxw/8JUqAqTBBwoqwXFffz+D0MTDCjKfw88fAwnkgN
kP+qV1v6SDzr1m9PyFTyv187cPTOgeTbRzinzmB9j2/aDndQFvvlQYTYMcHo8dIH
ofRXPu1r1wxs8FCm7AwCQHIuPz9YkGR3J0dSXNh8VJ9kw3QS+/V5BlnABJ7h9WQn
1VqHknTIpyPa5wxXUMxPqq8x0sXbIrPuxjHDEsSeffZRS66/cTn7SMGuSvyfBQzQ
N5KGIBiQaHk2rEmzT+CmGjLVMCL+3jZyn0VIFvUtL8hc9aVKAdWtJ6n1x5sx+qYH
4XMVpUwnVsNygOH1FBNaKKUxEMvph/E6OhnzBYuvf3Rlfhl+taz6VH8jaOqWrv9E
y21Eb/PeTIDTKzD6Rn+fuBBLurJsTgAp3EUsjuRELfFOj2DKEeC3ZtYU4PD9QIQ1
RpvYGbebNjwX4+rnBWONo/yyJM0kFYHzzLcX3uVwIdLYDip9ZUO5H+tQXp/Nky7P
Nb4PqzBb8INmLU9HQpjOWHyizead/W7AIntn2WzdwXA1uSFvkZT8l+1C7zwsE7Q8
Fuigw0PPnO7m7AYRFEvRvo0pPsYCtoDAO7Vqh8mZNmUbKM53BAzWJrwiztQTQ3i4
ADmMPMJB1qfMAnz5VbXUTtefUb2SYSrjzrPXsfWr/8Y6wcP0bP1oCB/aNJiMkMzx
59MTpMPveIzs8yuatTPCvH4vikbu6MUZlXSf51+chxQr3IpEwEkh04DHkupz1wAL
F0AtZG/0X9iscPgfcVQ9EYJmDVPxfCVNpu/MOIP2f3JPxSFAxXk2s4nF/G6dNg0y
LbxvzJipH+jLrz5ELlw84k7J/ErNFE472SSY/Wj9PblZOCkZ511aLIc4AgXUo+wk
QSA2zDdlF/qc7PSUPDMNKSS3296aV6ugJGCuGFAKS/1DORm8TvFJn5ZYy/Ps4JNy
/6u5ZQdd0sus2yh6v7q+RH4gQwbxKvngFN2FQliraIwHvfFQnXeY9VEbNc0zK9Q8
Nsf/eVzzH3sDUwJJSr9nKZsMvgrERZLESvNUVq4nW01RHePxU7LN+8OOfcRvLHhK
4vhEELmsaavxH443jDcDJ4OcnpR9vuLkkqZr2qDRroYbbaTS1nOJP/tb+TERctkA
tWO1tvX4KM2omdH2aMlTrm9DUxU/7vdqeY8MJJj/w1oy+8/H64eMlmFm6Mxv53nH
VaGqGbZPRfSObFgCSxmp9npxqBI1q6Yh6ZhB8D/AXrtaATHsr+8KgdCAlzIO10Pc
EtSTfmjeHB9rIjQWbJufvwTIGCX6cp+Cs8vRM96zBwf/GsV3FXsogQeRKXF9MsS/
4z3bT2lRXY0Ay1ogOUVL97S/iHmIyXoGWsOOQ8gezh35hiW+3OfPpk7rCT2uCE9Z
GoFM8ybinBzUJGTTRo8Gzr2K5lBtZ1Rw/h1+9D+U9nAeEjHkxIrckcuLnrlJVyKc
/7OkaQCSOEpjSSBVStL4d35FpeVkmkxKJjpS8N176WzNeaz58ZJojMrQDPJg+6xk
h0ZVERfmQ29XZwm4CxmG8img3M61pIjCr0DU+oFnJqRWqwCB6qvT0lZwduOgW/Sh
kHqbxfF5CYcWUuAr+TJagNelokLnYJQHiMr4nsgJJmcKZbKq8nQRdaIEWE4Il4vv
4LYOp8LjQ72PXDlUzwpTSd0aYnqv88kb8O/qhfPB82vifKOPYqaIZJ40+FL6NzcO
hI7UXZxs6Z5LTtEhxpsPTUn4kfUMwKmDyaIDD3wo4XI06uw93yV6BXLNpk9350pB
jfnaL7gHyBpcFB9nGhn+wi1ddrQg//qk7hwdF7piIr9RRN0ARTOlplc+lrWS20/+
8iLXUGis4VMtVafwIU09leau6nI2x25iD0yU7ePF46DmIVuy2TaMKgeh2RuH7JYX
6O/BHV39g4/ed6uxBVwR8lldmnhZvpSu0MF3O3AMDzAfQFmdaVkfe1i6+11rn7DW
vwCBtvwLMCgy8E5p3yghiq1Gqs3auVTh/cQBAdynpIAi+Wdh8TcKdgA4nhaKaVzq
E+DhqT8RvlCikLMR0wC+WEjKAeOycEc2tm2DmhPttDsw36bz9urUPXGS1rDhEoBZ
HlPx/vuFIj1xK4gKvrLeuaJPMEsNsKKCpqrOcvalYPS+my1Z0Ark/jXgSmDl+6Eu
5F/krQzr3g+4hPWWqAs/6qGwT2miXNMo2zzFsppEbMnEjSUXHfw46ab606/hLEjr
ywzmjrcSWICrB5kt4t238/M9Hvh49hZZKDyLvO6s1qBjX1CXp30+Q6eT/Yf7TC4P
NDM7+vSWDliOHj6iTYpVEKXYsGATaJUvRvGCuIMkhGWIQjspNhMtaVnn4PhB9eRc
fzRy3CVwID+I4GR0h8OAS9Hw3mGKJmyahTB3I5mhoqOKMwC6f+3Qd6TXHh/gdfWe
OBiqrqXB25A7XdJ47My3jMHmPGJOtdhGsq1gQpuECsLsPIvZQmdojsMtRupF20Cb
zFY+KKSP/4mmg8bgxp9vkNFjsCKsULBP/38NSgCA8jcoFUcKKlePaDBVLWwHVddZ
Mik6+Sj0iCpIzFeccvmEjFH60USWl0xqTx7jagz9ZsdfiORnti/ch7E19X8TQMT0
nawcdRO4pmUqIrnrKXA7TTp4Dhnlgxwt3+U+5KcihvrRyOwyylME/TX6B+o4SXUj
cWCzbTpFnAvZGu1mOGGfZDdKP8aZLkfpbhx+aMvY0UaKi2fy/xxh687QyDInrt1i
neM8kUCDab5Dz7MU9Tl5XFxIQZiy2au5t1rCefc/rJKrmyt0edWUMAHi9qN5gCFo
wGVPEl1GRS2PkVkMjKoLsyT9S6RvA+ETZLGhbJXKIQ48UyhsXY2i+vQ4j87YYc1c
7i8zVAFhliu9dbYeS+cYc11UzNZdxBJibzvfpIOzxyFR+J8ssnv2mmVRRPgYdYd7
Xy9j9RslfMyEJtSmRExssrXWF13d6EBuHsOGrGE0OcWKfyOu0XSEYcqKv/X6fpJ2
Utzx8ngaWvqArELcJ1HbtnDeRAT+LyyXxuudJgWYRiBeqSVwZ3r+kkw5/MyKATkR
NcSo0QfuOTLIKlEF5aiQh69B9ooLc71zLrSLJIJEl2UW0l3CweGq1or/V+VMOg6y
MzdRZyof4YZfCNvPd1nis77DdMIRpTeYT+0nLiDheGxLmTa58/zZo7DIDrFKIBIU
+BSSH8q+ONbpZYycWVvleeeespsOY9Zy+WYD5PTuoRHmG2htICXYoBpeZsjWvYhg
VgVOzjJ6DFldNG+eeQ0dzmd8s7yzO3MOOmaWCJoAk54DW293CRL1CjGz0T4jYgCJ
PCuKuvxsNmANtnhEwbAivu2MqPK2xbx2oMsjbW1D2mrsgg6E8BunQS0mFzyd0fD+
xdkRg06kmqZgdWdXP+dk9gqSvHRiWg/dFU+0xxm6vGJNvL5A3HvstnowuVFzcMHB
StB3J5DdzM1S/dv4hkXOv9gKyXmDwFHFmFSygZyTChpgl6oJEDoGJAozN9jYhGCz
8Xqu3zju8QDQTaCsYF9eRWQdrKEFbsZYpT06lnTjEcz7f5+fGK77oCMFtasFEcJg
CLvXYJf5V4YnT9WOAclBk50VhDeLRdkhX4greaKOVsVrTDf1mtNjBRPFEH3WBAVG
Elok48EZVuRWaziFuoWF6Q/HoRkK4i9q0neNkAbHwv0XgxJn+I6fIQlUKMfClmbK
4irmE8QPL8phI+g4YZuZOXyTBHO3Q2OryW4U1eg+oNnFyWYjKGTGP3pQhecj4V0U
HzwGJTISbOGsU0thDIqsm1Pbb2AkjHWVgvY6hrpjTsJtFifVuX04pRklK3zscNeO
cianjWfUgSgqI31LjhqupnFmAuiTZlt9ao/Yv2S9zJYILrZPW+aaS1rtuV7qcxbv
K1qOn+JAHuTMAEIlgHaKKXK1rEeN16S/C+Y1b0KuVp3ffGF/2iogeDIxIvAsuJfW
FBEY2EoXwqfbUr4a2ggejm8gTGyW+iJoAx+BPuZ0Z2tEjQzFE8FeLvxNPRAnUi3y
YRZwWMM+3HEgjLMsHxiWsFC0xv+RW1rBUCxNf4LGqPRJ8w3sFUKoAWcVO9tPfJFP
+T8dkuaTXeefVMMVpFn8BzNkW1WRkA6kyuoH7K62xfN7zAMqp+sXWuM2Nibp8aJZ
A/p+HRqKgncusKrsFgDuSR0vW+i/a8CaF/2c3SSzdhHxs+avDNPjGyvLM7NYQypL
JlBdH/8kuFgM9o7mUVwIotWBCABdBbSmo9Eaoy3ko/TVROjGjCvZEl4/I03JvY3p
WQyQrunhd7HyPOKvMwRBs6FUUE8R2D3hKxel3fAgGRszkY3UUqM6kAmrrQd3USO2
vwG8dzvADpy44yUPx+vEGvmGUhu2PsipIUYHJYp8gif+SuG51QOVeKiutsZFy+/i
jXbOHh6Z7oasa9xHY7uLuneE9xudSCAex/8u7UksUhoIJwlfIhz9NzUrjNU8SoXs
yNS6rfP6ufGnKYxa6/9VKEZBEwucMz0IGTkkJM2/rK+xqYW44w34CryNESI9ZBxg
oeKD+GaceVJQ5JQH+YTiaV1HYgZPS701RtWQU88ljbpG+SjvrGAoxImRXC7dBuMR
T8bH9MY/aGsWim5zZRSK9Egq9U2fVpScAmtKIN2761dxIT8rgw/9MfYXD71vYveO
VvPe+5IqVeNGl3xl654CUWD/VVuWyG3N2ergU83fsrb4woXAG8+Hd1Zswwl2Jplk
FSIi4z3hJIcqq4qqZdfOjMt6Qe/k6xXkp+J2qxR+peMg+fqGOctZaCLLgy+IQd55
/odae2Da3wOFRriAT1a6/eNwbd3Nj7jqndvJCFzzDlOIF4wjdg17aqewIqHO9cjj
4K8ORmM1PFai7UGThdTjl/q4Lm6sBRphtnn/IieO2au0ILXHawIce+qdFVu2vb2I
r4THukvmpggnudbMKPuwv07xk63jcONrU0NFwNcky2LFQsawWI2bz3mQqZVm4Sdh
8TU8zcjduF+Ym7StnO0Y1O09vnbsenwU0zxwklQRuOqQ1OQKOEE/f3O4M9NERVqd
jTCadt9p3KdvPCtC2haRfvCncNfqFMk6PiwodlZtx3Ezmp1nUsLM7PTfuspXhTwB
PNL6AF4buFJmHoCZFPzYSk7pBLP8C57F1lDSOGHQmlUIBJHc7RwfgtuSoUaxqNfu
BiFbAj5I/jC84Yyhf636BPHDR1hCkrwg8G7CQI/KO9uJr3eieb/vznk+aFuNPIpd
t3Rw0nwSn0a4ip0rDO4T8hywq4ZQqETQWqjK12SM0jIT/Ei2mM58hPxkqHFWCBOI
D+O3X7XVWrDvui/ny+on0uj/dftFUQpzMSbu76eDhzs8i4Iw76T1j/bReltlorwF
oCLepBmiOtQ9M7j8nTo/PPqu6YSfq08tBRBTo4RiaTYETbsvYGahlv7vBuulXZMX
pMAL3KX1AiuO5X9SQTgtGuzLd4hgVGIUcHoRBmPrh+lB1Lo1nXt7iv/G8wxYbHJ2
iWdlhRySheEUIgWyZswitEXlHA4JCqjX5lRsc9YfR2wbpHn2MiT6OiIhFdThK9kd
6757SgHXc4UJMW9D1WuWvnk+NrRWMQiIztcfP2OUlFz0vAxxdoU3Kv0aXH3+9g0E
pn9/p+g0c9jzIXIybESv/PmzeOKhTCnUCKkRxvJDqTJ1JdQoL7q4OUv0VDVhD9em
habVpYv9q3gnrlV4qYlbJ4AMVpv6KMLmsN3YHUfhCtBvU9Nyw/xiIL1Q2wIdYr8Z
2Dhs7sNwqQs/j0UOQsjpBK/++2xfR2xBhIF8gFN8T+31zRc/Mu5zz9vTjYktRqtN
EWZPDsej0g3208OiY3DIDR8Meh+TP4LCJ96uj4nCVnOouyLv6pB09sKWAsvJnP9e
jLe95BhHCXGroFHI2qOaKfs3yWyWzsw62ouXlsL3N30Qp7aDGgKHcnBudoHEbGNc
FPL/QDVMiqLGe1wOuj0gKoBe1IQAkR4SVjQGftPoVL3TvjYZp1mi3IDa5ca0mVfy
xKJxuG/x2YJvCL8z757aiT//N6Xp7BdlWICjK8K6Gs1uliOMTih2L5eXg6FTT8LX
Ehd85uW8RMh0wlzj9onA5xX4mpY+p/DnvitqEgSpkJatmw2+LvItqOpZAlRh2QFB
fWkSfkSNswKHLR20GKMIYyund8B3j/TXs/a8QNWZ2k7UDV3MgEs2Zm8giSpdXyvH
bB0/qQMcYyeEuBOYijbm4OUHJbutaMdZ7ec1Eo/kRnWOO/Gx9Z0GtP+BTBJmY5O8
OIORhe7VrAU5w+If7gneNo0rYS4hXVgm1wpJqyzUED32MVcF6z7Hw7TuQ6wESYxV
XLfj9E29G3pFAy1E9ldsXWkZ/TlpqJrR5npr5vzGrDBb2kOB3P8Re4ZmXutBLB1b
P6tIpuJMAv2MQnQqPBcaML9TnS0xjKT7XJT/ecTx+unq7/uguHK6uxMrxL2xFSZm
6U6NEjm1ptEjSATI3K33S5DYSuXoQgLvTVTIATgdtg3mVhgYLDLJ7iJcL6hTiEeU
W4F1BNj5SGjAbDlKFp4tcEeOvW9GNHRr/utGx4afGUDVgvqoY51yTEZeshiSMYNm
5vkA33YBlCE74CYKt/1NYbHaSS1RfLiP71tzJ8qXmkLOjG8caCC5HC+ObLzyb4Pj
20LK0MkGXFfT1Xpougzq+aa1y233wjEUq79PUHQhsTIgrZyetEQqiprOseeJ6hMQ
ig9YhZBJLJ3x6kzSw/6/S5XQx1LY3SH7n0e/yCcODi7bl/rIP8Pdi4Qny233OwSL
xMxTYorG9KicKtZiIuMyki3gI14DXH4Wmbttfdfr0fpAwjG5SjrRT0mne4r4dznz
pt8LfqQ9X3OjheHjaJQm3M7t1noTJTvtoQ5X/Zh7dIkYEZPQr07PAzfKoO+s/R5k
1EsWjJ2Db7dugHp9gpsoqDMIKndyh/6EvNJDtq256cfNv+zMkI5g3+ws2A5T0OG4
cc/nx4eKx2LRTeRMDXS2lFvPuj9tBstsONut/vj2Xg+ePuvrm2FXZ5BzNVr6/fYV
x8nUJOdP0BZNpyp0fF3mwfjeg8hv/DWCG0p+QM8PwWvWsPVOa4iCoZwibIaMLJmb
x1LzQfW71J6h/d0CxwWVL/y0QxQR/z76L+jx6iNgv6HWUEQWbHCmiZ+KksXcbAxf
aaUmoDCQOHMaD5P5lyI2I5Vi1pznw5TVzA21AMUhWltJSXjq9Pd+ZZ9I3EbPjQZU
LP9TJqp1QS4XScqcMU1jGVDjt0q1+HMzs2PAMKTGcgJaG6uYCqjIrle15azO5Uyt
dLb1AqBCUwmtHs60BXi6kjp5nKWI5x6vBEfjbI4dwW569x63+0WSeLDn+hs0GFI5
VG3jhFOKzmzpCLYsrZtGjjGDqQDcHmHGEUCeVcUeQPXnL63fiI3xUcc/GN+0fmu8
GQHv6FYviPhQKwKPlu9ppSA0YUsFu1Odcoqnz0cGI8HCcTOYBlsH+LTfSTGjR43S
Mfe5qOG30CctAijy8R7gJ1gNggkYboBg5BFZ2C2K30eRkVDrH8gz7shcTWKN+8CH
/kSiOO7znEfm40u+fUtRVWG//WzuKsX20Lb1YOkhT4nmSYuQcFBbilnLxLzR753M
wOq1aCICIri4/y+MIKwTOMfUjOtH1STqRCu27lybQObAdOX9t/yCcdTDSJqjD67c
Ubq0imzzN/X/4BVY35IarJZXGru0WUNs3UxZo4AQQZ8iC30FQ2NHcvkHNrWbwhSv
6KQay/01k1RxJ4NSv/UBTosYB6tQEX34wb+ZW7YCXiXqdQa+2lg/MZCaJyyD7YUv
gEmfBGRBJPswmVgixMtYWUq4yhlQG2nl8pGdhkWhra5Yoae4IuwJM8Z/Ch3jpbXW
Z91DMyjHYfo5xbqRWQom1eU/8wU6Ct9+PtSbVjs+sW7TF6ZW8xGzjFqENo3RNvgt
R/zPb9B4nRAH0xXb27l+5p8QM177OfkOybn2K/dkYqmLwiyVlQoSsFWpTEtbsHwT
5Z48wFm18hPBeAZNXzc5q2ig7PNQuEF3GMPauk8SrgTmCwmX81PJHf/IwiLO4q5f
ZrBN3nYuoOvQcFqQ9p4zulEtd0sSRFgCTT4FCbcryINbNpBo5r/cXW8Bhd9LoOLl
1r2H85Ks1kY9Qfw81C9S5l7YA93TFK9Mey057SjihsIFndTEG0apJcqISzJQWm4+
m5othuJ1I97sIajxFuw1g7wiQkI279Nqi++/zSpkR+fsM8/BbhyFcWgr9po5qmYs
IAbm6vEiwZlOBslxt5pIqriXbZwmwTqIe3LVv+x39WIhD6qLVDXz+3gbUkN0+kUd
SMUhxfloZOT5hoUiGnn73scUlQ0w78PsUQMKP3z7VwPxXbKtImTgf53Ciz9YkU2R
lDxxlv1HgPVSrygGIxtEG34UP2OpYsfVYSk3vu8blmhirNs7z0aJuVSUo+g93ouZ
3LZ/Mnj3sjUSZQyI99TFr8K5jK1TcOp4ZTH8MK6M/hX51UdKxBiAyyQWqx48dhKP
zmperT6y/Vaj0YffSEIkhXL5MhXKZUhbjsuWdrPq7m8P0rGErT+F26Ya0TVQ4cB4
wngwPhaOP6PLp8htzXZQVE+p86iLzd7yde89IHdBuh1SefNo4iOlXkwoyGwhhJRg
Wo9+N8DqFBwhRrYnoLmS7PJB4/2bNa02W/wkcXetY8MEEuFHtln9yNklJASL8oOT
BID4hISANcqhxnegp7eoVFNijm1hBVtBLkAdo0IqMLKCWlF3cXpWZfhjtB7gxif6
7vFStKXjw6+wVjyuUsePOkruyY12IUNXhhSxxQpG6LXOktiRehRbQXLWDHsUBhpc
gEdVYfzyFEfNEbVUvI3xFvSWByExO//QfZo+6kqxedcGPZnaYwBhFgeFq6yijoM+
8LJifTADJm1jTfSc8jUfko5Y8h9rJjw3ECK0VKcYWkLwR1F3PfRN6146yV1Gc6Sd
lTmIJZ9Mf9tu4BMCePtGtBu0ycOFrzsXHFZVdfG5OTguYjKKjkc7CsrsqNGoH7CD
nP1FvEU3/uTORzdH/IwwkPJZk0WNTrv8WcVI/wRebq0KmZA3PG1WGVwvRI4KfyBj
Kdnc4m4BG3eao9WjG4n+sb1WLINjs5tuCHiJMoy2BOl4NT6ihtnfkqgdTEV1Tloi
JTLWHKXIz2kv6LOOAl6EfJnx/fNYRsJA/Bj4hk2/5uiOfH8/KyXWgRxC25v2vk4a
ZSRKm20Jve4RuZtCeA7IH9vC4olKvzRiabyAsIG6yn/d8EriuLf/n0FNMv1wNo9+
OVAhaZjDrWCHbORpCGeBmpWYAFWjpDtpTHgOdauDIxy/nNp8juRJCqYXK97ZK+Zn
vjpBw7ji1Zc1aoEoLJdMb5gQcLfLW3EYQ4VoU0w43bnzp1nFCNj7x1lpRz4AD57A
DgZQBUFYmzV5Jt51Su1AUxZmfRGgBrVwTTCIF1jFQvchCgUjw1bD19x6H0Ku7veC
JYOrYjtWaW4TtgB76c5tH2M4vrPcKlV0uwHaMGrRZuIvycHVdHgGLKvWBudr2aLS
vBPwXGrnSWwkWmVGgZFp8UZ/x5vatqGuF6G/n0pV4RiGDXLHs21jDHhVfuNHSfQl
shki01cTvtj7B5cahm6tv+wGiqMoVjgW320h34C4/rXn1sofl638mxPlUiptYBmn
sEligVQ63q/cybRBwJk8jwuXe3uP9DwF0MBwdm+9Ic02+d9CyW761rRA1HVMZYej
kmzn1DPBxb74CGs87cxVNgGrFbNKfzHnG/z8ruItSQhT2iFuL2BqXOCAzt6wYdT7
LUdYB3jyz2dl1EQxO5SsVymhdnFMkBP+pMELslxEI5bWx4VEevrqJksCrxJXO0iO
0DEkFXjzdqv07LfmubtQXTmrORMEbiE3+IWtvRtzaFORMgxfcxkvfL24+FPpPkon
GudHxdMX+Lu9R/CFjxlMmpDLzJb7eU+lMKpmTe6Ec9gEz5MZuZf0XvRHmKNkzbzq
pTDPqxQnRf0BddOFjc99wrZzq7tfF7z53ACX0zBskJIuNDJ6x3Zkkdat0WvdyZfJ
lUE4fCcT3VTbHzv+zUhDhZ5GPi7Q03qW7n6LUynRKmbMkHZRg+fQ1/+XuDXsmdx3
cyhh/JAYKKm39/GaX/WIialUkVMcKKy4jfTRmfLxuexqqGH9lRaKhbZNUjf60djf
o2l1UX4CGkylWYeYKpez6r4Rud41prqNFIAUBKUt+6YwYQ+yDZ+2eneJeNRunkcz
BHsiMjDqUWsOJi8niS3jGi8gJCzXPymmEmYZ71cqLau8nQY32CE6R6/krCUiZ+e/
0szdv+vup89JI8MMLfZe9uW17lkjQerLB7LGsyFGbg0+2229De7G7zbzImtKQe63
0PinB6L81siPBeiWVdr0BrIJD/0Ql3qooKqxLQ414wD2UFS56MjLSxasnhUbETJu
pLC+ZyoZnzwsnSfR43bMToPo0UGUwfdJXPkdj8yBCl63UAmSBKfWtLGODTHnBSBi
D7gyHOL/OAUpSuohlZgH7XaOmer/qmx+gqhjc1czdIffNNISldTEo5mvxlBT8TXK
WSp+K85tf0iSDjs+EPrwtzrQrTS39Cz9qM7ZmZpVN8QBkVE693T0Fwdjau+Bp1bO
h9DAKDPEPIZtjFEi0SPjab3f9PuFfwTe51P47tdN+I9v0MD4ben9l2rt10k9WAbw
1w5bc1XQYG5YqfeGty8MSR/BYH/Xi62/smo4gx5MULC5M62sWrsSWK5m3Y4FB5pc
Ed3SbcpltzjeHAK5xTArWyBzm3BuZLb8lNWGts3sV53WQsU5ciowxLHrTGowOp9y
BwLx8w/dQmznXSdRDRNloYO0eFI0EuapM4scBIku3Ul1uL2oXQ+z1bET+CsmYMNU
mYGv/QMjsHWCgS7XOCbQPt0CJ+ZUpLnORnz04o6bysGD13zrNo32bvOKxsulyRuW
CNSLyRunvTlfZlrgrrZBY7ddFDa1OJOw3pQ6g9WNAGdsUQ8GjsAdf/heLRLXyOJs
EbfPRGAGhtEb0iiYhAr1AX0K5AK9k62OFc0gMn81+jAd8coq/OKQui8n77wYBMNW
8WtZnXgIgcJR+aI197HPAI0v+AxGXM01Kj8rbFCtXyFuCUtIpS8YIlbx4Eyy+sam
P7LLahpP6Mhd5kO9eJhKtofRY3j2aqIHzlsN9D+GY0VO8wFY8Y3MMY5esTlpS4zV
oMxtvUlxly9bmot4p2Z6xGfCWy9JIBEUwin5RDQyraG6+3xO7ZbfywviM9M2YmV3
VG1kKvdQk1dOyGmOXjpaeKphF3kH9MgB8qknJSEiBRpGvWRLfBuTwiNFClkR3BIq
lygmXZqB2x0aYYAdyIilKEC4QFddPbD/mbS1Ychl3f/y162ar/Sz7C5gKlO5TafY
p4Lqem+G9uWazfD/qR4blGQbqUoZfQLbWlcOdo0DGcq6QrxQsyxb8X4DqIgrzJw5
UGVidYyiE8rAnvW7eYbxVAmnUdYIYJP9U4pYwoWtNLoVr0phgYB7zWBKf643Zojx
uYaQf9Kldoixco13nLtQXxIHnqC5gCheAfgvu1ophkI46V5xbGfCb8VN1MGQPF08
J8Y98ZzcPy/pMui+jqjDJ5P8DwuRhNopfYbOWbMSzUc68YheTP4aq8Y29bNCVO6D
ZkrXiNuZqhIgilHytrAOKxvxrAN4VOR1hAvcHkhfUYfWC/DJ1zIukbG0pEAuOUDx
8cCB9Y5OMs7dZQoMty+19RTkW8p8jBVNxR4SifK5vJdSe/MC01mFd1Djbn6xi7ZN
PFcVTiuhZRl2v+Gl/VtuyoZtAhEo5QgjS5bS2lFKofuWmjMdNq7jXwCVC0MOXCiG
D8R99eQm0RLvAIKNv/O1R+n8DuuFo9YpDU0Ks0fHwxqpRonW8Ave829afXEaF3HT
y7ACPRvfE/dvHWxK/4KGej4tPgxqXG74KndaaIdAgZM1pwJxLrKZ4UbouPPlH/Wr
M7ryBw1BDVyACJ7E+CD6d05NU4CX3FT/VAbkxFXM4ztAMa8GN0ndeGeOpUQn/Ric
9ANym3s0roZe/GME3ukERpPpVySLgXGEx54EPCqNnJso03MKapi8Dm/IFBZNRCMw
yvPVrqPNrmtrtC6WZlaDyXnS/VM790JO8DCqXvqnxj59pniiiueAgk+gqJR/fAXu
z0LL9/2HT7UApVUAUTqmreLpzGfSW4yqH919lK2cMHpKY1Qu1sxFMg0ZLeLK6rYJ
ylrgrhCPjohBn4Zt0sWT1U1+ltn/Yvlg0RTvP1AGdfDVHeanoHJGhiRGzuKM32aJ
okDaI1k4GkbaXQd66ZaBEEIBcOlXTexp9kM933fhia4fwaHktBFr4eM+jzNDuXJC
Ly1RRIdglc8LWTyK7HBkC9Qe+/vBiQbh5z87FxwUsSqhdoSCCj6SILC8FSrYm7YC
8+2axXdeolQ3sdOeLqpnV8SE2PraStlecOHZzdTKtFhdNEKLdISz7+FERa+dQDT+
qid1sPxyw980btuhrAuvaP2ULQd2c8Zjc8ZW9xqFbLxn2PzR0jSyCnBCT0j8/X7/
r6CGtrW5UrwjBKD+SeJaCUjTNPwZTINlTHmvh7iPWRaiwLv9ysfdHJJi9eTAbDMx
Ck9ASXcCjcIjGBlS0wm4P+/kRXmSIZV53MO/lCkzzd50IztM/RM8gmSJV++q9D8o
ViN9q+ADViozwb+ithECouatsqon3D7NZ0CMfSykxNyIklkZv2jIKKvzuOZ7WTs2
W5gBR/35NdLBfebjHQpGdZoLdnBs+jyrQzQVtYivLf0eLYvvUyWUOjynon1iNWjL
qSrUntWyCUo8oayBWyxDs2HTk52qwwfdoLpRF0CEWRcIgdUaYhzCkX8zqVejm//X
r6Tf6JRAtKLrV4I2rhhSjs3FEVTNJQgxxiP55LX8gRnuZNHw87/dIUO5RxXsepeL
Ute7gG0/sXhfqiiOmsp/r72G5F5OYpHjc8lEayWnvNquJnVfcCZW2l1/hOM/ZvIC
BfydfKLs0Q2GjZA/5PqqrdBdv7H0QUghnP9Mapm80iZF0jVpb2DsrjUpEIOgk6hf
Oj9x8xIaXc7M1Q7P9puEw9dv2H976xkyxYCdIX0aUjaQa1yrnH7bhzA3nGAK0tKK
Jng/fIaUkC2NZKMJu3cNa7Zkx4NoO3HVRNqdWOT7e4DfzG5riWPPAnMrLeoSEMR8
yoaGVsGtJrvySXObF1AdBELgizx6axCwnxyj7dTOGLIpdSqvtKu54Gauc+yQYKPJ
b/QP6SW3ih6bjb2815FRcLKUC3dpUqGZ8J+xgCyWriMtvrpKgsTm1XDYo/hE00b4
e+WMDhTiQSE15CnUiFp5+827UgKSeNZe+Eooq//7gSDW3ZnZTsGz0y+rmL9rKXIB
5EplnNsWJFYf7w+N++hi11oYoXEszPuiTisFDrnuaXIN540mDehvdqOqNCX2rBuy
EI+PNU4Ksv57BnNGIKXMQE8waNam4pvmcoapp0N5d6dEyM6ThS9ukT6GPv4Kmeay
JS45Jxn80BdqKgr+ksOcVsM5hamFW3JKBaVZqbOEBGjvGqp9i3cUfF8nDmiM/REj
TrJrF0MHIhO8eAPcjTXq7opcdSPXK68/qh7Mwy8+fIz7DhRdMrMkkVfQPwjYigTE
kKRJ3BCARwxRYgdH7Mo9SiEpsHtVkOUzB4eJMzaWlakuomyoS3/ZwIADpu3bd3cM
pX+BwQIkkDHgHDJk6mm+yLeQ1ph22pKZ63PA/b2aHbBaJf9TmULZmvBf6GyeKvt3
E3tvixUk0s4aphfWc76HFOlDDQrfS/7KmQsrxU2CrwLQnffcfazmuKQCK6JWgGdH
EqhXgmOZv7nOtoEEvE7npMfGwjmoYylcAP0mjSTpGj0zWj011kwUgWPHPAc9gqNz
rw/WNlfYH7+//Q/Xk43B3suDGmqRzUwFLkL8a8rsoKGZkhmD0gFt38XfX5zKv6BG
FOuKvV044R3mtN4l7Ebigip2rgQRydUzK3j6ZXKLRh5W7kwnM5NB97uc9dmvKUKA
2BGqN1wvgzAvDW8T8oCBJiLmTdNpzmXm1YWhKx5aKQq4A6x3H4nvSlC5n3p6kyrq
nFpoKK0KVmjfoq5ymbgNvg6uycweXWDimC0GTlOqLx2zGIuOK1dDCUemaWQAGnyl
2B1qNpimQHPpA6vumnAC4AacT/McusptouGVzL6+CIK4DtG1ihY4JamzL4uNnRzr
y6vHD6pQ2QiQCK4FKhXWhf8rlEk5XtxF5B2kVbmgwytetdX3sc2urfl+7sAksZgT
yHns3srD+Zwm//RzpXv+r1m2cFpPFwOjVRu6YMjYa60wlvg82FZqkyYlZoHdHvDe
FAZL3wX4TAGyETpE1geaPKhPmbii4/zWwg/rJGtceOw0RXvNdQsHaOk1E9A8SznO
3KF95V1mcudOu5zna2BhrdNE7tF+Sfww9SOwEuBy1AgBYEYnhWY2HoQdq5mDsCOp
en48es3LdjgJ//2qSwbUP56MeHgPuOkffvpgKix7Z1dFRTYT7BasRGueueP4gHw5
3ZUfL8VF8jgQRp33R2uH2cJkrMsX4nxzk/YeDFyoJ1zz61In5DGQGVdPtz7RV1Ut
vYln99onGA8idd2CmSnsqdmw39VgSZDvW462AoLjFZU6QgPQO4/UhvuhV4vBU2c2
dwB0LkE+2Ry+WmGfm83TPCDpCHIZwKskHmemKLTcuIrNHkCP8rQTarYuRFtzjC4E
BjFllUvlOCt34pAaaga8jgCxmYBaz+zo8SG6Chr0GrVqnoYESp0L9T8Dvzhk/dmd
v7iLBS+iFNxQ0uwIP3wvQXSZgkyciq0yWfCxxg4zeYVYlUzoesEH7w58SLpwSUID
I4SW0N5xvTKdjp2zou/+1lE9t5ZwOAqNbJ0cQJrDzHxtn0xr3d4pQrg1uIG0kByy
aRGrBpa0NhdU2l6Re0XgCLJW4KO7/lN47A8gYoBsbZSc/lgDBAkFOE1UKjRA39Up
ojMspkQJrbidaf34ZuxX8ke128x0S8/vQB7qCahi0WSv89DCRydrvG3xcooThpPp
LmW3QeiMStsA0UlZ8f55VoRXymITDsoRTZjNzrfLL2TaEVyg5PO7XV5XMEnhauBX
h0VaaS4GWTfGNJ1V8zy7Bd80QKiyrkY0liJl4obzT1BOt+X9anBchWe6TfQDFBu+
dgAodaP/hi8JLJNi/w317oQH1gzhcTQNc93Gvgt7zdZX/8+focTiCyqTHLQSNvor
qeYfaoGcJ7Q4EV9QnRFOuOTP51PzZR7rddGcLfRZSmku4KzHatH+/eHY7I877Lmq
uraTfBdbyRuUUEtUMiZpUGBViJCHll99sV17BN8rBCh2eeVR5OQ7eG1yrkytXexb
fJU5lN4evC7xbPh75FukeQTk4XG5yoNzVG90xZYZpJ7E4Oznwb2h1JUQClLDnxF6
bdCbGbWbxAWpwOxk03CN/Zz/80Xjei85lwaUgLXKT9G6gHlG1Okku+FIPPyj2yf4
KV9xqVzEJiI+QkQZAlp9i/CBF5XJAKrL0algKeM4lYLoGrtIGvpOTeypjxNx8BZu
sxX1pWaAqNACo8AJq3auRTu5Qzl3/JWZNokrTT6lylzBE0uMiYP53o9eZtBrO82Q
EQWbmAgxSCmRnfN2WItNhm4htXKEqUA6Wvp8kt3MDASK7qiHEGfj1ZiuDbBsSfLO
fU3GDfpwdPjhuvAiWoMZOmHWpfzswpPt/+lPcBczG2DY25fqNwZ1xIaFOGdKHwE0
9p6T4p7S5F5tXinROYqKOBaB0UXDSQhGqIAsSMXOfP6gx5vGXUQdcy3gYhTEzZzI
oWduSsBovj6jghLNF9AC8UbbYdbkJQqC8jAlmb8FIfgoguRrqQ5GPZ3Mk7PZwigb
LlU4tB37d3Cu0TvThLaNXJe1udO3eZaJi0/JXuRTg8TB3Pj191ubgqoxC29WIHv2
hnodyWVmBMoRFE2quXJr0luiOnPlnow+heNci7IVKEJ/7U3Z5nS2Y/TcMV7xzy9U
BabcE7VdM/+pA6sI2apU8mFRapAyHXOJs5WBO175S68bSAy0LNhsasEeI3cFETMa
ZuXUyLiTkpwpaCVMK8stx7WPBS8W9bPIR0uaBTBO15lCZPHly6eT+rKJTe+Q/+p6
2JxCJyuF7vQhH5E4Hd1x3m/MnXbTA9rzsKOq6Si3mVtOHrEanIRLHFCS+jNY1XJg
vOQ1Bb32aGHlmlWKxLZseZt2sU03tBJDe+N/496gparx8XfkYltfE12c8BSU0QqO
h+nXAutJlPnoG5bUQ0bYF8jJ6gsh0zk3vGdMwOzKFwVlTGuxFzm4hTCNQo5LAbm8
rqR2VZZkA34IRDXdZehi/lq99Lo2xuFdWCaYJSF2bcpEhqH0Ln3XWCFFoHU1RrAB
JF+nhb0c9vCbxwxKVW/aHKFY/IMILUfu6ILXWzXiAt4so0wIl1Ji+RiYRHeISd7v
VT5WrRTDkGEber76Qa/YmC/3V/bREM6d8HwwdnE4rT7988YgWcA3SAnzw0+7QgBO
dmC61cuA/ck891PQWz6q7nVltr3cLPMp3Iv8V0z+87e1+Y4nvGr+Y6l1yd9qYDrZ
m1581M0vP5jb4XRqEwdSqSEKsIhMj+UunJeMYmJHS+jCfldhu795lQhEov5xKU5f
qldJn8K9fhcf/45KjawgUU3sXcFtJV25GF1G6EvlV2S9KYR/vmqqlV7F0EvTusqS
jxy64eSTtX0s3Fb26ACxxbJA8oS0lHaVFTz6rrg0i/uL2FAkiXgHb+ay+eqqOkQO
QSgtL4WHp5uDzk3FGEG3LaUR70/ZY2y+4JQw0bW7kMQgFGvxbJzayTUeXHMbT96I
tkLw+IIjj/4nFsZtVrDmcTDNPV6TPVk8vAkMwNiBY6Nm3pHW8+ZSswfQhV2qtGOd
PCcxPWV+uBaCbxEKmIjs5Vv4Ih5Nm1DlvuLOT/D0WbJTxkmzaB0Br84eAr9Q0OBV
9e5shWBRScw5XXtRoDWsTiYMIsMiy44vDBPEPp0JUe6vCwmn1yWAbuN6hbnu4R1Y
w8o75OBo9GAFi17EvaSP38Bu+HCG+mbxXHDPkJOEXBi4Qpl+ADjm5yeH/hAANhgc
vLgCvAK05virGzipBpRRaLnSiQW3XBNl7j80RmIZeQBc6bXV/sAVPJK7MA6KeIP3
CLJwoSgKHvbSeiYYgWkGPPZ9F1iGikbiAB417bcWBXUl3S8RqmImSFFuGsaguU7H
hy0B7ayue4zTKsaAJXGOHKeaU/F0uhFKcxpx5vll5cUQnYUcJ9JlAlmVM0XeiJ40
kkZzftBk89xm83zye0UoOMNpVMlvXnOjjWeYk34IuKg9auzQUmdPOSH/TVyckcdi
bBFKvcBU2k7gFHfxhRRXSe9oCrjhWkKhVThifCxMHbc4imvqqBinkf+60uMsZSmA
LfJV+86ORJjPrxwq4HVXjIfBmTMcD8OCTO9DEUy9/QnvIbvStLzmK4KhgbVfAHnl
bjwU+7C0a+4YUz9NV9gHTCnjElhmmUAJBOiL+McEGDvp051y8ZdyQdiC40Wp8LDj
shvZhIlEgbvN2I06/Jk4flGtX7lICqJmlQSiqn2B4BbLsx9fVVeOG6r21fE4rC4+
vA38hCaiuh5CJ10dkn/Y2vMppuJyCIr9yeAuUrjUnL/LoUjPHRL2WyPtMJyJg8Ey
4VSXtkw6patOZSWnfscUZAapQ0pKtAOzR4QzR3wia99xgV0yZdnrVtJMJRddVchW
UDAS4ZVH2xxF3nbkBQm+4Ow3N9SMzPopSRhJ0xk9cmG93bIW7pDrAhAoWPOYnehu
cCkI8UdujgPC3qm79dCf14JBXA0Gro4nYRI9khgsPe0zwlsXmS1N8SI83xzmpWCN
BT1g3TKMdZhdocR7yF6Sjlyf3r3a+3ng3eDyEdt4ICLrvTWHBS4nRSAdMzDDbH0i
9TDOXDa+Q0AwO3vVKM1tD4i/z+6GkkcuR2ptXhcQQs2EcVXu0vp1qZO/8/D1CIAp
Gj6KxJlKcbdNnOi5P5sIN7cwcLH/H0uM/24dlNVr4Li0gUv8oYCWH2pI4cbdJzMr
NTGpi20MDgcC5Or9FNBc5HOotTW7b3uJgGtRcpFudCv5yyjYavn0EzsEw3ttpgGw
SInjRs3Mh7vTXNjsm1U0kbrceMYBoIfuhEdaUGpwSb327C0iKEta1FazRKjCVqvq
9RJVBqGEq1Eatrb80emX5TGU2E7OhqZvkm15PJRCR00DqovNEL2KdgTzN/tBVn6I
t131SKXPvwHotFnghIqnEdhODL0buhxnovrbEzUWGxi+X3Gr2GrJovYkuSRqOw4H
hBGAGg7IVSAlA3JEMm0dxxsz+MYYcR5uoQfVOMKEUP8DU29MQZJ7SKW7fHbD1joJ
bfyySn/t2iOAgkOOuFspc6MlkNcmkJAY2bLPgiB5mwipb3r01lGeJzxfbwfexdHI
rCnN352sX6gdB2YE4Fe8GItL8av4lH0kSDh339XezhnHH6O7rYgTb8oXgu46kuFu
FtKL/m5uhOAUWtlr90tdSA4FbdhCZzgSRjxMxpvF21rEErxwfNAe3eZ2fVF4Wn/L
0SSwmEqEWBzR/mwfBsCi/OxD6AWF0i+gKY9IlySQ3RxIQo2Nn2P4z23xK58SzU1X
fKnwVk32YWvK6FBoW102BRl1dzv/30dNv7Nm7ywbIInHCCJFJ0Be8rxpWiBzSz+7
9EHRV6oxtbMe6kKQP8MxhaIh1wOAOLmzMVZUhXpBnz6eNCN6iJVHkom6COpfIkSd
/FZyTAmNeRrh7cBxjhC1F6Cc46r9iCUs2lgYOG4OgXy3/tpKwZ4RJqpfMtG3yCUm
LM264vXKn86kY+T0CpyoSwH44sROb1oERG4fQE4/pe3nz+79uuQZvDXg8Cd0my/S
GkY1pCa4CtHq7sOqzUe/GZQ4iZQMkprvQJXnagDZqrWs2ZCYBhT2Tdbl08w42YK0
8sbjAdPpu3ssmeIZImyTuakqKcRxWMNCS6qkJQUb9am2cIa064a1TEKO6GJNyHYg
RB4oo6Dt0uuAVRcROm8ZxYIEn9sh8TT9shpJHNk8a8HycC4iSnowEUpLQIx0VwgY
XBh2McwdKM9G+sMisAYBZ/tgX+YkrvIL9m0ZVTJu/8Zw2d1elYzvCyMlpKAUUpGc
ssKcpiBOFNMpRYmpxj7zZl0bV3iTKIeYK8Uqj9hCWh9V+1xBbCYzYCjBwvI9LvCe
yFZtt3kNZXZb/LiIndqdFWiICKKHghG7lTNcrvHzhEdmIH3eL1Z6cu5IdOSrZELP
a7/WjBpUDolDK07uzviAsnlIN3oH070D00IXri6JdA1U6dYupJlmbe+eiC0/I9M8
Nt7FjJg2+cXDI3bngEwZDRjU5MJXQiwPvW8fMb4VQP7FR1eSIFLB5bBay3gWw0Gi
AFQnWpZ8syvJKN19cdQNIj7sebbzR/FbJiKptHdfS6N1MmurEpPUMRyajlLS3zBP
DQfP/Blg3M5k9tVz5CXarUX6aybdhMykJtfhhvm06DxaSa3lx7biVPKIeU+O5WRE
x+Hn+34L8zpewqYWa8VHwpTw36TMfEVOcaPXryRl0Xy2NkM65Ms5YN/c2ayGdUHv
jriKDgU1Az6WMEzNz6snMY8ml26Ij0ybRgOlzSQ2QvOyYuJ2kYChkv3kiqwIn8ZS
pO0J04PYGueIiUJF7bkiTTDMdiODZ17t+NVBJyV8vP9Y4E/JdIvB6UZDGFXY/07M
i6ng5VR4LnImXvGQ5Yoo6cb24H9wFjthJo8c72ZGc/jHS8ayir/8oRg+sjGFJFCJ
2Iz242no4q0nsZqbT43EyEoY4bPZahAOOaGmcz3eqYmjZ18YetDmE12qABYWgjXJ
x+4DaI/AjGJI2X8mznujEnSGRWU6hkQtyB2MW+lipVDbhUi/sHXEyXLqqOSX5xTF
P/B0xoLSjM+hNRONpH7Db8jKlQWAeA0IS15GJZCTTiZo4jTjey6wQ0P1j7JRcgaQ
VyOMwdCHHrKVm9C6kkLmqZTGxgQ6bVIgU58oLshdBc5KW4rwg4bot4dM1QANfd2H
Fd1nt82I2H+oC5oI82b1DLCyh4UDXWx7noN9BrB3t//kSN2vsuU8/zGfNMCtDaBJ
5UfP6lxrM6KxxZsGrZFfANBTOCTNCj5gZvjvNw/xWK35bRAEWnTdHjrhltixKmug
3X69kt5E1Dmxhe+bwAom2AkAb4bx359+YpX8cekY/i+mvaA3JTACBD5Vqh3K8UIH
kChsv5wI0fahlQafSX/Zi++Kgi4rTRBzXL3gIFl0uWtA8UMgpYRAtfeMUvQnUG1B
fCHBJEarOxzhtMEXqcZQCKo4QD1lH+FdMu0jvX9sPekPkbLEj6+yb/hM4QmflWGY
UGUqAu5cqM1oUmbhVEgLTboF/H3kvGgSggEyuDHsP1hNJ/BL2ourMVfbt5MtK84A
22yPCb10YWiu2YUOi1yANHXiRthnQVDU0n46pEY2gJFJ7hmEO5Tp3ZJr9o1RVrfl
UOMy4B0k9Tu3ss7O7+MnTRojdGo9j9YSEb7Sq80efFNg3H1oY5UrXFzJ/8QsNTJL
6BrBL3Vpj58QR+D3Loamnd1igzLiPJRwtvUwh9Vb5z695bJJZj4/oLa7ktsLXOJb
b+OGWGa97O7NdwUUPtOsop8SiosLxMudwA7eBQQty+1/kMnDurIQbpj6T6lY0lxe
IY8Srg/IoGG56PCkDs7vJRlHZyJhAw2B2bwRDTkcFshF5IM9YOl1LKF4NbLWmXsP
sg8jzyBqXKzxvRIthn3I11lBErjV9a2/zdqfUHgPqboHT0N+oHy4koGxrtn7/rVH
1c4ASEcyT0XEG7xDoeu1Xr2dRDaVTCaOftDlKTPpx0Gq2gDURS4J9xRKcnJdOBFD
izhBb92IaqfCSjfmmY/2QjxS20uxv8ya5x1hTCcyJZ/tW5dYoEyVdFg5vg9Xi8ZQ
+yXmeq9tH54x/MfpxRBLpPFcmdRUWpGcE0oEOt/veY4LvJd30QblQcGohW/hqHdK
CG9Wth06SGnzO91ExLEBpSwWT6HNDUHohxao6rAq9oFSCqyoJcVTBZ4WlEEu6fdo
/X73CElhXm2Bunp/4WePbWRQ2kY3Oj2jni00+2l3RLeNYFQ6h8tbC1e/BNdSn0sG
o4huQUvjnWIcLW0YVPo4IIU/bwho8QW/bf5jBe6gErxsqd+QGuRWjIPfXn6ovDeu
7eZVNW7zUXns0H0WYMa66bU4x/je+442y4+IqIoHOZXMCxh3mMycoAOMdGfkmzO4
KvsDaxtELka5Gl8hIaQfm9YWeITyL9OAslfwWKQrAjEAZ7R3QlmqDaV2L/zvhXVg
aVOqOWvSFOAzSPO1yFETiR9CUR9zV3fFiP01obHVyfgqEHXmYgPKL0RmyGzFQlWu
AIgGDPSoFi9J1qJdtkCG0xeudz4jO3sJ3S4zvdTaaUcHvpjk6wf5+6pQVbqk+MSy
uwX3PR8IWvfy/6q4l8R56rzhTNP1KSMyjw18N/N8AAEg1n7hHeRxgJcCmCdcPHuE
TA6n+Tw38HXG0+AFmf9R5+/mQlMyqlwXfm/ja3mU0SEZPGTCXAuqOV7pKHbnqWuQ
szK3PrcbubWUD2kLIa/Kg0EHxGpgEoZnrmItTNo0VfYcNOlp8Ip1oq32Fe5NmoZR
KtifjWKpq8MNz3k07BosQIZX0QtZ3v/ViWeolmUyKYF1VdBSalmLm2Nwa2fEijew
Uus2o1HUTcxibVemSw/GwbmEXxZIINfSf6F4749EG56WqThQFIRje2O3Lv1K5r6t
VsVACG23DegeeDgnZGn5WfJ4PUZ/BGw/x77hijUQQf/Au2QUFG9vTn6qRuIQnB66
AxtXMPd4Rac4GKvVvDDpwdrk8HUL6TBbzurCKdeqxGwtcEODFlOCzjFTWvexYkoD
PxPe33fc4uIWpkkUzThKTRvn0R8p3ec9bmrzTQ/JzPhQAoegOoIwzIEnYJQFWk2q
Kv8FqKzCqNuyNxFd9DRvQgFUK7D54RgXv+UMCSavc8KVyJXMck3wuU1XN+LYKvd5
YGHtioZjXnIH6bQUU9XhFIJ29LGFiJXMMbfd/oNXF21cLHy49L88VEL3tawOUYD+
BCJrR+l4eJ37XPIXFpfVMfqxm6X+s/AnUkKirrzHY5MgDz5fktIlFcC+JL0zwESS
XQkbA0ddijB6sokaVhFPXTZZiKUMBPfHSE5MXf3sH70SYzjiqgKJ+BAWAGHQdUNK
+q24W2pBaHTB1K8ZbBUSElBjXcUBIOODW9IupBbM/AM2i2WeljkA8kGPa00bHK6f
UCTk9Ngr1Bq2S8I6YsGR2T2dHTF9e2YkqsH8IgR1V6ymnnq++z/juEkMb39b/Z/O
AIYmSW/RLw2HQNTwH3Xaw23Kqy1e/UEEF4c/6qJdfYvsb3gXQC60nwjwYmkmtGb0
MdjLgXC+mQ6okC/exGIYSCfIctd3cfFnYj/bbILpMkzujxPZDQ0FjlZjWMrsRFMN
krKFauAO6E8TY7C9onAVrtZY4fbWEuo9jIx1Iv9ZTRNI6VwerhTPQoc0VXHS2g+3
6fMMxoCXJWXjiUTRNF7b9+gekQXwhnL9PRiSiQbid1LkAtH9naMAaTbBsJ5YUaMd
eU9nKDKoIu1J0ClUEo+Du+xwCPp5nnlsRE1JUHk5zYguMZT65L1IuAYkm/X493vp
yUggq+PrqGbkx6sB63eOmTHp+uytWFA0mLQluFMd+WcADcUVEH6TVTIscIZ+v5PP
pU2+6lJteWrPC5floXaKitHjrtI3mRRlzb8yzjPcPhC7vt7Mu+yHlLrr7DItfDIl
hciXyVLc9hbIkb2MxLWiz/nBBed6XTTKd6QUZhYJN7hQE3oGc0h+Rhg6gpsOiKZT
QlcjlJeG/j6sbU6byy3O6R8+7h2wfBEOkqJVBsHMY5+CAVnEthUaIzcltL6OalmO
njZ7e18Em4RPlPv2caIDJxau4toyH7KMdBd1CGvWTBY1oQOIuWIl7FMbyJfM0E5a
PXKa51TwO8P8Tkl7aQ6bqTsN/QW+xuMx5+C67ktxZceRxn0Eer+1gw3HufcJjPB2
x81fq+AFr9D+HwXbir+hC9/k+5umsI6GEetRpYBlD3of/QAqw/EPDHhLP34u8my5
Qua2ZrSrhqwrHTn6JVDZaR8YerzoZbVO/7Z3Udg+5/T7A/g8Coc/neBG+D4LF8dd
ByXFqQWE0c9TBz3RDJY651XEino6bNj5sNpNsRc8l5yrE8SUqsvCKyR76qXYlIVn
o+jiBcKUuhWIOrInFIw0Kja7rrYY5qb3huontoOQ7/KiNfo2hI/Wooee9E8ipNrJ
hsNgEZGt1U1fWvNR6SnatA3frkI7J2b+1GC/bQQHHek4zf3age57Em+JM/TDLe0N
GgCn/zUDvy9d9tTthBOSmK/3uxH5Mfh5Yx5/Rl19u7wbbwD2P2cTVbaI4JAWts2B
LqS28zt8Z39FP8hke/f82mpT9c77gguXOZO1ud53VCLaoTadLXIwFmOE81nx8m/K
ogg/xLAujxKrXA0gqDmcrFF43IdwKgo9QLAygibQ2EeNS+Ldx1GN166rGzv8qaTk
MzbT0G2itzzfC/YDANaqNxb7MEHD++nbHPpjYwvM74aJt824dEb4vULwdNEzKGK/
DvmGK+3r/qFfe+856Mq4Oc/k0Pco6km9V0SGiVc5iOYLb/4QyIgfvfKlIwalugiW
OeCtcAIe40arcIBp2/eKBGyZnlLAwVSPr+xiTC3A7BdBBWAiovzK07vHooq7YkQL
VU9JFV4YxPlmYGe+hh/8s+xYb4tF6TKchx3FPFVsgaK2iplIu8zD8N/Npp+iOjiR
wabe0V3y5NkKnhhVJRP+6cCAz80gtuBc1fI0SpbdNIllrHK0K79gW88j1IZl7flo
ACoO/7iPR5rHWje5+zDaIFg5plazqDsBVFtV/5wNYfSBP77Bkx9H+EfuOzyIAihe
DI7cNK970/2C3M4gZsHTb5ZyMO3loIfjaBrfeN3Gjxlaw+bJzFwD3ONKtJlFPg4G
7QLBKnplGLetBFJ3UrkEPWTwprbImDt2+a3Q2PogigGvBtVfA1KrO4Zxki/9cJAS
MOOVraw1sAUzZCD63ishiv4U/OfvJIf9FHWGR66ianLTkHUj/bPgRkP2vMgBW4DP
xcgyioYnsNDrIRmZJZG5PyJpDYwYnHMwp/6I4ma/S4fqEr24b0dXtamDIAqKfMh4
8bJhX959uXVUWZGbdXz3WrVpjHYqLWtt9dOvBZQUXRlr4sPULa2rQ5UnAU1Dr8C/
mLQBHCftdBvh39kwh/uHgkYB2OsamoQB8msz2tfRFw/3otUEO3PJs0XLDQCZYLoS
o3q0NJ+cRZ1D7WGgzwGlyTheHVjG9hrg0OzqMKWjshmZs96SpuMmW2Gavmuehx30
SL/Gf/ZNMDsoqNMvFxSgyylgm8ef7aPj8wkTBsVMdipD3nP9ty1cqi8tFjP1I4RE
yOzX+p3GpTfvvJ7WHgEE7EmnRppIEP7GcFTZi/59n3ecdTu2gE8Qq5YJpU0jwjbt
y9G7VAnS8XKpdO5zC53AjfXx4rHLtRFzvdes0PimplDo4gs98GoxvFisjY+UL82B
Bs84D+fXpfHm9w8Tf93kSboiYR2GDhdVFgzsPL+Wo/HjKqZVw7pQFn/hRhOjtSZF
EMmcO/GqaJkyIf/cDd6fK283eW41HheOjIoggXtR7/RgxNgEXs7DT1zv4HoB1ocA
f+QOKErXjQYsAJSXHrUIPDsoi1kSfQc2KiNJj9PtS3Qdw8mFFinv0ZHxTH6QvCo1
eUBLWORjeacFbhnVXaZ6pH13Uns4UUHauNP7o50yhQzGXuAq4lE/HSoiJpPD+cRT
bY6sniJR3ExYz64grhRwSsmcOJDmG+L0NemCyHytYKsBQQ7eNH4e5Ny5TAjsCUoI
FQCV/dQmTXNy7Z56jidWlIyWcOe6dROb5ZCLGkBCCwbI3d7yqFVGZicDB65k/QCd
odp67KZfBTlZvbB2W7uGyLBMx2iP8MZnXYwwpKeYR61UABw1cTcCyOySxdNNPjKS
cYVK3g0IDzJyJYxGkPutog9GCkFdM2AzH9dA5rbW9lhfWsE7x0LRBsKzgpf56G0H
2s+hF5XA9LXGwmlbb2tpTul3uj6iu3NLtp1rvFs3jdNzaG3skj8+uarMS0Ck3K2q
6yBLRUTo5RFiTnkSD4c1+9vPfcEPFz5DM3O5U7d1xPBMvvfOxi7TMUjNhbsu+Hab
5Oi78IIqvMWvNwg8c7AZ+HVgwVz3DHCSgJct9LTOXWi3mMtnyi5/Rcop6aBdjd0s
PLrKm178jO502yBW1WjpoVJamQXf+eYwCAv9QooeeE6PJWD3lSF6zCudu3xIBpo3
nTlIEMKGWVKJ1wOUQTF4iM6RUNMmJAcIGAd4YYrM2XEFzdR59m2utRgv9NBGak7Q
KGpHnFJKFS8RePPu0a8+yVlnpfNF9vZBI/eF9OuMS3p0ii4wWxlDZT0pW4waFc39
KijkX0xqeqpMamOEFZGBNJgwgp/6/U5BYsEvkbKUAabkslPjApNcPp1P2OVpppAg
39napNgR2CWKm2I6QrfYFGq0cDMxjKNfeFZ9gSn5HXofcgPbm8BKNg+RsAKbXsXy
YpGRTu/w/EubIp4x9827t1uZ/Q+wCZrVpFCRBcZJdKO1GGFrXW4M1HAAZBwkJNB5
hI1TcOLVf5zXR1VMilJsP08Fkx9DOA7FhYAjY2hrRcz6g9wrDTO//3WWCcJs5BV9
qpkzZZ9BcgfsL3XctLKXSk1vNAwMOMDRcZe9X9zaMgxLXIK+/HToOZr+aqvjoZDp
+dIe1i6WhvuDUmTkfLYNtE1oHLnN7+dNgN4RIPa4DCSvOx8Sx6Su0BiTX2ZdfO+V
hiN4WecD02to476+kRJMiKPFH8uktv/mN+aJZaLwA5HlBKkZyGb8C9wv2qriKM2o
BmWlRKTh6EE72Sk7pYRKv9/wkeUZmX2lxX9PBJ54suQ2jrGvv3ZPXzUEZjhe0Dwo
aFR43CGqaMJw8Oy5kreQWFNLkFDtVHXm6nzLhvW8qJ6+fkN76Da+12RhYFXrwLmN
GyTuiEZfKIfD07Gr6oidkBVWa9rctIg1Aep6na1EqAI80+EROvfhb0bg9y05QpUb
zlddUVop11OJr0w2TQFX1NWFAw6bsvw8WLlNe5LAVjy2B95R3MpRJfDxuDTvZJdH
fSStbp4V4xJfDFMK6cQCB48/CzU4q871MsBT1vXZOSKszxmTqrAfry6jrFSfG11Z
Ua8DrhuUGacpmUGs7SUvWkzR5bt6iHBrxzsbK+bSqJdco3s2es/HlV7ew3TOYHi6
7t5wMuIJIo272d4LgulOsSX4sYXWtzZUDIXwz56RCHxxFs0naohSJy0VPkzPEUuI
h5YDqF8h+T/O4spoJW96VpXkCYMG29TCrCcSy5KHxcoQqsXyECVLcgMpap5GEw6p
OwzAHDR7AfBnpDAHUTD18Gkc16fMF0RaEi68mNESaSs+S3vsPZYHltA8pu59WK0H
xNPzFVp/y82ijARHhQv2fVRzYuc1lha1RIXTK/YcGpZowcVi5yxC2k/QIlZ+3/v7
jzEUTMykivavKiN45bRdEzS8RqxF9HHtzc8THrwh1ilEvNQ2jDtnXgaTT/XoLr0m
Uwjn1i893ojG/TJbMOT8+41lqHHlWFppJs9eaCleB0HvrgJSAczkwiPo2DoZlZ2l
G7DqGrSgbgfQCGE+og2B1w7YDiYcGyZ76yO6c06EJhP/JiBMre1B3n3Ze60sGlRW
jgmUbp7p2VyRNGOV4iAOUSa0v6gXP8v8SrkdBx61pRCbQ9sEKbaT0jUtT2OvP+4P
PvIlUkbIxv1JvFQVkH6Sfv7A4q5pWimdCcOnFIo2Yt8RyDV4aAbF51W2bIOBM/vu
4g6oxybaZVLQsG8s2H7CrEvf+6NklboJ/OYfCloR659mZBVdPH/64FDmz9VuRVHR
+j+kPz3NKq9wDdEOyHujTExtN5mxxbKBfeAqoyEzWx+qZg3gMcezEH5LWY1Ug+mO
Jtqd0wY8aSZAMkEJnJOGpffx3XRkMk7umBRGzjuYl42awGJLifX4QepeGXchkYQ4
F7CgV+tAcLfovzKvRMAuOOazJmawUZk5zbJOsGKdQ2hwLzwr1JftE126wyQT4OCo
pfxmTtyaUJynjoSOWqia8Rd6mKVYrEpQVbxSkYt28X0Sfo9gTXJ4713lai2F3/di
pcfgf0eFikhGvPfGgutPhAyhPBhgrDXD08m9L8vvYdJbXQezeTq4GTEb4FR/9UXr
InJT9jvlmfY0g/GizNySnBqqhFainSviUV7KBhkVeBCjPmgopzyKQ/DxM0BQITV/
FW2RsWz/hiw7Lvst975hP7LOrhi+x9uwQPO61xOYU7mY1rvy+YV7nRKLnGtmeB3R
RbgV/KuUreY/lq+rofGrkg8P0NWUVVsDPu21tn5DfdlWPjZlHXfRZIsGHpiHbCks
ErOeQi8JJbIWEn4Yu+d+ru48EAXo1SZR5s29gz39ZmKMK21klhXaH/XHYJ29vOyp
fjFmjqDL0Laib8Qa0qpT0xgucEtPLB1cLCszwAf2ksk7VYaog5RS1dKpY8VJq8eY
tajWt0srJn/v1A8/qUry4fcIBVRDwnho9qoT7NAjsuE++wXKZjhDm0+0a6N/C9wQ
wQ2xgWhWtlNu1Lvho3GQfZCs/FIBRrJa9pn8AZuw/k2SdWkhmEJ+95cvLzp7YniI
f19xnWWBYrC0W97J+AYKaXBvX4o8B0V42ooo7FRJ2CyPimQprAUHrNh7oGkNVwTT
na11hFIOLIFSnbTUWcBYOrpz2Tpw49dfZ+W/NX3ETbPdHnAQBKTvwUv1HzxFQCY6
rwek1o5Ie+vDQoSmK78XtzubXKcV4DOS9T04UG60iV7yBg1cHc+OpPg4KnvklNCE
rx3WpNs1MwgMVL7dK5xURj9s9mtwlZN3ZG+VBlUTxKwML5FbuuLuRbEyYwFnsrnj
bKSyomkueq20c+1s1Mnko4S07UYuiekvo/hoe9biZg2quKpmPbc6MrgL6tyYF1Qa
GAOh5o+8X1NuqKkctGhvYlJXvvVZFS1wq/YxNe9WazbcCjv0aMy30eFu1fiEuV2u
AGF05mcU1G93wYkWwwj3cBwJgucPfCSGvAdApW0AR1y1D/XUAPW/LVp0p9XnGNWF
mbgEdf55KIF9NDTX8HNpiqKu1hOVkM9NoEcFtoTF530RSYGtxvjlKuUaWAR9V3wZ
T748N5UnYGAXFsM/D6UOQsCgFcb11MRn/nBKF4+JYSq0dyDXlnlaO72hEleN+2H9
nsp4KLuUFI73LMc3/uHWOTNeGgXGHyt6Pv+C2EDdDCMu8JXDYjBA8xREFdUVt/wu
m9sl/TnmMecuFEZIhwkQm3X6A8okDRlHvGeKUW1iyhXutHt8KKOOdQBHuVaW2TXF
yz0D/jKpYS00KrtJvzM8j4uJ8YjzlO+dsjvsBXnYwzXiMuJUsvrhstJP1jMuLBDZ
KnyoGRFKDF5QFFrYAOBmw4xEb4KjuK3zqeAFR86RP7cHtID0bq8eSVREO8d+EQ09
/6oTwLHjfne59hBSR94E0w5MFd+p4F/33GFZZTQIYNlSJ/aBBAOvmWDFyetdxtN9
TLIurVY98yFHhece9pGzkjNfff09JaPv6twDO404d9Wq4q3zTnovituspHOtV7TE
MgIYxR7tjWFVYj3VcvfZqOuDmSCKGUVpwYq6K6seQNyofftQxul7r8pO34uKmX+c
v4EMKn6F8s+3C7JWa86CzAs+aDJcprbT+gwuChpsZ2yz0sgHVoFg03W0E5t2F/8I
VLNHtnPlgTGwmHujr/CceU/tkwGGkpHldJf+jen3YbR6Bj85kWsczvfM6dxsd3Qg
J89p83mpCImFNVE3Xwf5dq7tCP11N3sY6p/UdV1EtupcS25sjhVKazxRUd7iG0Oz
7WBg45x+SS7pzpgk/JOpBr9VDCYlrRIAF8nkUHJWBL9tlwsMygeTllsgF4FY1FIk
46AXXZmj9Cy3TJX3DgG17KFZH7+X3rn4Sl3iwLX2gBG2eIcDkKm3PrKHJS2i2lkH
wwPjsmRcIdM39KRX3Sv9T/EeDJe/BXADC34xpi97sFtqtc30r9vCrdOKmawHXgG6
qQl2C7qimPxBRjoL/57zz7tqFG2DAvoYuvilmZNwwkhUAQ2b396XiqWZx2PqHdu/
S81Se/maTikLvDNi83e0OQaoBhbz8NxknFArov43iaUS/qQXHRN7kA5SQqE11ZV0
bBwBQRobY5zaT1vjE1FH5Asc2Lm9ljt/XPu8L9ST3aQU64IO8xJ44wVBZ8cWbe+U
8uydV8ocxiAaHy1nUxYLaUNldijP5fb8xM02SqhV5LxDsb9+OUkCl27E6TD5oaQL
gEvjdnzlsQDTHH7b9cBYh2J8mXpzvVNOBD9XkD+cEEF3S0gLMThMVduXobdhZ9oL
NlCPVpo3vjsxjF9FifqMIXoIkTuW78ob5dDohklwQXbC55DRIfDGOrVfJhPxn6sN
PpSsLihE06Spha9toBKSUpHh2/cccBaQtQKfJuaBjsiyKBHJfjXW305IDi5pxPnv
WgEj6dtmuXJ9wvybFhMd0ls5hdZitfoycxUBrGWkB30Z0JhWLjn97OBY1cOmC6Sb
LXarvHJdls7PncJI0gPDSHiusymGuSOGAVmMYCV6995uWALW4pRlpkJ2jVw9j+2l
2EVUV0ySelx8uiVfh4yhAiFwfAs1raIzcDq1wUeBccPz7lcqFrG5T/eFiHt6HpF7
gUJD44NMVN8B/x83uYplEDUZiGngILIK0jUlHcmuhNrGfJtZJEM9fsFmhBW94zU8
LqoUUFxuQmr7hPgGkBRhLKQb0Nr+v9AIgI3ivLh+w1WdWiYHBeQMKh/9cnaZswgc
ZG1Gl0Lyy2aOH77dX2NQbsaO+UYsbndfTUoaktkPUdOxYaJr2qBERasy0lPaeCCK
6yM6jl2w2CstEjbJQmKN546yOLpbKeeqnwUXphAFwbNbYxgZH4shPSNGYslp4cHW
l8L1m9KSshvTLEbU49O54Qc81sDyFq6gWdo4xSnxp5TBMOZsQkwaCNN1/fqtC2pR
HpRUUWcwlgACudcOgDNBEex1qKJb8uZxX+ZN3MJl0cPj2zdn6dq5Efp86d/5cJWF
InP7gMoMXRVCJh4rlnYG2IJkn+uRwWG5yDJHm5tzluHFD3s4arCwU4eECRGAR6Re
QcrXsVDAoi/85HjjD60Vg1uo1KoXduMQe9TvPVNiG3pwzg99Z3eP9JoCRrfqFCbN
9vgZs1DAt15ltviB6AmR3xV0Yg4l50+97KVu5PJ+tPw7ochYiH7IcOeUoMJQWJ4r
hbpD5Q51yTgrSrPm263d32Eqiom2YJQlmclKcQ4tZt3CHqrRCokaUNt9SGUFsKBj
kiRFtZhtPeGOpVpRQ7ogiwqtVxMfz0ZPzTOkrhXZBBWf5JgVKCE1gHpvrA+Dx86v
T1+FZFlfkgfJntZ+BJxX7QOJdz3Z8knW/7d+fWVXgROxL7DJOcUBiPelcLFASE5C
9qGU/KgvJr1aYQ1M7keKZr0oWTHhdVvBhQscBdDevpyCPAroAKeq3mvR9Ci1G4C1
sthY5zmjlGrAFPyef13Fh7UMSuwnJnF5VXhbe9ab5ygpXQgqoy6DNAHuaNzrD/Nu
/8UtB/UKiNMZYwU1x9uZJSKESVD4aJiVrdlnqTH1tj0YxhNsiDNZ9Zftg+Pkb9QP
Tpxf4dc1iwcRIj6RrYar+h+1qm3e4Z2FTGSv+TG3Sd/FiWQe9eenUSudCAqowXMn
MXFxy0utAGXGer0uQA70FnlH94j8U53OKLHUoXTJ2yRbxEYDeXZDKohJIzL36UNQ
eIhip6AsVJk63QGQzZbbT0yGSxazFDwIvVrfnRh/aT/udGegl1MXbdrNJp5B/TLu
yT5p9tBRGiq+fP0Z7mrRGJvNb4QzA3mm3CjFBzcptJkdijiVMSkEzGh2pTYWy/CP
CS1W0pxnNVmO9CUOdeAs5PurdnY7QZe4rMwinWFvxnmge03ou4dHDeKrYWSjOj6N
Lwp2C6B11OKWinjLFzN+zTDDeYliK8Hby+h1pOTauAZ4khnE/VoULuHEMwDz8VO/
Iu88LwFASLpwBGHFnUMEXpEMsGSFtQIkcOjXnorTCr9BYaD1RweTB2g6/YTLL56s
gKzvHTlYrWHuukdeB7TFng5Vou/c0cBWdEzKh1uIQTt7qIOyGVmlofAGTDFHYp9J
684HIaHhpscko18c9rUI4hM5CDdDg000M0nrAPaFa6pzzzcu/ub3wp05pq+imX0/
mE03mKpzSnF1y7G9zexGfigQ4SVqSTk0i8mAgYeKlHz0I++C5fmP+b/eCv7Z00D8
7jF2IMNyIgdoMfBTDVZvYpKtXhdjSOzfoMv3UkN/ZVYY6AAOBFTEtmJI3g3E47ov
/dF/TKl5xZiy1SHwnhyuKE6/XRkl6mJ0Qo3J/b3YQOOUzOiSkOhQ5fYmj90e/zsQ
u+c5VXPEZd0qIygYQV29rqHvndwfU7PSRkheJe4rm0SIdELT9KhFpm2nRR77wpzJ
pI7XFhIaQO+B7mk7pb6aLaMY5tnodzAaOyt7xsug8ajrhXjbl+mtTR+i7l9hOouY
1Fsxp5NYb6+6Bk+U6v3pAsfkPW342cCfBu8Z3TZYYzNp+UHqIl7KWHW9q9CQK0DR
+c/Qwn1x3rszPvvJB6b4D302/zDp/6DAQRwETe7WgftoXN3nvFKLkCWVquXeXhbw
KQUm6lV2lLIXDHD1EIUuZM6H7+UMem/ktkVfGoktxLMk3fUDJ2CZxyFGf/5EIBbU
mXQfyr6dTbk04Jds0pYvwZqdKoEpIBRKrH4TZP+6QVbpYgbdmQBQnnj/2zoFL5sH
UGxaxwlAvPuNz2kA6XSbi9MilC3RQmjg0ljG2wR3+uMCbxAAA+f6VlrrVy8ogKoJ
rJrt55HZlT9Tl/GPoawBpQViTsJC0DV0eN72wGHzVODDjj7i8+BiTF0s6sAkj536
nNHxIsIQLgM9uPMI3xE9J8aKzP0CkF38GsR0S8LRha+jCGWmcnvo1n6hJGkou5ZK
ouH8m1uZLtqolo9FDpdGZ96NYIcF+a7INjMtSheQNIT6KA5OeV4tZ1RJhvvJ42qp
iDDbYsWU+WnNtRvyXHCT8/jvK5oU/gVAXj8hFZz7d3/X8D1oSrPSs4M1Ax5iqPlJ
QOQr3JMKNq6u6i0g1ezgOMuv3qhNR2uDth9JOZKuvR8A1PqtvWx/8kU6z6ovATWh
ykB5iKYbK42WAPDpATZ/RULxWkFZs+zVHeUgy/NYIvSOLrg2tpn1UCXKMp4Kl9jn
by7LrQJ/ZbNmRJrIeX74QiRUGVyvpFJ+sApukAr+j68KxaorxDiO/xscKrYZpRGT
/PsVQsOX2pSrtSXlSTt67eWIxnVsF6SSXsORawQniRdJWV9voTZcj+F5aIfXmrk+
Cob9E+zq5B4UNUhVo0QneGtsxFrh4se9rM9cXj0C9k/Ayg2rC+tkwDcUtZaI9WpC
8eHW+YbLWnqWnvhGSyIw5CfN6N5kPu6sDBQSOp9urMMgNvFWa1W8STkFxcChWf/O
DxCoxvxVYkr4Rf7ngszS1jVtpESMvNogYefEKdBXFn4rXLrOu4M9RrbSmybhP3AZ
KnSLx16gyuZs9O2ByASZGlK3kVuWTE8xKL1BDiQqcnvNjITtPz97SWygxKte8y14
nFoYP3Sql4qEgiAJuGeCEq22g43y5mDnGNZ6I2RSaQp4pj8NUKql9zBzEATJdWPl
a7hEy4fntrEXq/CwVMTSJMT8p1kQZskbKcS2KP9vCTHfUxx+jTQ9aR/S26/GW8sK
ghRZE6owJLWX22R6LAddpP/FPqgp+u+x9LwQPJnTbCvq8MghsNeqa/cyW8iq53oh
b8kwvPMc9CdAZxdyMgMO3YkX2zp9NPmwBm/F5JkElfGlP9546Y29+GY/q/aguxJn
fUQlqf0WS78BLRpS/ZSShVPgVAaMshNZBjm4oDecNW/acoU0vf15Kk6rb2bj8lmO
F8mq8uX1/7NEUuLJrzFVBjnvIubukcyFomi8Gfl3ifcAQuDbmbrVM/dnajLX/adc
vnVhsVIP6u3YFgQH0AjFbROWzdFNH36i44z/EQmEumCbohGmK095G3E0AR6McNYH
S0yZt8LLOAzlGrkRJp/6WduYW3ElNTeZWoikJuwiaKTUi6UB9lEGm0ejD9iQ9Mcg
qU4+fOfykqmHFHEA7dbdmXcIuaQboWo8jv5n7MkvFA1zf/LrGTuGao+H5+QY2C2h
eEu0QZuO+UyfY7N6uzQuYy4oudMS7pfDBy4tKR9y48ZiMstFrOYL0Dzlm5QB6mAv
PTqUIrK//3Vhhl/x1OswSGIKKcFfKlhGfJwLCesKAmQlLcCDy18gj1F8xyfyVsiT
FKmXoMaLDvp5yRW6FVw7mk8nAC+u7uRcOEhHXc7WAn8sIsTLGoNk6U5/16YbK78W
slG5WDdjPI9po8sbYCwutzDmoJ5Ci9/EV3MmViAATJMCdyQVnwYvkP97VvPeHSNY
WKMIeuyRpaTcKM4x9j7LIENa9E0AIXyw30yW2YoP4BLXTZcn1TtoyfNZN16FGbjw
0BGThfC189AEkb3484mQD+Z5rlCHYb7TCUkiXJAyS2G3LHWwQiokkumSwirNoGcY
g/op6y7Hgz3CByEMXTM4DLsxfwq47JFfW7K4OBB033rPNhGZ1HesvKvphl40sWz5
9sWv0ngx1mOERfYDi/NDOGpdbNtIhN1PvYhzmLnWyxo6MonOWnMmZFCqYVJSDvya
54mmQBbWHNzWdjTy4Nmjov5lBkYx42K04zUsaskMQO8zmTqIk3YtTN7CX5Zqtd/k
B0wa/5I8mkoQ0USQM4IQXWxovsfLu8KIQFXGJyOdgElynipxhYlwAy6fzYJwhRQ+
kmG5AjDv2GMgjOF4VyT+8vJvVHHQP5fzRNsp64BKq5MJ8BkeNgfvqCs/a2+UTOCr
4BdqhGKXSDHZ7u/EsBa5GnQj7fxPbzZH5yAO0DVFlsxsiU/HYLjEXGZHWpNDwyox
F5p1vSmyZJ4tP06EKWZOnHfULguiGHBrcGIjouy9mu+ysfU57SCwypdmITuSftWv
nHRGApXVfMg9qPI0Hydu/iCXJfTL4XByAfahEu8sXyJai28/SqfwTDcWyIuhRIZT
T5NlM/XKrRtUdxJ/pZdllxhxUsCcdgMPlPPLlwdVNReqmlK08w+xMzSZqOGD1dKj
00nypTqeQwI0ae06Iess4mqRZYqoeXnasi7htZczi2JHnZwYpFcxfnNm4W5XDAEP
JF7URdjoLN6AJHny0VMi8+EM6xapQZaO5vAFoGt4dIyODLQQZXl06ROUisU1WQij
vXLOolcDjev6Hbc94WfyeCH6R7pOl8O1hnwrrrSkfvJCQM3XwP6v93kYZV2LlC5w
6pv2KUfmDq+fsXsrLPAvY70NiA6nhh05ahDu/Sg1W5mVtawFE0vTEz6YHzB0zZZq
azJ4QNoD2X6WGVaLFJF1JgpKvPTdz+VDI2XC009paAwiSP+vJXerRLkSW75FMKt2
YD/JT50VnWUiTe5W/LPHdYbSJEMH6HpjuPSwcne8HrFrVzMl3wyFgpBUigzGWlC4
2XjgbBIA5SayNEdxMBcUCFgYhnkf/VfYhLLYT/vzP6NnV7VlcTYBbZRIa/j2m2Dz
Uz9D2S0NOVVPeNdmxEnWmA+mv7CFPSQtf9ccn+hRCg+1+IVFqnOnDPch14O3+flQ
6jv1IJUpKH3d74LmJNGmIOd3a8Utzqjp6g5xTYNGr6z4DuW2xh2ym7jvBmRZRO+r
WdBLzoUkKrUViLHUAjUWcPDEqNQvnx0u2ohG8Gva3HFwKD+8sxowATUmRrlFsLBn
c9LT3B6UpRMGWtRYULaUAlzDva86BEppTwMn9CzoUQDf1EYUiTb3TPonxLMYEJ0c
8KCQz6DUiQ+LZ3IXtKOJ5eeIed6Y/1NUcZnDY0oijtJJGUdXed4F1sJWNpS2XwRN
7b+7sM60PmRTJOaDc1WyWynjgJIWB1aY1dDFUIYCrsOKyrvKCRVdTffM8YF8PUca
8xUyvfCMl223S/qoE1E6yoGFYYnXaxcveP3n2zs5WgBBcm8enSVRd6WfBxq7rmMW
6K6dY+9wnbHBLozKNioIyGnUXPgMQ45NHOBIti/qBBA7/8+jPsSwJ8jr+jstxerB
Gtr4WIgFQ/gS5cNygbFJjx3BUg5ks7R1omrpdqX43WosiMmFb4P7xNyPun4Z5b5h
Y3903TXrCtonBcXHM+EcSbK373mVi2qQtKhWNZ8Aaab6XKCVzZDc1nmrKMZvLHRV
CbWo+BTLPWSkT96F17oWlMo5NUCHBP6YdqxPnIlxJXbhQ0Cnaf02wVQcUiqsQ5aB
y/p/E7Z+Rw5o1oU5L0SZ0tFmV4mC5uZYKbE+V/1UAXMiWGdLPFZMncGef4BFoJdn
3/506SpEK8KS8M2//sTbImy1lxGIn/EZijzJ/tfhMNyNdMB8NGtzrywrz0ixiehW
MwTXLoZzuYQgysdmJ6Q05vkJ4cF1px8nmaBAXia3p18BDM5WwdHvK7LqBqaJDbFG
qjn1sH+JhBoisyPxFIKfhyxTJ5VSgRRNRq/7EkMfOD8PPuvjSqFsR1lgW/E0/X+1
CEkOSGiXPbBmbyF0Nw5KBbZ8uXThN3cOwVhUi4IS2T55EC6ovhdxhvNe8t33tFFE
VfDOVUlXnY3ZMx5tlGOw8wJHjKvz8WZIHePZ2V7lkvzM5iIvkMRajJ4nQcBMimDr
dGk8piOkIkQkYVhUYpyESgKW7hPKYVl75Cet0uPz42CJx9EgNinAcgw7xa13MgUK
ApCfXO+H3WFvwNNjeFzWI4AOGHylBHZj9q7uCeWUOW7lt0TTx6/qwtpa5b3C+2Ug
fgWwfOhlTfa8PUXCPGQwDDh8e0pug34EypDhOkbaCjt1KTezi3ap80Rhh+H+CVR3
FiW3wKaEBirQnVduEs1FGxbh8I1M/+THZfPEKjyWdc2knCqtlk2fEEVnETAiOzAn
o+a5NE5gEHbyz5C30DGuOuyeUCUTLN25oo0rmaIkjCt9fZA/UkygoBCJ7SLuJUx5
xpBt8GDmBB20lSGZv2YdUGN1remnNHeaFpupcPnlFygzSLB0Aj1KlGllz1Hbl0Lb
VanEmXBMxGbP2Ks9gBAxgfUTi1qOJwIfV2/pMCENYavCGNVzumw7JUQzOGUyNmyt
LTGkIiZl8jq9DlUE8563xv9eYoN2HrPjUWtRXO9cfNZiM3TNQq3zfAZi5YmgRhOP
wztj0NZR2YXkaPC8kOWhXg3vP4n+jrpswR01D+L2xIX/oxM5Eu7K61MKZF84oBL7
DES1DKjIo9itcxC3+y1UVEf7oELuFyTa1C84W5ZeBktL0oelxt2/usFuG1KMGNXn
ygWVw+WEMafpwKLSDa3HCt0VsuZGW7rh5w9wSb8aB7EAL+XQyJh/YE3N+TvnPgA+
fpseB1H13tLrEGdia+fKMPnqj18/7Z6Lh6ysV+zq54PGvw6/HISmJUYUffnSmEwG
KmEiw+rdLRPXPAddjta6J5mP4aN6+d7Tsa86ySul7vwVBESbsQvMlZypobFSJLlh
gJS3JNS0fG/fmx5xS6PXevzHxr+zPuWueIfiQyrAhPWd9PEWQhlY+zNXOFvIANP2
SSbfh5smFKtAn8Cic4lOSf4zB9yz4B3vX5A1pQMxBUGz/uk+pQZxWlpXcmOOdhh/
7JhSUc9nXBAuHCBzmwMl7gfMNoVaVx0OGkVb9G45gOGuBPGQSHvdXFyYgWN7fmSH
FpuoFUPDR1xi1SKppq4HfcUwASY6hPQSuX7n4BfwnKOC8f179dYvQ2PrQUNd7SYi
zU25j+Plt5VFrzP27kFLIk1t3Wg+DjLS98tLxdmBi0Q93IWqkPo7iAqCYSTvAjPw
tUQgDGyOOi1iNtt5YR+VtmDVnztdjSXlMHC7bvuLzK3Eoyrzesms9muOlmhEHEpN
akk1HmJeHwJg1E6m/FFMDOYkLCj9SWv2K30qZyvhZiZea/vsVgSO63v9n/vPokZ6
nbLL1E/VtWDfHwOmXj9LkEWjwMHk5MCJ1aThhir79pKH15jZkGTgg+XEWsrB1dle
Dld4hNGrcnfPh8paNr08DbZumcisn5Jt7SLs8m9NWhiD0lFR1bCD3YJSuMGkrNUf
wPJRc47csVMF5ttYmjN7It5QDNdYhVOlZlwCyos7+bWnfsww19hdyDkisuqdIoJh
c0BVc0643wxrqIRYsw12/K/1ZflzprV+u1Q/FCZXaT6r90JFqsgERnyNn0pwwxL1
7W8pEldiwJNT+XN3pxvaFs5HSJdoA6bDzH5JGymxopGzRei6BCoCXkoUdadGPRL4
sUfIfzOz/SKuAjqrDuy4ZaWEw79O1oRxUBS9QK8MwzS4FhDXqS2PeJxcnRi1cgws
pp87s8YjbgJ/hM5VBF0pmznWRB+VV5OOQyxEXDagqyC98/BfESoEAe/wKiUKzSMg
9gsLJi0R84YDp/Aupj0QYFO+/aALbQ+tMc7anMBCxTZ6mjCJKJQDutJWm/AQJ+yV
IFoirYso8wjPtxHGb17iUT3EHSGmnUoiUV/C5M1FHL8oGzy4mBgNjoc1yS8lJEL3
EUIHAp8UIDWNQZQiglt92vifERPu95Im95uyslKK87U6sJeVPXNJ2Ylgx+6kOtoq
FtYUt1x8mzb7TJ1IWF5ZtXw5mqdnYgWs5BcZ207WIAE5AsV42uKpWbAgsJppTcDN
LTrvO5jeaSNJlB3lfVC23hSgo5aY/ho6Ec6EiBRUUsRiEBiLfxnoAO/M+jRbAkb1
EKqO7LSaoLYmvAYAaMpva3f9KICvcbuS0u1dL2LujD0rwk6JMrYZX53A8RG0lolV
IX+t9n7HrWY3NMcM12gXIbjW7NP1PW2H7Lb8Gk4X2crmPW9JJqTY9vQpDlPa6oT7
IlG/XymvoNkc5xvILJSHgoWfU0hYtjOIgMRoig0t+qoxscHnze31nLbWGWW7Spr4
Q2wVIl5gO//u2oGFOqU/MPbIQL8vqhLt0j9Jg6/CklYDpLL+ah0A/ODLE/xawBHK
RIOKE4iGdiUd53QWcdliYmD1NRNLHTfepXX4rpDZyFKGjm+OGcU3Ic7HX68svkAi
0h0n+493OT3966DjfnVqWdwAAViizEro/OPSX5Px8uYNt7esSyVrf5LWK0kG7JmV
oOAKVnkJHPoDKvXJt5gZFk2aH/rMVYvOhQOc7yRbZowr92+thuYMQO1wZoga+nui
PBlx/buppJmV8wIRMIH/h5T5qD1jegJkX+gfbitp2P3bp3ropHH28i7j5x5/naLk
cuHN+cEyZ07i0pSTyI+l+yikYSXOPODDvnElVEgSQ8w7sS15lCcruS2sv2CFzrX+
P6mJH80v/pa5YdlIXn25X2fnvlqGoBr2tTUBHEnmV6ftyvSIzbRH3O6jB7qXp3uO
8offP4t7BYD95Tz5Bx1ZtBPXswvuDKnkjUPVN3xZEl6y2Sug30nRzBcHXHRKbI6I
d4dOKKCy9mgCEev8YkTWk/hz2nN9dpItpglceSAbqZbtO9u44hi3xEL0fpJ/9Lkg
llQTO+wBlVa8wYZx62kz/sCxm6WqC8xQ+IpRNZWrlpxiDXzpaIuxRZhvJogYCEUG
4hSrK3kDy7M3z+ZNub0M3kuTpU5fx167qQKZi+x3Owy4qwLPYUrXFU4FyRFTDi/U
VoJVCwveoyilwlYPlqCuP1wJRdCBjVdUXHzBQHnQgfziKm4vS36XJCAPDaF9I+eL
QU5FM5iKk4CYfX6K0rMUupun40L58zmxWn65nAVUue6uBM1YqUX85eBLq0HeGUhq
0/fdJsMsF/giNssGeLsTuK11XM5i6613sRWrgWI5c8bImBHlG8VXpm2hJtHvySmC
V23EL3hcCbJiZGuahXJvHG12lS/UV8LHbyLZPGl2OQRI4bN3yX/ApQSW+QDDZpsy
0O1p37gtMzykSsL7pwLooG4GjcJzqIs6NpTQaNnCGRIpx68/pWyljRP6JBfdrTyX
lDhNbGms45ZCvUo0trfW06eWsPjVbIDw0jdTlYH459lAoQ9FdLQMz9qeM69/BRPB
uMoc5nVsf9lS85gE32gXKHvEwDO71ApHOo40YSBUp4bwXHPDaI2U/lTdfTn6aNJL
/Cs5RlX+p1KQYPjQ1IP4Qdbe5G+bKRgXzvDW865Oj6bf+D3G47TSpRWqIsrnqY9U
wzLUtgtsUXoKWl1NjendsViV7L0NJM7LJiEoEsha+m3Nmkju4au/lqt0uzJCkrZM
wSJSZYgC/m0ocO22ZRPqcfE9ai+UkWNJIFe80yG3DvzIbH7OifiiOuHjxRhRvmiU
6sHGntDSaH1EuTQE+EHshOyvL83mlz7LDGPfUNZSuCkGDHOnJnc3ZWqJm1P6Vh6z
RvcGLoHF3usHl6zsRzv1VmjDEht/tIaEqHY3mZlJTGXwRgAkONnp/H8eLQKcJrxk
mLHydJm3lteD0GDVhAV5DSEWdapPe9YYGR0WwfsfL/UMnUpn/t/O9aA+St0lN32Q
9SDj9WQ0mNkCSKapkQYnsRdqJlhtqC+oAoSbHtb4WRHOknRHlf/kBt2c25GOfqro
ou6sZdUIrk6r14th/bX0s1oMB1m1M6K1GsCzILiJFvwoadkT6bHcz+41PjUc8Xbs
63XRnxrP5z0Xal8yZMES6XHFcjOvWQ467z4RqVam6fW7iNiLTXg3uCaxfkHrHQ3N
PiA/2WvwC51cqaZTqbzvZtFwAnAwJJjKbXmIcC1om8ROhrmIbvwScjo45D2vd45O
LoFd7zxz6AtD5w9s6zQHCHXNNm9BMExxNrVCI/hLH7uaD1euwLi4eKH4X84OiBO/
dmQYTbLQu6QdtaDlkj0yPK07qcG5WJufy9TwbNZQTBdHudxL/lapDAysXPRGK+as
GH5TGwiWqn8kVqnwUSv7Z5mFz7SJyav/JF6IDW48eaKbzHl8NDojJXUatcFSWsfz
JcYMxHh17DkUann3wyQgsvG5eq9QcuKTVPZQSEiXRT89OzaFvb0f4rma+X1boS41
+9VEccHAKiJbGcBYwtRKWZ4bA40HjD838Q/28cDqwu08RGlHkhGPZu89li8zAlxj
k9bv0mmfjgU71tWx1j2n0BwApTzBto50/m/7CfV6XR7FacXwP1DAj5o20BYz8gip
sc6HjNKS3jPs8Mtcx753PGfD68wJ0kPwChbgB2GV+ijnAlhnOSvxdsgr9FGdAlVA
LtCubSq4ZE1TXRIaAdcHQeyhbvKn1KuhprnpnPvprT13NNAq2G0sgPRr4Mmyji5E
TxPCvxcxxB/CXOuzpSWkmriFry8PjjkgPiEfz0iKBrjKKC1hJWuavWA89p684D1J
tmNrvYrlGMlmd/fXAaHcK+ISYHUvdnxvZFtG0+TvYKJGQDMYohy4qu3xk/vo9jTx
fwBMmPNCyoE+5ZXehmHmv60aSJ2+fR1TaksinliwUc0coO0tgdggriWmXFomrFWo
bvx7lgu+tDnlqW7dJOYYUmyuwmHO4fcIN3XLFe/DQAXfrvPebjzZzeeSJ+H1mNQQ
rL9TcHX5aAqvZKJLruj7GpBniys64q0HxszUpYnAIFmrhyWrcanSm8/8A3nTJfYz
kvo5f3z4KASnK4/f7M+GmSE0khg4EshZUFO5rzL188IVYpmps0QKmDfhwCfKuNfD
p/6xzus4omnSKXSKkaDmR5f7qWlZmSj8VlrwRHwEqr7040uVEDSHwbapSWoo+dbo
7OW5KawLgSLHQtgPSxi1wsyuPkZbGYmYj1od8XYlxtOYGNt5z8qizF8twI7wE1oG
6QllxNkZIlqWwIEB4q9pTHZF4R6n6Or2jYpfrH+SdtjQOT6uyfdiYuZJV9Y28k0W
QlKZB9fF0oYCOlJYYuYT9qrzuNxW/tYLx46ZfjIedP39HlygedPi8v/swpPVPznp
mFtd4X8eK+vXzbsCLIZzu+HywWGVDp1Hq/G38LXB0O/+d91pJ5N80Gd76hkic1UN
PI348wxIXDodRfpS15WJsIEzeMtK/6B0XKZEYRZKGcH8l4bXFCtHFT/b8BtTxfcu
HJjA+L6XX7eadOhrSuZ4KksOp38siX2gAlIhIfdnDAvlnm+kYE7QF5iDpl/TZfVJ
YaWXF0Nd4XIw/vtOIdiFbh9nl7Nvyabjm4Lrf/l2sAymKRWqUH/CoZI8Uw4qngKG
26IxQlHSP+Tu6VgXYeN1HjYFTb3ZYQ9n/L/0EOxi2GjKUoxTZtHZlKUfNpm98G7q
jCpYuTcOY+j+nw5dV+YRgDHBP5KR3EluAPzE6atdbreqELqFKBf2/rUmpy/PM2B3
PFjGHghE69q7f2h14+KNNbGXSNch2j86t40z6VteoFj47bKHplOF7GH4ConoDKVZ
Dr6Lwpz36bnLu4rw1ltIj1brFjVKQYYcsqJmtKPAY5Y02ryqHbYL7fav36GUigIF
WBB5lvymcu/KGRFnGKjy15diynaoVuqzBecNpbdyQy+HJSrg6njUYE238ZOm+1HG
N/xH2Lvpifa9XUKugPjT1A0eXNVAKlkG+T7d7Yz6f0pKWxMGxld2U8WE/CVbVbNl
LmtNdCrej66dL9WMfm3og8jxmSP+eleeOEfHSCT37XEW2y19/7qfSQaPgR/lXV7z
U9DGHsvRu/x/TDhtNdgEJa9FIiJDU09xczF5V6Esphk2Bz9CLG4CR/lLgBlpBX9O
5j3gIzdJHsWGv//qhAs5yPHVfyqGJyT8aevvpLlU0M7b5mtWpboiHMLa2ImFrbtQ
+gRN2hVXC9vj0x3N2ztGkOizc6wXoxRvlKMiLmSz5soij16sF6ppNYlvF2HJdCvb
unMGYpVgqLTgyU80Jv32VZf5yWy/CTxmISCQWepFDjo3OHy5uWUpi65+SOaUecVS
blVHWXgTCIkYnVTMQND6mlXgd4EbNIfAUSIYBEUTufxkKl9968eevkcDvZ3oasH8
UMohhFuJQYnPIpTYLq0sPsK3yooR54QoPM13PQ04qkUlz28Cm8tGgoPIhcnQ2XX0
r3XxKFRjpg6s1/iNhFH+kI1azLpVUN3iouq7KHJSQAIpfN+a7gFCOrMZS0oCy046
QlBjxIiG1aYjj3XxBDhkl/0fc3o/+lDPpOOZPpH+yaaWlnd5qhCAwrecQKEcY6XA
77JcdSSxGp7xbpP3LBQC8SUwSq3jZAJeNNA2H6/FsnPNrDG4dvqaHJPEWZb/ono2
Zh/gLXjvYm51OPAIxCR106gpU96g1aKWcn71orYrQ0t8xkd6NOEUwEfNwPjJRfUL
gsjzcDF99CxEj3kjHI0talRNGRFEoAbcAtt9++jlyxa7osbhqutfPYSfm059QUHw
AB8xp4XuYiEhgwB3BO6kcBUie1n3lLgDh9N5m/zru4M79XJZChm1GeoCRlH2Ud/O
6DhZF0BIEk2Ay8slmkZodFW8nAelDVi0UxQzVa1XMEA7POCaXCy2/ASs3Xs63Shl
r/2XN2/avVzEATfSdd22CCsH97TiEnSuwBcUloDM7YFdIkmT0vsvgh8xu18T8XFk
+wba4+pYPhDPN/hxRObNKnPfuuDpvrEIFa213AhOTTCpQGOeG9vX1RIQ+zvZOrrx
sfCBpUDn60EF+YAQqFb32eAC1JJRPZ5pmfFIlOquyspg+BFzOGbfeyWRSI69o3EA
mlEhIesrRUhOlf8hZTLh9g/FJIzsT3htMTif88qMIaNF9nQ1uiaQxd1O0R24xyTZ
38WJUOAkpjdYd81n8zyFBgLCXoS2ixySnXagjh4FCqlhkrCvXMCVxh6wgCLt7Lk1
iG5yZgdfPqaU97UwP1hPOAzhnKa6bV9CNyK27YG7irZDvUUev3/GfCqkIGtxtdNO
T2+wZyNvh2abxcz64+XWxhU+VN7u4Rl/9+fgRNX7Kr3M6oWQ2v1Rs5iZqnFA+8M0
f5M7trO5YX7V9oayMpoC++4Cr/MXc6eOUitjqTWmgayMFxoyZtfq46GJ17COvZkk
abalxa3P/dT5ojkNgzYqpZrMUCzxlbfmrevCyFaTwJGHPkHo7ICg3tXy81K4j2Me
hHUGbPHsD97jOjvXwgli1AS2T7f1ZxQjeEGuRDkMCg7V5xvpcQdjpU8DOes2mqpX
p4rZXUEqnoiZn/rTyMUbeCCscoHTXq3s7UYfZ86+5CbjW0CpkgyBomRAQd24xIst
M1HSeq6q+s07WlAV38uxbKx3f1RK6ylC0prIJlVLb49ya9ujoCkC1JaPidc3q2eY
HDGHunYDd4QcK4qvKdnb98wZ7R2Pv1FdbMzWJoaKdek19FGFouguZJuyjF8FvUKO
Li7Yj7RhhDGj6lx12DBfrVXkIOUfsCLia+zrCuL1eILqnzAT3Cog6UD10SyznpEX
c5m7KSbdgpyNh9324q2CFqPqAc/M3KTpmQr2Xwxqf0BeO9QO5ZFKlkCCU0BFkabf
x/7xpQH6NBX1lpLzaarcOINLaW0Qsha34n9CNqJI3LO/ih5CAKgMiEqMiLuYHXoI
cJ07TiVWHnDxsGtSc9346JvvSPSpkfLXPnjA1cOThqsj+8gWJXIRWI0VFxsQiOoq
kWvx53nek71lZhoTprNy1lp7R1P2+I0I4l6W2y44Y//cRBmv7OjY9bX8gTtRJYVi
pJnbbJiagj5W2CDudaWeVBOg4sgy/27wMvCjCYoRjUkQk5dpEXbYYNah4yE7BuZU
/iBpwlVeXrpVAPzfbIpKW5WA8ybDP5QZVDxal7QZyO2zZEyb/oLgPKR+HEJzQDed
B4e3JWdR25j5ygLVwGHOA9qDpu1etppNcBsxbKSpD1Dv8ZtFAsZ1y33uA2k6iv+A
n+7nRLZW2ZV9qeN13JkLpnqJKXIklztut/JBXyR4jTIQ+r9AIyXDna9v/N/alzzl
OJOC9JoGhmkfZ+46otbV1ac9jo2GHOWKexgdpV49nyjut6AX+h/BneSlC6UTtPam
NTO7vjTTZAySO2WHHNSKxF3EGB6wRc1Z4l/FGR/OXPtJgpjSkXIvvV971o1awCaG
/pJ2S/FbzNnpCaEOYkDxNCcUcDX/2AoxHWSLgGrYBZviK9wAce2uJziwAgeAlnVG
vmN11D08/dZU/QhUnBHzBk+EqE/OTrQdMTO3XQbgWUrPMggBzqTUYa7FjDA7URcj
9Rv4WJTlc+tNlx5c18lSJqNiUgORdsqKJKHAYXpszB0mhZau3wksjv2z8pMdaQqx
Vcnvc5Ta9ElxDrdKy/nQSLFR0ZNbLRXy2isMULqBbBmwxeN3AYik49t6aPC8pr0E
dXC058vCPoFWP6fwG5rV45ktx1KCHsa7f6r6ygDSd7dbAMK8bp8jtz2aB0g4Kk7A
HIJTQ7xafyblXiYQxgg/6LpVIxfsrBHYBuLsW6FpkWUhD5iEAQm6+Cr78CLMs+ze
MRYTfc2iWBKatFciC+aOJhtf9f8SCuExKlX9VsmtaYuqj5sXnJ8u2hSXwJ688t8U
voDDNV5fiopQITNOaRzsO+LVyoIShQ4JTglX60g/Ya1m2mqIyiRGWCTVFQcjgsDp
Tb1a83MSupVJfygsRJOtEnrD2XdZJul3VVTRNIgL8vsICk2U2MJ0mgZ7WVTQ7Ecr
tiqIHBbtviI9e+/5TWUWNVdhIh+Pf8N6eUTkVMYo9jcoG3jscm9F1q81Lu9H8Qft
HuGzwdcFSgBaeNFuPRxy9AHuOdZPvL1C+vUbBMjC37i6mgsM92YOT7Qfal60rIpQ
Yz9hSTkM1kFjExjAVgrm6OLAbUGCg8KiqZheu9Svz5oekvSfNIwCfGq47jkyWJPl
z+vpbbgXPPXpFvKMProTp7s1HkK6H4fbl+WI4YN3lORj+gAY5sWdjCJ3jbOFrkXX
k0YjMN3e13m2hVQKNcTfUrbpiE3/YwWjL8kas/bDq25o5LkYYalQz+uIjn+7zz44
VXiXYp3NtzwebmmEwZ097Apnks5sc8u1UjgJ9uKxsSZOUFoeGGbLRBAUMMKtb4ZI
mj5adpaz3AdlK33nexsXOffWAbFUykFhgn16dpzO05xAAYi/XCZ/hQmEtJd3K6RL
H/i2s+XC+IwQKVFvMyhkLOYurpq3tU5SlS6yQXEbLwHInnVkQZqzYjSa7NbLP7kM
GLMnkSjcdEAtlOYz8Ht5/a+fngsUf/4qrlGbeGlVMY8P0/2Xn8dcjiVL9jh+suIl
ELN5liTO0kLjrNUta/5fd1jt1Bozf1vnk2m+3vHLpEdLPwVBEUl3UkPnBT+gGsES
95hfOQc4GdoO8ovGT6uv57889oQcwjwn9Q41yyLV4eCfy72pwg16J3PNyT7/yxEa
hH3HSAVOdWoXyoxjMr+emK85DCFSc7gjWcJYY2e8gKm/B59RZtNix1NqeQpxEAvZ
yNRojU9dd69eJEI8395mSi7Rurh2+fqMnS0VTYgC4LuZbHRt2CyzY5duKbK8BlCY
h9gXCUl2w/AX6bUz0kfSLlKNzvqNFscsAuIEUgfwOic1ByC04LUjwFZb1dKAVbdt
2b9UfFGFCNnq/5S8EBflb37BPK2W7tHn27fHGUsNNJkmas1tQ5sg1ceq9WpdoGpQ
iN9NA6k7iXHoP3RYYEa2LD4wh5OJghhbPiO/aW0EfazMeNIiBjJ1GoaYhMWVdSiN
2bvYCad3XRSvGdH++mu2bu5/BNYOXW99T1NC78PNrh1mCGbzlx3U8GJF9ij1gta/
CUZA4H80Xf2pE2XY4cadnmf79PC6wP/nsc2n5z7uvTWpiKwVjYUQQf1+SKuMDNI0
b34F8jfJQK5wTSxYsoIdJXSOZOa+Lw3Tq7LJhogJvZkPUZdldp8r2V3szOgCI0t9
S65hwrJaoGmA0KQ8ORv0HBFBibPqt7mvp+DSPL6SxmsD/bwZGMG7OO2JdeqcVZA3
vQa1OC+GX7jS9BH/+DePGWJHaLCnFNcMrlep6JoUtEBxtQVud6evELLxr0oJoRKi
LZNjLoahC+0hhM3XAD+l6BWf1MdBjbX+LQhDpDY6dvyY29eQlCP3LZ87rka9AB4k
8UgeMFfwSYvrhexX5yDCJSg7uCc1rSuFIK/yxfPFaftMK1UOtpywfrijK+Rpuwo2
KL1xUCfUlPg1ybxLGGOCc++Q4hKUlCVQGncdt1xAxsZ88AOHDek1TaTzv1TKoVpe
jhKdNBojKjcXNodpI5HrevwZIn9c5rLOvXtpEykD6wsDcyek3Ggy2XlFhjB9MxXu
CVxuCtn0oJ+jYJM51WLkkb2Jl/5CA05e8cPnCiqtEXtt8FFz94LiFWXDYYHKTXuB
rkDzeUaTcDhMc6vW1IVdYR26R39kMkaXCTjJPgj6s0eFi4FXxA3tgrIbHSCG6Z23
fhF/pcpwzQyGs6fGgMNx4ohXbvxvHgAcay0zJ+x06DGEw1TOia/PWN98iDi4KX4m
QNJ5d7XdVHvlVMqF5u5a7uOekCMSRn2aWfVz12MR4j4fnc9GtpGmCdaZKXlx0hs9
xFQ0Gs/lU9m/lHWzn1nryFEDaxJAMaF7fLp7hNYYdxtAsrFPZywojRvH1ho35G4U
iqpoUXyYOUPwdv6hM9WOrm8GEuvRhHFS1pp5f8Mtldc5Qto0JKVxSoxgant2fwSe
dAGqrYfQwM4PaVK7pXbtcowVKmqR3P/+UDKuslI7o24aASjdpafOKZRueEu8aWGs
1xuX2FAxQnVATTS/5aI6A3PgggJuOayVlGVEFkfohB3D+cUtqdBVGKyfvIIeVVt+
9JV4xL/VgTOPsR8ZsoIjr+edeBA8Kxv1d+lezT8OvXFCekR/IvMsZKIZNQT2MG62
XgTho2WMvfOzroi8v/8hNreoiApINBlXTJEeoudJjV2wvBSOPemJc4UYdWDbzXXh
HG1F4CevhtVpOZK8QZVCNzIJ4pB1gS1YkQh9kJlQi7Pqesllsmf/+zYzxLO55SHw
H7i+OU8bDp8Jzt+d3aH+INUQufvH9o+okSLYQVFC7I49jeqjI1zpLB7IxNgrJAMM
dFgoe1U5Ez2SBLh1pcrUXns6ZUQVJdZZTf3gHNjy5Lht4Y/OQ33uvWH8Uc9JBPjE
4mA6q4XMREKmdXlQenmjbbG2DOZccN6ta87ljZSsB+rBkQpdPeZC87Vd7txUlqQU
8jlx5oN7bf6nhcxngCQMXjRgouztow3mwmHTYVpl5bhbejWMvAwTyTtHZpOi9QfZ
qcVqtXIMoKen0bM7aOcIklstM6gN3NaNYoTFbbO5riE1mvpizsJX9ULLADHQsyo1
xSDd3adrPF3Jo6/cexP6O/RNSBO2T8UBxdK/HqDlPUomjaRxSvglyWXIzk71w1vg
6MYmgooPUHlHhOVWyjvEpJh5Q0ebIxgXY770M3d3Tvj8ygFPdrbxyrmWtHrsiPXJ
u9HioKEcl5dmLmqDpU6yW472wq7/zWTJPsRcXejr7Lls4kaWhWih4rKkkgwZkJhJ
y4Z6HLQJ+Vu0+YBL7PGLJpGHUOmPaLo4mwdNKS9OLqvDa/ZGmmG4Wa8xkHwPefFf
oQ453TUr7OfZA88XpO3XabyPj3vjRD1VFKnGlh1uEoEyx90s2bAd12y9TtyH3gUr
9/R30Ijmb3fBv6tw1Jwl5VjLbI4W/274bIoePBU2RhqbQ1bp2LgqUea2YzB+11yg
cfq50Gv6e8Ck9zM2ZLO+sINYEelGv1pjkydFPWdfPfnIztgqWJAhbdYblM3AodLj
iVgL0WDTd59IdUGyTG4u/Vdbjj7xkOYpp6D4aUT1CKfCDHR5jQLyodhsv/LkpBlf
anrB+0fJk6IhVmQlyI7Z75mVl+x3PO7pXMBuxpWOAqHrRK5Bc3QVWrb6mwtJgoNw
2BE3HyLbwuKQpmb9Em8PkA2Ix0YM57/zRR/NudwDy1MNAWQC+iKIUe3UEWZg5aSR
4NM6b2x05R0O1JILvRCK1KzLhZp88VaZHmF1L/TgLLjLnIX6JWU3EovsaGdRlDUH
4vX7DW/ZLbWlkCxsAkgVcYSXOBffSq/wi+UfUsQ5LQm4GtSodkhVXeO35z1sIY2A
9H7dEYUSkhepvzY9Hs/3JdlAgnHXxr/iQjhDBoMlG8LKGxzRzO/12JxhTBls0qUe
cZNBkHHVgE1nM9h1isqMntYlbv3k2nYrH4YGFJeVLKvKh74nA5BRGqEZXsFnUfoB
mh4JEyiafDUNUoo+OUVi85Yd/ALrgVUHsK38S20Y9VzCL1cCfqraKY/bJLeoknSM
E47tFrMYLxlP3FZMn20QrIVTmcBGfJWQt8RJlG4t+YrNCvMQehDBt3ZNg0v39jB2
gVDL8RFyQMNUUUFZ78CxwlHWltof9gsGQEcm9jp0lxrpljXWv9h8nFAG0wHWViZX
cagS0XQ60Xl6i3Iw6HbmQZmuQTYpdcSriZ71Pc9DFGThbMmES3Ueq6yftbdCdv0K
o/WJej3ur2mlbdaHo3yVVwuu1cU2/PTWe/LfnrMZ832bObecgs+eID/lNjgOuxiA
qJJ8mzvUyOC8ZTAUskQN9q4pnasFxv7Zus7VVWapdDPzEjQS3v0ZV6KPiXMOXKHl
rBAjDBZ4bO1GqHjdcmS87zDEvoeX5UFWCyTcoAZmZk/pHt9Q+EY/Ca2UNxlYnToB
oB6tyk9S9XoeoweuboV7nCNs/JOKHGjIPuIxo3f0RL98pAae3sBx3k0CqI2kjBSw
qChnt/Qkx32yJv64iHxQLQmcyn/W0JXuFDMUSMpHeil7dJFOj+U4RofQIeQqvrVI
ScPUS62AhkkDMtKUwc6O5Zso3VMpeM8IUmr/rWt/qsAtdQNp6cXE1a/V/W6ijKci
LPwlVz075tk1qFxWTMJnIxOZolbgsLssBOy3aILZdaTU1U4PFqpGHvYW6CNJKZul
WMEBaqLg82Plvb4npelClPZ3cHecWyqtBpVoVWnA6J4xGb2302rJ9bUt/e5ih2qU
jdWt1IIt1agMQrl+odKPdN5hjfAf75OS7SaGKJe44V3c/j2H3UUebGOQB4Cut26Y
qQUWBmgDxvgI94gI61DjxE76Rg+9IYtg4oHbJztdmpFW269+D8FaggYiaog0N3aS
fOQZ35djYirsiI8GkkCPL6i6GlB442U4qVk6lAhHKsDkU5FPvuUN8LazCgUKqAP1
hAZy+NfQBC53wIkiDo1crzYKRCtapAfQNjfMTdRqp3BpKXLtYXCMhqPBw2UbFsAg
p6DFDo9DiZ5AXh+4ah+7Jwl4gd5OPQJSIjmpwYhkLyzAR0OUbAzGs6Gm0ZElSyCT
PEvQxlE68cUfeDQwF/L1jvMEwmG0R3d/v05IGSqD9LBmvN/9lJU1/OwHgBIgQJWh
XHkaQhRFIevxgu5/Y3oO50W3wpKW59FJLGMVz9dn1zgNKgf+xCfObmix0Zk3gUke
feuCqyuf1TH1+t50T1uo3COVIaQAwvBMa74EzJsHtdweETLBIVzgx3SZNwbYiP/L
4hAFvhXAxGYeZctZjVbJIqu9DqgOEMLFTUloXaAnU2Z3uqoqIiQ9t6mkSDaoigXF
lVuMWYrc0K+fms34+2pKVLYG5hJ8yz23bTaNZe8lXRd3IhhOVRuCu0/QJ+b0cf48
7p0WiTni+pvhTn9LqxUGDg5NVCr8uKYdWHfygxEenDfbyvZZSKGO/LzVF26w6XGx
gJpRQmHYf8qj3R6dege5s1588Kf6uFBFdCJlFLPbk38Z4SNz411hQrJW7SheELoY
Sb5EOA6WOHpDA6AfdnCWg+dLGb2rvfjremOU3kHDJO4JTGkZTBMEKgThxErpj4nz
Dae6+0OtWC3INh47tzgW6YMoHLNTzDdniPYTPIEfpGPnLz07GOLBgUXS6GcQR8ju
jX0Aw/UigMWP4oMVPlEKQyNTzeNl2SKxml2E2RQmBdoMz4a/302LtpDb/gijDvSO
m5R+ofODUCaps4p7tqv2I/EMcY+cJLknZN2ngeGSpShik/T37UYmVlncILRgFZCF
MibWV/gScjT7vCDrk0VpTEVFT0Zx9Z47vV0AUixEJExzNGygPEZMLZRJ/q1oKVMw
XCCYPmDZ7e62unptc0+pPu/pkknQ5XmiyuMq558HfxEbzCFWLdhhA21FgP5vPpB9
ptKSx9E0agtEXqaf4V29TjdK7K+b+cSVTLpREiQrxDtlg9AC8ZctBt6RaBhSOtD1
hiRqrSBFKi9/ZTASCoMPBpUHO19Jah/wFlqMDbAAn4QNtxZ+7wgSjKgR8kOcMyq4
qTjAGdNRcHc+KacEJnUM/xTzEPGAhmeejQb6UjwiCkN40Sd4T0ZEg7J5oXg4VJe7
GvodBEUUIe6A+UskKo5QeYfyWsv3u2qkMTvmbDFrvUoSPQU7yrTZlNdRhZ9rmhgz
9epDsKjgXDA1un/mB+F42ztvAA2vRSaK6on5MjAPRL7r10NRhOSIWlL47D/Jgjfs
wYNI2AOB+o97Bv6EfdPnvP3a+WFAaZ/8Hts20f/I3lIrah8Aip+T10Qm+Q9X5tKU
klJwtoNKeltJ2lGSWXJ5/JPRJeLEIzV0lnLKj4o7WHems5xXe5dUmdSvvKYQu1sf
/X4w5XeX8nqV0EKexYJbubISC3d1iK9bHZ9uqEw0nsSfgElf/Pcf+EVZea6BwWwu
ETQkSSp8j/nZinw0OT6jEyQ+T1NGcl46ktk2CitJXZBGTWPA+BrMpS9IOSdKEbH8
tNAxciNlUz8EDD7bNtU1ko0W1/xRqtID/sTUFXlR21s92l003wQnQYUMNlgvRYWW
zjc82EWJ5fTEZZOyjZ7LgMFb6eQfCFT/0WmpboXwz6cOZaAGILSgJa0U1Buy62o8
31wfcCUg+nksp+hmxl7gEVU6WOCMsgarFs8dSd7EHIOy5eYRBwEzTQEhSSzDxirM
6lf0suyaPz7rODaVYwP9o7aAmnJWvfbmJM+JxnKnvVkEST/RqzkeOSMB/f1rqdP5
F3C+ZZMaulq/N880m/j8Gbd+S9gfTZhu1ovDX2EI5We9sDTAdsYvV21Sqbn/tZXN
mX6RXg4zexONWU9uudSzECT1Fm+/6fty3xwiTgzHINaCYclIU20DV0KVid9jr012
zV65yyPFwiSTtXCjI1r738RAVD+LeKB7jGCvxYRDd2CtxlGo2C0LYGd+dpHrh8pL
t2VybbAPApvYbNXJUA1iMgs9rqu9iyiAJ5YzwnS4n3Xt1f+RoA62iEyUdkZKO1cP
xW+slRiyiGKsNL9TC6AQ7uf+EOy9N083zZp9uyPC2JFC7XWI09oDcS1/QzrXfwvw
mAk/PHW7jR/XvUmTMGkyjCQYMb7HVCF01M7gfB9tUZfVcoVkqS4NV6ZE0ljNnOLe
+DISeBEZYaDp5E4RR5GSk0NmqV39+8jLTf7ytYU8ik4bQRApyuxkBAJaUfYlRi61
V+NHau2vGnwnLbelT83rO53jYrrEYyInvKVE4Omp+TbbK++z7JW9PzZGUPLpYSsi
IH/YPq/LyZWrWK9koUcI3qavxt9pbnx2ChgA3vrAE9byKSYkiXFU7je28dL+NSzM
CeZituwBja59RW0OoXYqdgoTb9NL4xras+7kJYjzksE3md0R6q1GnSORVBSzY4t8
UfTuNoi2RkxyFFwqNyZWqRP0bJCmF8iWYX32VAsoEJN6QGCxYwqw4vRUx99BX4Kt
Awi58+uU92ziVL2+/pbxogyHAm4Jc2/WEXn1rto2D2dZzpyYeP0K65ILhCqqXjfw
ivTsdYs0vQL/Vg77WOJQpdVkFbUupVpl+m3AQBwqh7Q1TyI99ltK3U0xYnxwUP6J
BBWBa1GLjMISWXqOkRuwBA==
`protect end_protected