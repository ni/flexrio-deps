`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRmRy9l4xs0tB8DLo+i6+lxmZYzbZylZkJdfpQ1QH318T
WITs12S2znaVMaxiQ0esp/5qpHDSskDhRML5GRAKcX03Uru6RpHzVdPatAHyk7kL
x8wSRsPVMUtHHA4MbLFxv+fsDiyG73muxsr7klH5KGX96jVapDQji9xjBz4RlZbf
mWD2nmbhabHcSguet6jujNTg4uqLzbBhAWqFPeM0q886CCt5vgYwZeqTPow3Nz20
d/6zx02nyLN6s4sciR9JH0clp5cRTzqJvszaCghpNuXQmR1DY+BLFga1352oO3RI
k7duAKhgRkVgWF8gE1uqzJAIeiRL6ls+2nIzt4nWyR55vcxBd/y4qUKULiGhDOAP
nA8dkywRVZ0UWgJ4SsbGzOLDC7PT6ZH7qL0cpC832nKadcRHqn3qT6AHIaNpiW6+
ExFGT/WK4n3ut47MFmv4UVcHYBcauWXltfQfvRZQQj+1IXIpS6jFcPnEa6GuJDfJ
5WoG6OlHylf+iTBNVLi1zLCCKcEbrUX9TlKBflP1h7EZjDvJpquWSrfbAWYhUdDp
vhS6t0CnhZE9ysQnDh4TGGTCqjLptCiDQwBvS+zkQvDWosIV5AUfKeAasN6qQCmY
LOnc2+1JZlweJ1HQk3VeOwIm++3Lu2aG7/KQLQb/pF+3XiVmZJdaIrcOgm8iw6UF
HFYegTQXyn9xUFqlxFQ4kZdAggDeUHNZw93aO3l4si3lYgTmSNZ5SaozA5wkuG+6
okifOfbDmc7wLUZ30yaohDDa8JSkrTsvsz9GA8NsOk/vQ07jZum8OQioQCNPm0qp
MRDeJTgZdDxZuVdXz5XfuQQ/g5/JG01KusYaIYdY/lkjOo30K38y5zrCpA0jMvOn
tf+wGXqYfxq8YWsYLZ6LI/iaBVrDWvXq+LgOsD54JDltoUhUKASlAN+lfO6xHmKx
nS8Wv1kWQqUAXTYwSTPGTvGrO3WeTeBWgIK6l+KOy2p7sexFQGLGaPNJivOX7mpg
8VCKLggopdLHgywA7iV1huJwJvCJSD7FxODYspIUGVhpSJtHYW1/fK008y2pK0hw
eWwCY5X/eCgb7meMUvArNi74tRRn9d10foGpkKCqtBYfdBoFodZldWASGxtLzjM4
meGjxZc4lJTOOvyvaj3NDMbENVQwzKGSDaQoa/ya80X9oUfsuUF/Olpi084WIzqT
qwSWGKAVrd7zZYZKKLYvMB4xhpwztfiEIpbJ8TIgbaP7xTPn7o/r6iM1rGSX2DI+
beyR2mroNnL8LwAFFHM6fklyqHxwkGt1LiXW7QrmmJe+NoTGSOZAlksQu38rN3gI
PcqRBjVRQcKpHWaWqrzizq3xNOYLfpXEYY6Gzn9k8s775yPRyVomnubOx9HUi/3z
GduyB9GX8v9iFuKj2nUaBtUpPO4TW4sn3HrkTzE+53qMFf5suM70KGK8h3/2nJC1
NYz3gFPG4PS7pcs4mtoHSix8MTmGh4te7Uv47Os0SeB9gvtNCsEEYB5Hs8UHzwh7
SCg+2OHNac2cqnL0jgY5Xa4Y2WhSOiIphHfFu5S1e20AIBidv08bEK+h+pPD0iSs
pwLAArpLjuL4SBlPw1NRmlNKFaBsiwg1kKIpyBKg21zs+I1eT0iNm+GnZ5K4YQ9Z
UGQUl9SfXGfcy+ys0gAhiHYjNczkHok7Oy2Fo5Cff7yKtpp3uaigWyRMND+7abMf
KIBY1mjIY/d2dXSuabpOvMKinRivte4bifvug+jRPapcH1SIHbii1B8NQd01Hcg7
BnBzvm7ImHidrtE2UCINiSyhRvcSwwgeCMAB+bdNh0GHwbyrTUqe92MX8xGLP1hM
aQMfptJsSwtAy2waM1ZpArj5yM2dPe92nvzSQkt4DBSS3zVQol0da/pvEruV3t+z
XFN6BkdpYbuqfNpsIB+/26co++puQbXNsFHRvsqhOAvRFCQkHNFwlOhtkejmSoHR
uRVEZ+u17xl2auhbAhnVhXs4zrqY9gj5/Gfl075EWeSovZVmxB4XUmpvbrTQtG+o
jFa28uJA8aBcZ7XPv1FJFAE0xVIcJvy4afTwg3pkCTWq+5lqD3b+CiGqwlPiJ98f
50dL5r/TK6WWz9H417kqBQZIKxo5tX1tCQRc0O3BZ+9Qwjh8VfooX18p2ZU+/WQM
e66vA95td+JJ/q8zD/GN9aY+hGpAak1xV3ad/HiyMlvBdmGu0D9mUHjtCuPseKzi
0Tr+wnFK3h6b57NXq1q1PY+t4QqgwjVbfkBv7cApEcUb6wCgLLHSqE7vrchZLev/
z0U1pobCHjBKx9/KGJHPmZ9u6K0V70q+2isMQUDWbgwInwmxtLxXk5JaFYAH0TXh
SWDwZvZ1h08TJT7fUW1yAiuykPRNz/5NeY9IcpOsKAlQ1r6H5cYvneMJiuLMCg5f
2z1ifvoYHjrcl6XluN8c6O6eHQjVsOkXI87abiYqlebQv7BV+UfBBv1zI7uXpXzv
l81k08TDB4d3hxXNE1ybIHR6sfP3SxOI3W4fr3wHh+tNeWi0gJF+Oj6HTiXlaqE9
P4LECrxtaush9jh8lIw4AEWjvJz/Jg6PyaQRFs78fqbFDr2LBwVHRMnJluH/qKjx
ShNcICvGcFAIXhecmo8GqcPeUFv674rhRkA7ZkZRINRssn2Rqlmc7ff0rcnzfeK5
8EogcFq2CNkB7+0fPt/5MjNgKj+czPVetgfxR2VxDuOEB5u4OpvcVf5b4AvVFgfx
qjjkv6nvACFfujN2o9OH2CeohE3Qq34mHOtmVJeMYGn1fZuaV9A80wc3RyhKb3k9
fBoyGXkl7dWVEBTaongnfWsxuR0mpNxl/OqrpGHqzXhVqIiOUYsD1uv4ETxaGTwR
7K531cDwBQHYj0LOG87gbntXGm6ls3W+tpzv+9dBJhY6clF8TPllkxePDkyha2kr
tPpcTWigYjlotLhyoip26zmUybyq1ewJOsYyV8SywcLXOX4/ckH4QLZhsiX/scgj
8hpvWuJmbdb6w+3MmoRktLWj+BRX6NmJN+5TmqVlHX5XCUQIPUl7vnrLNvrR21Oi
mte8SjMWbu8/N2oj39MNnMDR86dvddT05aiIZwSlRAtYcoRZpmrKddHm0hoIJAZ9
q327a9isI84fffZCa2iSOA4JTJyRoPm+kDBTTFijsA9APQ2HXMnugEwgfC3/tetq
UZpP1ghqehrloKMZdqHTPRG2KwKc3RDag1xIHZrFHQelZ2CZNnVg0N9XNJhoQoMM
NicSd/JMy9uSBp/V1bGRXmW3S8hA1j+jmZh6oKcdaTmFKA2Ur7oQALro93tlL7R8
TrpKflxV7dFLoCBOX9jZgig7n6TfucMu5+yWf7mWVD87YxBFyCYSlM4h3cgk9cjo
yFquhG4pjL0nSdFUVgaxESzovyMeMkNAazwterp5iF3/p3atQZpRZTaxCVyTva50
I7LLVhVO0gZpYhj8TpCfL3j8/alGfCbcrDNobBXE+Zcq20Wj0fl0fcwA7QqYyunU
FivzNNQm0OjJvhczmW5kYE2r5oaWO/fyFmvATyAqtKVm+mi336ZMqFsTkIBcrBWU
a5OQOoinfnN/bV1uoiItSX6wvqN8YMY06xGq+/8qISpBShQqpL9W2PsSWpmQdjMa
upCg06m5J4uenEpZ04J89DY6BUC6Lm5qPtrOW76rgu0iIUnVM7cYhr/I5V718UXK
Hwc83MY2KbgyHKbbyBOK13Op8n4znjQdhHwBkbORwUqHQ5QZcas52UXgDWfqi9KK
WmwoKsWyvR5lGy12TDPkd5hOU32vHmIkoxguie1Ky3frlTQXEUBYYxKumSQErh+m
AZq2UjOXk6hxiIZEZb5z7z4uxC5nHODqSiGTW5qXAtEI8cM4W0Pvk/Wjs6eFRDAy
vc/OHAaBFQ0u9XNq3ywPyF3r+cmNdVWoJSARZnoyaZBhy2Cn5sDS3pwMsJUemh7S
+BjqmkWC0r4Y+K77IVxgc5WbhxqAnM7ROClmvlNSZBIrTcv0r0xK+i4nxNYUbPk1
3aVJkR4vUpFFbN3PxT0T8NpyvHScyGsOo0xP6BE7vB+7VYt1LdeQIVhk83Z6G6rc
B11sYl8cRyQf3qAPyaPWWO8Lt9fMt+zeMntzeh/yqDjL2RfHCDZZ5ZiofeEMO1vQ
Sx07Gia3cYsUErAkTCsXsH4ITuXBiqYVGu6dpNC3fZb9r1yPCkqFG8NwECnoZ/FA
tE6iDb/XP0uRfkCHPCBVaZT0MS822LPPDB3lQIwF6kXl7bJGUn9BMhq+U5BGnOTa
m9LAtkiiPSmu4W46Ss1bHjFJHLUPzAJwf2hEz8+23X3NcvcCu1CMELcF+AXSZL62
VkJOOk/zATSKYEpS1GfO0FHzJzWfk/AyKg3N8FGeLIvcmNe6ir7FOYVycJRWKWUX
+LaoYdXlsq+knZ6l+DJlZm2piJ+X9fZZ0Q+hMjncO226zkQ1TgPCcB1YRHUgaIon
scDOlb3FiFWmYAlUvoQhwFiT8ugdMHSCChpzFdQvHfGh9nl6stXkks5WhKucLj6E
kYhxa7QgMxTAKvXWjefoufTUF6E1e5pFVneBOysLbE2Z4bm3ta4dcKSTuv0cEZ5y
wOVGZU8cA66comQLkTnS5T9/mTWyyMf7qzBFExzXXBPEKneeIeJyW7odh1TOt5yp
rC6cTJQL/8F36tg5edVdqVZejtCgaFL7b2CZSC/AlDXlVSo+FfGBWxmRnkEkt01E
fPq7qEtuZLOYbAglTYDMYcaxSuSHPh14hZwWfzedEG6ODkR5mSDwowi02DLEL6f4
6MUrRcHDDOM/bWH72PxJSWsZRw4D3v9dC6XOYyuDcEUXc3PHSLft0HIJ9QO06UDZ
gEIPp/ud6S9cTEfD8/mjiCVIFT07SzSBWkPNq60xK4yGVYTa/18dZBXQs+JS9/aE
6qI3FamCB7eTl8ybVQtl53aDSqOm3xmXsfyPGBw78SW0u3vXhV4tWbE7g1pWdYmY
vmQIO9E6hyiJgCoAS8RUvDvffqqSS79JNOxkuHm8lIC5qv32paL2ZCN60v0mAiXV
X81kg5qEvI2uT6NFSq7H8t4g0OIbbKa9YDceqSb/nUHiaV9yqtUAP3OYbA+4HF44
pyh4nkCDklMRZyOMDbXDdCXa0ZXdROkZFo/LF+FnB9VHAuXqARcejG20oPQKJWm8
vztGKmahocEV/skyBId+I/u1rtAYTlRF8PJrTEJR+L7IGnchLtpe5UD1ptmy2Gkw
NFhD+8LDVqSed0u1wgvTJdWTJ/t1IpbKHr3whpY0wnmzDLzxHHAgm3yBC3wxjkNy
qQ5ONclJIrtUboQ6xWFuJD8ufgDARAqQTkEIr5XUs557BSI+7l0WTxvWbwzKiKO8
DhagyrHLQ5gmPdZmTzftwuXX9oAYkoZluyDAsgUgaKMzCqJMFQ1Y7HiYI4vCooIi
lU3cLig8+C5bYyXS2Ssr63FqlWuyaNvpdNORXdjC2O1qqqdUD+3cK6w674FxtzE8
j4v+Mp26Y4jVpXA8poDGwT6fJGkFXMMmjT8CDoIKw87I9SWZpwBgffM8dhji07ZV
mL8ZlQxo7UmmUy++6LqRMoKWvWw27N0/hBwLy6HSW2lvd9ii4XJg0nuEOrqJo1Wf
ORu1Z1DRWVBQinsjF6vERVNA/7CQTtRZOVmMhMMqv0JHvPYw7M/2WvD7KxIhCdt5
yJJ7uyEQkBeVV+V4+RrSwnQ0oDIUbSDcIC5gAFg4RGm5wJf2v1S0wy9nm/ZveaGV
Jn2CFdxE748crYn5VkkrOkLadFtsUPo0hvccv0FE1XozGtAdnzYRO25Ryu4C3RNe
e7aPVZFqNzBJ3e29pB7njOnzBzsWwu+mPQ5aLpkP81kGSsmAF2I8zyA2CqbME2OF
HsIfKaKvVNhonUu6ZaCqDRG1VWfyiFYrVkEGaA+KXTYDAZEhrCKWgA+yURBEUCq8
41ub2RSL/PYIqrvsVsa3wDofHa3MF1KMCna/X8twjTe6vK5jAlmoltp3fBz0fQgs
dDoS8q1dbVcQmhY4Q1GwtHniAulkWUpOi3GMTH5XXgkRPgoTxYkN5KnCbMytuN7i
Q1mQW5yFec4uqz9UOsnFn6NIaAPs4ul/JhCWPO6zmIs6Snwcp75SXuj6deGDGb9T
LfEBn/A6raE1lRSU7ffOPG9BHXuLyr5Fe4MM5llSU5D/VCMTAMth0CSXL6xRtkF9
aUlC1aRao7oZosZ6wk+HMVO9vhSH9xirg6iTsYFl7Jjiw0RWBOm7I+f/K+30v0rg
xheWGICib3sL07hnDK69tHMHUbD8se/3LtBNQdjpz0o3jwioXhNIH2ieH8wRwAgU
Q6mfdAUrbVpc8D8elhFS77yF8cSjDkKLLzjmLCGTzXUTsvET7n4ZlUvo9bMCOFnu
447PPnmbczvg1cH747rXD8U1IknuZGTDD+BJJWcCqwMcDdBM99ir5OGKpyRLsSUu
8e5tQmkY4hvj4/JRuUWdjH51c9zF9rve+lCmB+MclPc+dHiEG6IfNNmeIb+HFfQ/
C6I9DSnzpQYCINORQFoSvs74oyco1zYCN/iUsExvU0y28jx/YrwV9+OIdkEES8Jd
XjubFb6dSk+z3iGd/byZBQ7SXfNx+6/mZRtnx2h55H6JB1iTaUUBsOkYPM2fm9UD
dPjT5Y5tu+b2NSzmPIIJBlmhSR/mvcHInwzUii4V3TrQV2ajbpscFlXGKc/kdAa6
cDP76dKlI7rSWqN2fjX54OuvRe5ntvVJUZcQGbcM1XqdKS87S8pZbpl5EvKKpqkb
Y1B9jeQRaXcpGz2dzeCdTUL46rMzFPywhGcPUQA5KIE3C4SW7p0G1VqGce3/mwW5
9mPPJLp2cV0jNZEbT0Dkm2sr9ExJzvlssUagcX6Tb1rxgmsbEgUDdFzJnfpMSf3B
WQZ44bL3alD9DEwxIKweDv8Zsda4D7maV9P0hCGuYTb4rHJFtaPmgU6i50C41NwP
vVlFFfPw9dSOaJzMiJ27fqbEWk8hCtpLBK71JGqb3Fqf46eI54z815x9GGwbvIZb
m25YqnLv743rJWpRJCV6kf/N8AP95fCfGTe3HrlJdsOgrDfBMTBuB9nr5OiqszKn
ckqVXv8t+eyIar8zx9cRWRtklcuvhS8ybE0oLpJDvcJdKtVFosUaWLBSwzxMEvE9
2/gkXxukjigZ7JVS9bExynNTgeEU1baSRcJ+Zq40ViZp/MutPaVGHZyKuvcatUnr
sn9bNgZuG7hHFKiqXr2GFgYSVfbn1qPEoSzSjfjqFuN99Mt4vwOpfOA5jN8v08wR
OdQ/4K4aNTPHRmvCMPSgIBsk4p9wj0wmw3KmE2uVIddip7RAD+rx0TW94hU8Wdor
55VYu0N+12XW6xYvK2gfgkKdMqhg15MTWnFWfCuwVjRAQVV0gmXNXOGE283NwRcA
dmPvnWb4fgiVScFNPkU1Hq9yidsHExc4blSXWfiOpO+PIAtJRb68Rru9u2HLP8RL
9fKmx43WTFq8/7KV1qMM5SxMtN3LpGUJaDKcktF5eILHLQo4ZMs5MQCogLjyLtFH
aXVGS2f+ALj84Ks2ygEXHqMjDDoW5oV0g5LtjQ2C4JUwOg35U0GGKJllIZtfbN/N
NNcgbe79+SlLYADv7IOeX/oBT5m6EG1yNwYGL8uuY+98tPZpsqCMnBPWhXun2+l2
UbL+RO15kZoewA6Apo99lJajfUTKAiuj/GfONAzMJHQD1J1+fwhwBEp4Ud07Zdwk
nkjizEaGZ6uWZcxpG4vWtXvx65wHWDjbfec03F5X62LLvaYGsFR1ByPHMJk1IKV3
z0d4etWpg9SOrbMnWKIFBmf902nJKy6+arnXZFp8T/FKJdlSk/ghW6oQL4B8QDpw
ztQeKWCKZEpaTs1Q4iHxgn+nEm02PAp0b4P6vTv05FTirz6B+467R5leUal634Bg
ObxyVVDDNZOkjsd2d6QOxkevHNkw1/Bc0kyTQSpBuql+ph99dy/IHkb1qZ1FR0E0
Mgc8hJdJa/60fS4v0+RGKCtdLpj0983PcMB7OKfs1MtEJTyWU5hDHkrQcy8joCGC
MYkUNO6ZxuZIyHecqwv5aRVQDSe7A3oOoFQwy9edgdSmidzRsYhtBHs9m+jEUhnR
BLGZdq+rFWOxTmLa9VMaVoHqOeBz3xHSK1bOT/K2a5YHTrlQB+Yl9Pmd0gvCWJ3m
sNHZ/C/82UL0YKyit4dsOd6QRFWhYOgUk7A+Uga2qdqfdV0qf6dmj/RAB42ELs9/
NS2oo9/2s8gd5w+ttNvP0qvqNdJHhxuUy7BSHQb8Cz/rYCW4LwLH09uVFGGDO52b
96o5LZy9H+1kug2roiMXeMJgEWH0lV2/DUZx9ztX80XWqEkTh2FyWWNt3/Aq+VAO
CySO9dn1Hd5b44KeARMVsB1g/TVs9UMMckMULrrEuG4Zg/YosZG8NytruQj0N6m/
y+TY7jb1uDDhp3BKuafdfoH7DhbJm7Jq+bBiqotKH+ExBoZUHH6voKTn5ryR/S6O
drFK4+DMLr49Y/R9FZ8u3dWSShqKFDYBhRyOnfLCClFuW4PBTJxCRKJNOiBmCDaw
CGNnI8wZ5XAVGkmdWs+4wsX+g8mBP33HMBnhDZKrK3JO6v7ljJmMWKfzPKRyQOZE
ddOrTPlBp5b2oet+Sh/ALVYAg2rUo+IrvBzIfYiI5S0Tu39tjnoTpdLN3ee941km
wujXB2XQWHaDPQK0wgFOPnC8rV9V4+I36+Es3jmMtzqsGtE2dJr0Ixrha18E9lRP
YejWk6BuzWV0fKfqIq/GjH5A9esr+8fCKBsNgLsJMGZNgJE50vk76TkfhnxJL9bp
EcNDICWT1bndkFw8DcS9dWs/YA06tOjeyDuf/SwK8l4rvy0otfxPcAGdVpNK7q48
RUIPaVM1aJvNSpUg/QT1tTR7aiVlXXGlyRCwnCiR8tWJ8rgpB+kgqKixjK9kDPky
8D3PGTW2tAgWxapKKXK783cO3V1JZbxksTcF2jP7UjAhFMAVleST2mGD/9qvA/am
J2TP4NAxbWmj69k6knZecbUe6M7+zvFslZz0zL2ruaZErt0+oQnCMCZ5XAt5bxY4
tpuxb4POROOUy8VwvWRJp+t5MWCqLfjgq77fjrrLmC5HgqBwLMmiTDMoFiwKPfaO
qox0mnmVT2WAyd95XWb6XfS9S23ZL/Z3YYxa4CVVl5aakstGLFkD0xfx3eThf8UD
bjti9ZQk1YF4ZV6G0AxEPZBInBJLLkFsH3/KGz8z4gIZNpJNVJ1zS+esqI2/HmSV
TWO9PNxjbFsL/8R65im9oYcJRRilF37dAMBJBgmDMa7PvNzkNCkYKFfX8hxTVKQb
alfx/lfL7n4w96S3TPiOmEY9f+eyAZQ9WFA7hhu2MOEP750e2fZyO1DkVCtaE6RJ
uZAHmuantOb8ykXzUUkgV4hCOhqb4qr3H9XSSy8TgMon0ednG4cxoKqWgdgO38dq
2QimZWEBKgzWYkkyYwN26SUFU1Lulp93xmDMQ8Z6Bw5zSnbXC3Q9TTWom1s39FqX
Kcf2+/Zve0k9hfgDERG+avIseP4f4E2NGN74Bq3gZAKdC8TWwx+VY4GDR+sSl5UK
XS+QbM6LcNbOExGCC2ZwibXBMloAFZeHZS1F37OSAGdXDVZAgLz+nFe4AbQQUz8a
rRnWhsu3YImCLA1UvyQxpbC2ZcZb/ihvQbxlr4I0+koVnB1NzOqaub6C9d86yzQT
72m+066ux17YOGvHDGXLp1QhkT0j4hl8f6694qd42EDkMaWDl5QeYTWhsbCDSPpR
E7jy1b9zdJUdZUU32m2Y/zgpm9zU1OxGkCWMJhcExqtIEcPRgawXTRIPxPVK6LnA
xgTUCq9S20b4jQpLKnVHvIGX3UxY/3f+7/dQh8xEKvHhghFUUGYlrVqtaAKBxa4a
UTMNGKBPmMhZlLrdfZE4owhbcw5eH1IfjfM7MRKqh3+bW5yMTFckw6Ys+9U8b233
8oqfH1m5MRxN5WnZ8uRqQiGSvfRto2ZWSWcskoroxS2eBDZLcO1OClo157INJZzd
cvh1g35G7ztZCGxBOE4MjQvOGgz3Fyk4Uk+oChNOyUXdvUn0KZWQOu7Alf4S1Xug
XSpwPiRLZTA/gSJp9pU7hLCy4YEYkvynR5GWpoNrSkTu+laTwObF69u7+jJudSEi
VKF44vGOc0xPB3cc4Urj0TfDOJdS0FeVgbuyX38+INs7YTO0iopddT28p+yHrPSl
23xvJAM2G9wSkYYNADoInVH0f0FImUtfvoX/SnhuCUnCkfaFPh85Zwn6eaQrFGOz
PsFx3+oZWsiu8hIZj/f9tYcd6OhmN3r6oirtNjpLXN7cBXkHJZkJpxPl2Zz49l6T
snS838KpE9nl3yGHAcJ5ViQHNZdllyygnDgSE7/PToePxMYvfHmpI3f3u1deO208
vT/m+rcll1GRRaKkx5l4aLrVS7LsXW+pQtobxPnoqhzuXYb13an/dwhCTzVRb0N9
ZBYV+6QasxIthJZzDN1/yPhSOwwRbIq+lkSAQi4niC2tp4TSbPi4FGuczDlRm7Td
ezBMVR/SUV600aBc9+oRvUkaJRJGFb3ltIGCL4MIZpBziRBPJdkHfVQPAUjImYOI
dURaox+SKPogpw9fgtm+v0ygE1/gu8oxXVU+fvnN4OXLvrxSBVBSW7l0Q3PVOE/X
Q8Hsc8Fa2MYetcZZm7Y+/8KhpDJgRBEd7knl86a52V89Mzb7KYv/ofnqUl5ygof8
xWnG4yu4vAEcQWpc3wXcJM8rCX8JGpCRnCvXnDXvfCSo/YSA9h+v4+WbIAnml9hB
tUYnmWI/TUHMdUFRE2XExOqtPP6uwicUIKWu7JMWPU7os7QiFQaeYi9vsMqY63wo
RXc5jwdv5lGn3+0wFJCFexCSZgkDD82aNTVeYJbEd9+/xCFrABzGZ2u/Kd+OBBNW
okUg9Atrzr4lRWcR3ny/pmbWOaBFsQBiPNhgB7oPYwbHOIBocdZhgtaNmoAKNO5E
6+U2vsDzsmspdxrgSg/HzZFZkQ53XxkiQ4ak5orCPg9uzAe5AY+e0CWlFJa4yonU
5o9IYZAxWbX1WIF+x136xtRsEJcq6nxGUdTgdncEVCWAqmMo3LqaMTRM4xqWTtLJ
1CSbfATyM37yGKicNjjH2JHNvU5boB4Vp4h0C2RWPo3N4kP3jfadeN/ILYlx/YOv
4+oWBXAFSj2CHpb050qptoGT3vOttfup+vFqN/v1wmw/6+gk88mhz1Yk6YOxn5jo
uK5e+QvF/Dha/YUopehxF5Lil5rf2WDSlnVWQ3bItZv8e4CIPJQqYSQFG9ClkJLP
ccRXiYsIVbvBWbVusvJjARNwG7OsQfTKiYneTvp9A6Q9Ny7TPcqqy20ZKchkFmsD
nhC6HCl8fVMCOzq5/xxrTsPd/XoxML/IxtrzBJX6ky4u/24H5jhmVYSDBklskbgU
JmtTE235K/K3xyQANfi1czGxiKxTZh8zBLyEJgOgaoIQEfVW7Jbx90aRYqIPx6rq
7emKpaI4pV0hcD9VcpuWNh4pFx2T9ka/ZxCosO3ZIDvALzV5/f/zo/nZLvq1qCBo
YqLjEhOjRWoZh31Il7K86ZcxddzzvUwKCeEeaQkUA0nKMzDoNR7DfscvTcLr1EgT
6NqIHPFkfwYcXlKfkzYLYWNyehT1MBaRvR9qOtYhduIncBKnzkP1lP3V9DTiatsr
cIscdXweBHN15J9b30HyTFLCQQNo3niLSpxZb8FOjZ8h+BdqNoh0PxoKkuqLWaUJ
30ZER3lneJ0v9vgv2oXR/17AF+Yg7fQoD6cZMxVn3usUyE+BdcSJYTuHJF7ayF7H
mLzzcV4DabqDfaEbPY6j4tDLLUgyk1jaAR3nr2+/lYaJP9hNyckV7e6iA+q8fPJ/
UbTS9LZbZf/MyZh5e8+yX/fxCCpOPwkulyu2j5nkItoMcUl8QrU538y6sH8NW2HT
MDCtXfUbtPRw3afI3/ciXZ5YfBGtpCTgPqRlL+RXrh8FKKyo49r6vtSTDrV6YoMv
9hmcGROSLeD0r4lYodYb4XZ71w1pGlQDPRNG6IGcebFUeauFpQSoG6Fw4RqSI+//
noL1kF1gD3f0pD2z7qdB1fecxPqMgxkCKh5pUmP74UHN/HiDnhu+RmAHp9ekFXiH
5Lt/37G5aLoer8dC6yfYQJR3kMh6zW2e72D+NeHa/czc6K5nPX+MADPsLjUbs/vH
euM5d5kkMj9l8E4h9Qgy8QOtd93dUXDa/BgBAdg6ozXKO+2M50dRiABUx3x0bAbJ
/0QFtw7P3o4ob4FJpCwz4HIafPHZSFMn7dTMgb2Pf7C8JYZEIQEaXLxUsQAi9ME/
Fr2PN0/nDg0J6GHg9gEszt682MHdNbX7BM5AmEmL9dxikjk/6bwasI3LJkr9J9dP
vrnuVChpdwfY/bAjTKUmLLsP6QPbRlz+DImhjMNHUQnPh8JLVzI08/gdY4zf0+wN
itDuY9XJuKXUMprhQhR9jMe/DfPpQ40ZQl+wR+GeS3O2lxR+T3LceJzjEqCWK2ZD
s1uIfd207DcIjo8HwGH7wk1XCGhsQFe0pDm3FJihSWEfORUpkXsKxEMSKfEkzOPr
lfTuHSAto5Oo1RkjWmivFj5IpPhUqEBT2kdh+v8uXZGnIINYYy+wg/DPHFuzayL2
B/9DbtujSQ6k+xCc8OmCnPYY4V1tbjTk+9iQ/wp06Z0qo9YPaug4cEkk8YffokPU
sV4wqsCTttavfLeg9s8ulDP3XEu1juBynBPFzAPNL31LC6nBj8QqhqYi/KvKoDdf
I/66aRnVph/CvMmy1u38S1DHrNm4gvTCT0Vm4YmJtoBHbSUxCK9TPLZ+Yzo1+RqP
sqnn898kuPlrXZxRqMg1dgGVQ8hu7QkZZizUWydKOI5y0L1F8L11L/v86P+l7wOS
FDIGQfo/8DT/ZBW4koZGBbF/AkzLnmfbgPNXG/EWlLr98bAz62IJVWEQXmtZo9dm
9u/19GErL0t0x/dCcX028qx/2L7W/qpbPGG7UBm3RWH0aW+21tqxwa0Pdx/oUns5
8/qX/oeAajQMPU6PUtw5tkS2OMy3H+XA2A8QGPL4P2yEMVFeXTnSyUrqDbpl+QbO
GNo2trJeAB1s0/LSk+fmLBsjLEzT3o5V4l9FoScxcqL46mtC+FuW0eTkLfWMsx0f
3R06Rdm1FbS9aCDExgMTSrHj3KBJdE6FvdyLR7DOmKWeIYpTQIrjrCX739EpwKNb
0W+omRIzlC8iqk7+8jPNeJv3P1z6wmuzNYe9+1EeigBGkwgEiTYarhaOacsktlyg
8HOZEXfYoXfSQK3jyNpGf3pUiexg/Rbjkjj29ToA/M7E14CoQtksOK3RC9Mg5W+j
F+p9yrmAnW1co1nk3br4oAxl5zUxSEKglz9ocmEQn9OmRPh1tAbOr7lWYeC6i5yw
TCE5DQyPTITfTTkIh7c5lepAjoAMqPXCl3zsdOhuJBcoj/YFjpStpaUFQmJ88n+Y
WPVACBIncKD7J8/rDUaa1UzBw5C7uY7tZoL+hPO4jjMrbM0ZT2fTJWQ3sqxIkiVA
9FCpJ2JZdkr+qly3RiNdAYKFMuLpRkxC/WnfUrJm567qUJ6dWot/rf5iKj2W7DxC
s7vOugI6iIiw0VNvyXRzctC/FdN4ym2xZTbG4CPlLbtwFLRt1YAwfP5G4ZxrntZW
69ZssXS80bbpmcOHv9MrE9eVAdjhywopNllbo1O/uT+AEYiWIxzzy/QHjlnNaPN9
m7Fg/RDxoLtqqikgOjWr1Is0IQ82PQU63+r+8hqvu0ZyC8pMjq5/XjrB03b+BmOk
XVsxTs+xRicBmXv3Gh+7RmvMotBxpAZioNM5ZW2l+6B9R8jDgcg+eWD85UcTuahj
b8VQVZuCfbMwfXvm91hbwggRMyJLWpAJeabk/iVU8hhMp2OpqJr+z8LI5Til51mW
03rsxuP4EfG+wPWYB5FyjNRUSNdH4uQdGdHQL2h0sqt7urm0Q38TRAKbbS9hvKiO
2lP8MGt9mCDOJIKQULLIctcwU44TczoiIJRnZEBum45+Bjyl+3H+m1yVli01wC9R
mpFEt1pKMSVDRIk0j0ZY4vpFbXDvvWOuR5HycRCubenw1pfomxqlUx2ROdBu8Xzb
5EYDkjfn/fP6wJAqm1oPUgqrQsmLuMjbB1URinwYaFFBcN5rliT5q5dSN3gpPlcf
NAw+DsBrEMg9FLtqFotehPRoLaIyAOlBO7fIPi2bNxiRCok44dNShZzUEyDUEiNM
J7S/ijLaEfdKoUC6cUigTkgyOuIVQ8QzeCjTjbv7NivjTrVnUHFb/tsg5P9v7Jwp
P/+lxo9o4JHxAcqgr4efbhQTJZYNCcnOpWEk++Uben0vI+qlqhg1CxQkxNqYEbdx
hviORWSmRo/5eNa1x22rHcuICaZAU+CGk+KRPUUSW0NNn6mGG8pjP7OUAecRw2O3
kTblGcrclVfuKhXEW+D+8zip384i/7/zUDtJaCXtK+1f/3K/z9gRu9gL1xURs8dY
AxdZRuo/eT8SZKKkA5VTV9ZxDYc5z6IYaI1Gfc31tpyUyI/XRSIsfeDcQAPlGy6b
S4gdgKj7ImHbTMaXSRpiIlR9wPNJnu2PyGznqBKew5nYqqwKASS+tctmVs5Wls2c
e7DDfQvbFApugitU4ejn3bzwSSyJwvJ/j1cv6y7bdBjKLl/VonyKSp0yl5seC+7l
hpR6kvtEUS7VNaWj1ovrB+UHh76mRu/VTYyRajy6qxyjuC+AQ7+52ptkvNWzURd/
N8quYOlWx/FI74OJXapyyc0iD97UPYL3VOpv4fk2z0clEh+J5EPpRA0tVWeROznZ
lh7/pgRobo+/a6gl8QJW7Z/ReAkgnhdptDvxJz2uyjO+BrItNLD40bQq2tT5AfSq
+OZrvsq8WeCr6vSOw34y0ZxqOJI6UU1GuiHnA27Em2412VM5+b4p39C5xosSQeQP
SBEwvb8rUGlq2y59wAaQ1sb/QBon8QSkeFruRdUG428q3nyr8SnSgp7yVETBkd1Z
SDykX+nk5WAw7XP7xjTRCzQjnK+9Ul+x3D6CmP603pPKQUWvdQl933W7ilIASkSW
uHnFmymAYUuzgE1+xlLN4m0H+jOYiZFBDZL0gvl3JZbTSoEmS9nP/OVj/HU1gryk
ciyR3zhZwjq29sls8/KJq3jAhUdlVsMGDynZdj5oSGRueGlcYiXFIupGDD+lz2Yt
uTr/O3njkHsBob0MnNlJPCJIUMURIwuJQtooXZUfTHUrHEYlQagrtp0XPcQ3I8GH
a3aPX9KoGc6p/ihYsCHHyIU+xx8117+bZN0ntNaFiyVECFPk2GMVNaRlaZHDz2wF
Bd5D0cWAVsKO/BvIce/3nwDnCsPlutu2GOu/QiNHaWnHdQUxKElNgrokHR17YbZr
M2bzY+oiQTzwRnqC+7k3RIFynAaiq8H7IeMRoPZvqhgtT2Rq35iYFuYxbpcgUCkN
l5x0Il330P5IjcJP6N6ZqFGu3ZN6XGPLbR/3araChJb9uDQbqjWZDnnnifq8Xkzx
4MasknfBiVRtgiywPtLAAH6eiTSTX7JKNjVpq/+P4qlnJs+UUuw42W0WqGzHX+52
Hr0BNTVSbfBXjMDy1k7E5E1sqqBQDrgGX3tnKYgsb4zvWnBignXUR3MUjZ6xDJ+S
BtuBVfS/RWvrrP2WIdJB+Y0XtKWGg7/4JPojp8nRiEY5G0LNsX//hL9tbDoUofWG
tXdszP+70W+9Y6dx0wDSa1eCzykx6ZJqA9tJmTgyseVSFW1cp26o4LA9AAtaUCvI
cKkqP2tvyRPCUDAaLSI8as27uhzvFKof4EXhcCx0V9yT3bXgB04Opgb2Cpyvdt0b
bx61RMGkeDofTVF9ibiHC+ByE+8Dekz00N2ji1DjSpNTkDOcmiPWp2smXKM5vzqN
uipohbtON/5FOCLB9S8HEbVo3IumPb8oDZQunynLqXy8ekXUzNNn62fdqMVhgjr/
Gc3PKBUMm68Om1zcsiFpJ9qfECcz26AsonO0Y12bxUfue9sjXK7ccD917X6fE+Nx
jZJcOE4tznJXB2OFFy7sCN/mZQqLO6nqDVCvNUONiMWFzVq7Sc9CcB9XV/Weoa7m
CyHTehjpE5iHMv/n9rL2AlwBUbOWsRBUUsM9dxcn6MHPkXXXsXrOmZD7V6ib724x
4o18X3CC11P2ypQQOE0eWWiYCC+++tOcup4nzUlnRQh0Shb4ZhdMfFGmKEkzw9Er
Sb1VCjNuXxF7A3iMNw52gRHLf/NvgUG01aeVHD5Gz0yfWAogwegl6PZk/LxAW/r5
4WMfcEhM1pZ0mK6SANtGj9iWZBKkjosFmQpZpIDO5aarjmddjCHtNvK6L8Ef3jNG
mtHMyV8nXpwaeiZCgNYXGX1eW8GqEAU9vpAdiigpBiI6WOFplFbsdnIJA6LKtUVC
Mmr8ouV8YhtQ3fJ6ascqXdJlA0b9CeFP0gDxuwetRLPimDZBruor+MjNIXn4QGJJ
5R76AXbJjYcmJgHg1/51pgIW23nvTznvdYqyzlbisvPrInsAQtDl/UJwqAtxedbU
X9JySg7zgACXxVhzwjcXgiobcXRVJm2WN1by3UGRNsNEJzgybuf209FBCDUrDvzn
uhN0ejCEuj9BUVSM4YbRkKh+MD23R5HEUmBbYByX7IZRQDYhj8YdQhr0A4UAdfeZ
JPqckACd1m3/EpOSoZUjO60f7qjJh8jqZEQNHDjKJZivtqUnwsI7pZ6/RQTXf20C
fbf8QCZkJx1oS5FuZEYM4MRixeLrtnCdDW7Kf4llu6yqdmwUYRovW9m37AJtKaDB
1UYtVIbAy1XhKc1ornKXmYdzaJA0x+blYdW/kizeZH8aCoMlNP+vskONTRVLTJdK
mfKFrcmoY6ZvXq4SivgocRlA3XPRUaXLf49WwIM6YmSIP2F5k8hxH3HrPe9h8pD2
iyaOR2577BPO6bHCD/EvOtY5DaeYhrF50ZWA5f5S0GvCnQF+9W/p5IBWYsIQbYqz
6AOEdd3vCOOcy2G7VX+5IrPIuS1jXmxDYlQcxYLW8Ty+8S/XeNZ3o/+hpH6Elc/k
4j6LDv9qjkVJCRNzTYqahLp97jfLm210suK9bAZH5Cjt8Q0sUp+q33AUF8BObsAx
za0cTs8NqaDUlk+TD9ynJCvHftySP1DKzAQO3O0VcAfLThNsckRe2dJJ2xNav2qL
HpEEVYpv8mHqjRx7sk4+Y8VD/Zod3p4ubDEx2ZJ1vnPxkK3Tel/F8ZEjmRVnU9EA
z1e6uCHBC7griVO91oQpPY39w7ghL6LhdfjOeYPGGKiFT+HMHsbO0Uku0fSuzszA
Tk6FZauFrPBMslor8S3ohwY7WyOM7rqWYsS55Ls1VMjHwFkf5Og8LLkZyvNtOAf7
7fhr8WstjD4mHDnhb1jwieBD/U6cpx88mOGiobYZD48sBqihi6ESel5cwbWHOoGj
uCo0Y3sVwcRO968opcnzQ0lBcaqBQmtnJOE7uHkHD/qX/rHzWRrJBeB6KjD0chei
P3KQzRpubR4CGm8fG/mshwwwYPkEF0mwZa5/XePuRfk7GkQjXJ9urT3mcwgIGNCa
WemjPgeY5TXbolVtgoF3PJcrbcNtlI7Ug0vobbqqCtkvwaKmzhDIlckVy2zYP43o
cz9b1s9tcvSjF/YXoP+Agu6ywUYqop9ikErZspRJ9TyqlHRyoXDaRj4F5oojY3kA
ZY+h0SiczstKx0BJzTbsbOGEKV/52xLVGwSpYLsVgoHbLcFA0V5A/RfNhqgPV/JV
al+NYhs6FhHkUzdAbqTvHne1ByWfPvk8d2bwQQscpxbxVVrWh71Q+CaaHIMX34+V
xEue7dlPwbEL/kW+x5PgIrcqsTXnH4BeLHolO51vaxf+K8k+awq8790KuIbHkLIu
8ruMxEhhq4Bi+N91UPiWZvNURKO9HRm7Qp20QO0cTcO77KCJa0ez9iEzGFUjrDSr
ZYQOK3kvwo5aI8k9I1RfkfzaxUjhfn7n68MyltdpLtprRr0013DBdybrFPAk1oLZ
1t3tBA+aAdtQ/5eVhpNeGIwwhG8I70aArKl/vXK5vAaR9zcWPRY0NsVoWwl8189J
ehO/o4TsZQ/dV3n0FDOgBFatwpmalNst5xAkWazzaJkHj7e5Iw05+Qah9PqhQH0L
rCYCkJenN/uhOg6j6g5mf7HDU60QzJFMtq72sp3bo7tL0shvkVbO22++nSUEc9Sq
oDucX+0VTy2I83dIJkO/ts/P8pDdH9nBALHC5WaLe0anGrd9PY8FfqBN1Xzk4yut
w0HysO/6O1pnY03mCqdKufKjIJyYu6WTLMBoLaM3TieuO4khL+OANK+5FZtI488W
sQ0eQH0cdKwn/wAwMJn6P/jEoH5MzRFcJmZ866POHtBMvZwPQlHAGB8LYQLI84Lv
arh+ILWrj9Oe1nTIhVhCmO/W/V6/xMT2eBB5YMWS99z9sCn00lr0W2BpzIpI1LRj
2XDay+/KJSzPMTrh8D/NmwFKPAMiAYL5Jtnroq5vbr6uEUBwmIOj2gUtpRnj8qTn
IBiI2T1wmlpIOHkAf4ql3Gl7boqgNq3f48U2k1Kp9L2iXMjYeYa9QpMlQIjdiw6R
EqYW48expT+WXH2kuYXVK5xJ3rUz8ihbTLH4IOZNCPSjDs/b6Bg6srE+y4DpDy6l
LRARUSyNE3xkNxpp6vnxyBZaFuZNUPpJyM0k+z5gJMDZfVKsoF7gzDfG3LoaA+pn
XfhdY6E4fGwDtqK8jPcbr5PscXiCBWafw7vkeWy5D6hJuW3tPdgLz147pVuNETbo
XPHFVPs1Sy2GZri6c5lkQWzu5NRvGHLEATbi7jueyVCx/umV5F34gVEQCmkDtEI0
vuGa7jUEGTh4lijHEeSRaBNOfpDXEOIXnpEiT001gm1N8OugVPiZu/WRJLcrGj3y
rfYRuexMzxGhVXtrHmwWnK++AwyEv5+dmK3yPW9DrmVFjygK3p5F4quNshAH7MUQ
BHDE+Ht9ArZDMxlDPKc2uNPPtPaQMOyCjQgccgtL7j5T1U74ymE/TPMPtICW4Sz1
1wKCdtDhqPXoGpYgZyO2rrBbI68k7uyC82mG1Oeq3+dW9lTv8A1ypMcL0ZRTS08K
A7vggR8gSY67dMHZhyOk6JrifpfdtdsUCQWqntF5ZOrPqteJ5FM6e/4AvdQPIomL
RS7LbAcxvVLWnfnGhaJjolvtIMxiVScSlB6XUDhjwIISovZLcbWkqPrGj2dcRyMs
RZqi5J0GsVp/KHr/6BeoBjhbPrv4eL2ivjjFicWR0AuoVf+DLJJZFSKDeyAZMafx
unxRUUEdIy1slQQc47rXD/NNMpHYT+ph5/VmkvYb71c6XvYtKVeVydVC5/S12cxt
TqNGBq6peMZ5HPVvXSPXH2zeSE+XGM2urulWBnyQBrGl5Os/q+0W8aNvZ7OuSzL6
HZzo8q/BkyAXXP09UVVRaIzKsl9DWt2aZk/J/fzY5bc7ziXAoP5yrFRMxh2WvlM6
5EDkpMPVkOhlGkOoUerp0zdfn2APKXu0+gkkcXEo04OkbDc/UL000AchWvq4hTOX
dAVjdoxBlx9KErg556jzFxgK1Rt6Tqbts5fX4+7FPjR6pRLWf1lBYipU9dLTk7hz
472O8aaij7Kof+YdQZxXWXBOzST9ze2bddkueyrv4+xJZDHS+jt1dOXJty9bxcQp
4Qjo1r0E6zzwTk39fl1AAT6+bCDjhYRJOBXZbh0nKyII3BI35LCmbjxV1KuYcTvT
y2UnUGwNjcOxbn9tWaAQICr/1fK79QF/CP1Jb87avkJ7z/0qQzxMu82h76CAs1qc
2vMmZhQN6uSY5tznEOyJqDlKyBOYOnimBwJ0Z2/Fjy5YE7b36KMdCL8PTGV3jg5N
uEVOHBhnVKNRfik3/TzAcdrgTdBGm+WfePBmqvbd38D6GtXTZz25/8chKJNrAmj1
el2+6ySkfyK2hdqU8REUXhbhl9zAHy5w/TX300lqc8S2PvlNciS04lYh9GHaw46f
Kn7FVMjf60/EUaOjREleQ5Lz30WJdBZEGXgjdkfCCQlmYNsaKWct2pmwwB2HHiN5
5VNFiEkxlbXMgSucVspm7OUlDKOjNg/8edbHAeiVaqRKfhvaPdNMErqN2Q+A1VPE
6JMR+CHjW+vROenjA2NAvn8a1554Hp+qSkeEgqUOMsivIL3sMLpc2SIsInwqw106
RNMOw4GPKPJNXAwuzwkvPp9y4Sunj3wVXLp7W/6qEyT2dibDRmzULrubfGztvJi/
rLMZJ8eqtBEKZFvsFCodByPK+D0/rGeZ+USp5rS52yiQkjmo+Hip1I6WTaobUQmX
bCscFAiWGk1VTnwe+DzMFTVc7JYJ32otLlJEXV15JETvWWHMYG8UUM1nHGmbRRRt
0T0dP2iRDgzHOiHm00BzDMwQt5V5psWkLj8kfs/qaeUMtUAqqsZ6jsxxT9srzAxK
WH9iaoHeSNYCYRbLP3ZCb2PpL5Lb3QaOvSVO0qi467KCPSwayD0C/9TOWkTypxfz
Qaw4uHUtFVROG2fwg+AiUn9GIutuDQX4VKs8eB9XZyum9nik6JOmID9TCAiA9slo
DegAvhO4+Ai4zRXikelwhjclRxwoEAgjS8TqMJxi9MSNsZ3hFAHsXHLzp0oUOMWn
a2xLA0kzLtCVZ0QRKiIJqYtiEoa8RoyYwHoo1oR8OU4/PZukXJyVyHzR8kKsszbY
7fXhfXaZDnR/N0sxHrelTg==
`protect end_protected