`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRagKM/nMpyIo9jq+/KCuNCGT
x06bhTtDgl4AWxu9m9jPLAHIuyNRHe4Cn2D7jjDFd9yWnUnGDgYKuYNpjO1TjnLF
DBUWrElcOV90HfWVXKXoyHGYjibTdSk1R5me0KGQe92ns+cSsypwQPBbbfYTQ771
BrTGPDUUxTlO1TtAJXwvD1bwh1w/1LMo30DmapAwlYyctBbovkbMd8Rd8YrcxGr+
dmiYNahlgsn9f19IFewVrEDuUd7h6wisHINQjtNBPyEhwthBeLAphtYDPT65r4AP
u4Q1TU3TceUXLhHrXmG9dvJB/8nha4IlirLLmG3UsTA65wK5Ck/fB6JwwgTSjGFA
doMwMYyR+bMU/h8OHTT60oAN9ekZXr3yaKiQ0KK3YD1Lh6QH2W74IQtIzlvdyLal
/iZWBMjaKWpe1VjGgJazbzFdqGXi0YWNn6RZ59X5xfViMVvgzJEvsOS/jS5KxZIQ
rScR4K7vD5qeIE6ZCD1dbxOeLHyFWR2Ejx+BpHoyDMKzJtj6serTwVvLBz6q+iR1
oi8+Vw5n3PRNH/lCGJgoeW8iWiJ1E3fuLrn/T5Qvg55GzedvCeuGKlgOI8PVZ1C9
rglCS8Md+fvN3mILBaadoCYbU4Kq0VWuZKXJd4M/mK9hqmWrhhxN+LsyLJzyiCpm
CKbDLSSGrZNfXxD8F75denfR39sxrghYZg5UeGgXgi78E1eHT/Jf4cLDUovaxKEA
2LK9OQYt9NfL9nD9oG0t0TNNyblM+e2zjIPVUMEYb+XuzR5r9sdgzsztLXImnv0K
N4W6PbZmkvfEJDJ0Rl2m9JiHZjmrhxSMBiw4Xi63hEOO1xkf1bhmIxVmiSRauvH1
rRz4RA9ypIYmhKI3ZLmpkD66ULnF64IB1N3MFdLQ1TubR9Yd2EeNSjsDxAB9uZn2
68k4ayQkhe+IqlR8FX6bgDKWo0QS+YpOv8DumkpRQ8F+hcVS4SDhsZUJL2WgYXlh
uv/Lyx7fksVbIWKb9l4YNSA3+XrINDe/dCdCBtRIwWGZo5lr7n5gQeLP8eBcoiSE
gLPz5iq10WSig1UC5cblHbOY2ndDJPtw0GZvRvdD3GKsCoQpilK1h947RYM9cgGT
4bJsmS/qyQ3EI3YPVrNVI0fGRAIIZK/Gt7PWpmM0xILy2fd9uCkpJbvOYENkKENw
rKAFNsxNEwQ+VB8hNfdqQff8l2jt18o9FjVrgQv40ddjqBUrP/e1fMZKxBKMjUdL
5KuvvhqgB2GJZ7YiJvOb1WG8CZoYcwpbFzdZOGAQ/SkeqBja+erMXNDL/6vH5dEp
gWV31Iz2KHkogdKgOJff9y7fet53sZCkh9bvrNulGfip2bR66VDueFQGXGwGiWlS
bgWZwrLPIPeXfSwX+us4+jGLq8ctJbkoAySGepN6E9UW5xMgq91KNvmX/5c+2UoB
bGF6qLR7rFuhOkYKvrCoDtWJr7RhB/2HMH95rfgeeOB6kqU0N5IISE0hphtNHCDx
gOa41T4QlFeuTqnaO6jZ3xCfMgcetkbuiJ5rJ7VLWZi3mjqO+7GuvXP8J3xicY4U
9j5KdlpotLWyBYkWVqBdLpxDTvNFUQ9mMU2MAWs/NCOVkwzq/LHdqBxC13Mh6rR8
Hj0USurRDloKcBNeWnAgnEBTqhP+CbHGDQsq1HonU12jjK0VxLWzHMNKP87/Jdib
xdYkV45rYfaZcVDRjjveTJFYY/IaLatO5vv2fHItCUg7HFW54E9lPxhSj4EtOazZ
1GxpRDmy1ABlcK5KNKmLJf5uLmcEsWWULpDgcsQ1yvjcFy8q/pXu/GK6vQGSFDvX
ylwdwEXTt/BTq5MlAqnfOVss+xRTvq3JYWOV94C7rvwvzcZjjkKiJbl4kccfAU51
27Bfle0ExLa5neQo+AquoDfX5qXt0tbkokwtXC+ODXEwrxt+h0pWWDOeHnmpnegp
RLZRgGjww5INDMVWoHxP8HT6DwYQi1LAC1oYZsbarO5dnN4sjHiEjtpfl4Z6CDPA
ntDVoHdRVryuswbDOUyM53J85cIKJHCM+oCblzzbOQo9Uaxo4TR7jncWh5Npjbf8
Kmku4jIs04so4FArwlbWKgiGIAVwx1NMEALSpb8qjvx2G85QntDA4QWDUV6rYM5s
OBqqAvitncL4kbvBDcKPGc55SDQtKB5JMlqZdhJTl2rZ1HraOzRzGSx6aHdo+T0n
jgZotUYVRJXBNjan79yl99xWADvHh8vLjpbHIMG6YSOhPPox50t7KQDsFxNGI2Qq
KEbTQrs3n7ijZWk9w7RG/UjqbOam2f+sRq/k9gNg3ulE7szwtd1EUxLvoJkDRxzB
H7E9T/843lC+58ndzn5esWAqABXO0VqVQhfzAGqgErqNf6zqOeSevQigaJMo+Nfp
lT97Bx8XOlxfVOa4FoZNIgbRQngnfHgX4bY2BwvzLlpBDffBL4EXud+HMUgaY9ML
5ivapcYUice7HaeaanC9FCHgxmUBv0mGW56xJsLCYPTd+nnYe5EDXSQ2IQlt9q8h
47cFTJwzeGVusqOVW/+PoLNrB19gweLRpoUcJmVZi7GTjZ7n/WCIb1DCWasU+syc
rgxN6wXxbK40amxP+bnE6sb+A7Mo8h03le6/xfzcxka27FOibcXGZ5zeu0+sFhsK
xPKZmMJE928M0y5pi44ye9nQ3UZP7eJn/wVweg37dOnNKU/BZ8aGJBqyGvt4nzeL
DpWRl2LLsKVchwiuTcSatFDEcuziHyMfJ/bOsEbofbyONldMKqXZ7rEgf6/bUZ+R
F8DidykQwQiPOa7D1lvVMXH8h4uSlsjHWfW69euu8ZzwxAof9hIJ6eTMYfnG0zer
vv+i8c5qKOiQmiwnAcxXa2A6liY3BRr1ok4oLEVBgMAjImWN6XN3kfHBzQt/WLus
lNC5lU+nSPHEvRxMaE8Q4DXLnuHn20rqH7n49Wl9c4nstvsEcF9L6y7/OfIVk8Fb
Tl3UGpwv2JMtuuZQXnCwRVZ0hOfK1tqKW6BpTapeuC2TASIvqFxoFATZArkWXoDl
OBa++ORH4uHCi7hiqHe3efkrZzRW3M9HJB7MAi49owWPsIXL6J6YAgWCFRS0cN8L
pLsavzc+zmyyFsv4rm4EZ8n4WIyImKigjUbpF7AvZ1/GuoxTZGpTl7wmjoGP+pf3
dsnYRLPgBIda6/Jrfhv7DowPUqUmZYCoZP2IA1oPdeXagMoMjdX9BrI5esX0Wi7f
miFa4f3a/9NWrSXpKu80xauGAW4F7UwX5w+PlL/09YkGMcIxEgesMO6ubJeMsu5D
uNR+floH86c4R8LQSzxnwmrJ85DN9NUULb8OLKMxCemhAw/FYpwezniP51X6XkOn
8BeAqr1YzY/nLFBKgyV7ZG82zzdopEpBtwZsDNef6OPpDTQZEwjkk20aWRCSSdYE
zZ6PjKUSQVZqjaF763lHA6it0y99dWapSsa12ySnOkmHF7xawT8HSiiYA/QgAnRh
JDx2OWVCjREYvt1WrPkL1HaIkfB1Ge3hiq0EFh0EeBMV/UJ7O+FuMl0VKy5zIRVY
g1Q+2hGf4H0CxnvzJtgHvMwB9M5ve0kYlwuJCvnsS2W8oVZk0KzmCd6QNeDs7jGl
LD4SXYdYqyR/dB6x+p6l+T4o1TctXtNGGW1FXNLly2gydj2AnaZgK7cv/yODU0Es
Dh/3QgdypPnx0gA6b/2Tcy9PU2YxPkM9Y+x9F0dvSNRL6UQ4uXdfZA+FAjY8Nf+r
2XY5+zWqFMffLjctDHltnaf/h1egP8Uvl6CEKEiR/9zP78jkeXjegc0D4ZiV6CKf
Xhe4uAWLh1R4BgAvWizPzDBu+cfuJAWxgOR+BhDx+TH8XAHsPJCku8bH7F5yZCLQ
lIDMyDzE19s3AzvkQldLz/7bxzvOna8zvk1PynAn08KTfTKfRybE6glL4PWe5Vb7
+InllOBnLipoEA5IBnMpayH3QjZgogc/q4F67JUok12eK+CBPH10In/x1DVsILam
P2fmayzYH4DJHQ0QGnCSF8Eo6ElKfYgXkpVXac4GyMiJfsZztzOvd3OHAqltmY6s
0nb0JPzNWxlD3I2snroukkljWw88L+kcmlbydwRQpWofyxJwetxQwTFqyCROQigh
puI7oiJYEplcrWBIPVScx92L7qkpk+1nIhS6HLS1DZ9/Q/0t4xqUadUqLvOinMAB
q56dmccln0VS/jwYVg+1U+x+nst8f7i/I12lNaBIxVX+XB791REb+PsJDXpgRbgS
9I0fduNs/CYu2kShOxkDMgL8b06taA30SnNSIJezIPkufCR4X/q87g2IrD8bDALI
APi/bmCnBnU3oPA07Wkk+HG4GmeSvA9NI4QI9/nAYwDgyum+tbJb2T+Th3x6Z0jf
hR3MdSTsygWrFgqVIPnlAsJt5qNHqGUiblRus2i+KpkZ9i5mrZS6z4JF4+QRWtP9
wV2fsZvgFLJsDqb+goECTzmpz4jhpGEMo6IpnoetlCLsEalmNKoF0GF4ZmvYjJhg
dq45+Xu0nWCWFy3sCK8ZAEZFtLuFA6SVzWpbdMipDkSMM2Mxqd7ZhQ0Bhud/DYSp
7IQWYR1rKQhLjohfnbhxQP5w2qm7qpCZoiMPaOo596ClHC9/+z+7v/N0wZ8VZFAO
m1N4eiu5NXZQMx2yooAUnAOPzhFdZT2L9IFWgf3WOPLO/fYAPP/lmZTFh2V0rVKx
cPR/MKY81ITJXchd23RBlXQEjJvWLdCQckcGi/2NjpjQ6r4pepACm2x3LLO/jGsg
Rs64Q/p8vBCsRLJmGOuM0b8Oq0txlTnfOorhqdjhlTUNpCSp6Iai7jLVIP1mQqJS
/2F9QQKNtWwH4n6TBlAKy+D/QV2gjZLYbDwIsX9hI23npifyFlQvV5+js8KjrZXP
iwN6kwQRWviRS/F9CFFSTOltcdp+H+26+EAmOoWgw97WBj0Dlo02AN8bnEs6tKUf
Si9jWpxn02MSFAozpRpzVRefUB2FY2iL2usshKo2nW9JUjoprgqzyrmPY/qWP/Uk
L1lPStiP9X6pBtPTLmTtbHLfk4QFvb8sa6hqJOnUu2E5KdYTyskU62Oruu8MOGXp
kwK0VBUfvJ5tp4NDh61q+e3l7MI1UhRXlw6liNOLXdWeWbW0vzqdJVf+w5n17yi4
tTsD7Al8SA3LSqeqbOmKdAp+jIFWWbLEWhh/4cRs6kfhogmi3JZGLSPRM3XXpMVM
Je2NKnPEyKybBeVlAdjK0PF2gSfyFeUjyYcuXQ5+tcdktQiJ4N/IilVJRL/55oWX
fBExyiIPexHNNVrfNIUznS4G8dLe/m+zgIg6e0Sjtl1sEPTUYlavz5KXy+nqkmQa
5p/AlbkGcI4izbrzk54tC3VGS1qunohPk8EbtN2I0j1IHnJLcCFb+m7ZON23chpy
flod+1Pf+zHYORnhTDIY9uDF78APgdmhBma0TXlM7qHX2Q2S9MiodMURidxE4FZj
G8+kbhMbgNMlTUyJHpthr+kHk/0Mc8KItA5Hy5L9ja6JdVvvgSXHwy3VIaGHI3A6
RCgo40pEhmzgYLYPDVT5PvrFkUYphCLPt2sMo03PLnXPHR9CddlnlSbKAJ+RuQsP
RXQlvU/s+iI3x2viO8UNQPC1JW7M+S+8Hc6Pt5Nxscr6mw0v0pAbuBGzAq0IY6pw
LxedBxwiZTpS/UtQFbZHBq2nlS8nTRpcNkpGUUVo1YoVu55IBMIWd7pn6uDhcxoO
heDPTDYsQaez+rixvhtXgAM6Us0zHV8Ttjpb+v5Q12WEjrUCNGc9QhUIvnrhnXeN
YOIwG6jc91jRWb21aSudl6bjh18hk+nQYDndw1guCWkPeb/LdVvz/A9u1AMcSNt9
DnL6q1aBT2o3XyUwR5/QQFIPlQ3yeSaXOAHDd8Hlu8Jr+EUChvZBGZuBYUqP2ESh
m6xq842VctXap2Ug8/DSCMcyjRwf3yPF8kc5/6SI3Cw0ykn7RvwgQYbRVh9hCgTa
643WGvsgHdYFaI9ykCPH4yf+QW5+4aB5yhEVMP+ytTvxlb/RFwD2fDC4sr0JxAGf
YwNga08F25SZBUWbeE0WO6kkWiRlfnwpesv7nfvRNxy4gAtCi1bjOH9qxTY7oKET
eilUgzT9YALlSFL0z+GoAP+DOgJbEp5+8l0gyjONpQ1ou9vreeXltUm7ZRB6u4yO
o6R15XOVkoTkNi9jDfc/zaMHbaURsmGhVoRiEh9YcFCJwHc9vOidOxWsqnIO2Do9
xaoMvkVzJMw1Bjw64+/klA==
`protect end_protected