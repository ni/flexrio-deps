`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
lhpPFePStMLIsTdmvDdSWaVfQcn/5tuBN+1RufesQw6JSdQKVXcL1InKu+/77hKY
BnZvTXDrjmE0Sfg+QOSCHZFBxygNgVddOYWRfcAdWdsJ4UmZw+g0+D1jWh29yVZ4
FKmLQkCdLzrmG71bsAfMmDqkIgsXnvuKHp63jX/NMm7Z//sOw9IQdva9zgRd/hXY
xTNXHn8XzOOvsIqMBxAXqD7CuZJy+pIu/xIYaihmPxSRGfXFKLq2bRbWn93Lr1QQ
IYfNz8ofWWa3CFzNbLTOtcIr7gRAvQ/ci+eT9XE/lYNSvjGp2+gSdytG56YhB3OJ
E2myEo7ttRouFq0DK7ln0RPtmraZ2GGF6mKj2l/zu+LcVMIJ7jSdpNVMeef0NdAo
Ou0vSp0CC7qBABsVPnBAa8p2G5MArbRIDf/og1Y4dFWbVTxpr2W7gDyvSnRGOQwN
bp3q1fVFunnFf7y1SrVApofDJJobQ/VC5CY3R0yVtn3yaL4SqtY5d50bu9s+2Dzy
cGn/0mXxnSVBqrjo6tTC03n8oMyrwBsHWra+GyxBPZXxhtx/uwHNIZgR43X3C2wV
OGKvqwNAbI8mJWhHRHYyn7JBfsicKWjsSrv1i8DtRdZJ3wVcUhpv5Jnf1wm56+oN
Rhi4okxOvHQH64BJNGmpEQr5Ft45mo/XW4YYa8TmhjQq1Q1r8pbeu0oqMul3MiSi
Jf5YIaMir/QHoDff9UKuxirCNCZSIhm4WDyC5Jq6GEi2Id0oEwbosErdoReZaJWK
sAxuL72Xa1DRlZ+TZnw/Hhl84elCh2zzeK+sbfaCmfX1sliR+CbfXCAH4Zv9j+b7
S8+59drpCc2EmO0ca35jw2HGvo5CKG0pH+VXyYaJuA7pGjbdv6mI4cGg+tVlRCQy
8nlL1tVcTS6bye84Jm2V+W5Cwk4auosVk1RUN3ooQtrBj8CktvrxE+AGpZO5515q
nHFN2qFW2y1Pz0QdkN+jfk6nx1Fen/pl2UMUNsxr93J1I0Na8ZBLpWiOVKYlvypz
w8s6xkoQvA2oBJoNuU0ADWf8qjT4gXNQQDUHllTX5+9zH0hs7olyZA2kA/ZORzAs
wnKYqMq11y7NXTrvTI0E7s7qrqiDiehnJqxdYaCkZumAi3k4f6VXp4q5VPTBdhud
ne4ZNx34WZ9bqyBx5+ids62k0ZxBBvwlEE0fksYqJRUarU+ldk8pb5RZTBJM3ONF
mB1CNcw6f/2DBJjcY+xWCNtX5Jrm/ZEnVgmdPhyGOOZ3+CbrQi0xxcCCXExRorJR
s2r0aCL9ZcRjWdEBuiR2O/D3diq/4EchB246v0uQzJkHbV5j+faGpbK6rpRMF2hy
0zIJoPmIa6055wZakocxPdrstVqzCjutkpfZR7Otm3rPn0LMfAto7v+A4uBW1ALg
4QbRdENT0s71o1Aqpz+uWJEncrZHjJ7fdD3PRuchzd/hehPnkyVVRk/y+nNt3JXn
+0BQR8RV5VLvO9dzJwPeZtEBUkHiScpLqlWErV0vzqa+AQOMvYukFnmkhsOHmBq8
gV7GJDW/1Qw2iDfXWsNCULy64Smk2e0jB+KrHvcIAuzrYvaKMcEjuwTgv/9QxDeC
uDIwfVbGUpOYOxaLtOkWzWIiGCrFoJcex2qJhw3SAAGA3eFy1H212aXso+K+Xay+
J9XTHlYkiDGl1IK8ouzbWN82GFhkvxs+XEICJ+CMDW0swgcKe+44ozfZAtttsk4d
vIedPJLxfos2ikeRT80odtAn1x9MSPLN+O8wlS+mrXmdPrxnhn45wdx+xXtwoTkP
CAVX4kdUcUYxLmSHMyhaIumeiEqbkAIKr/CCrJ/KNeXyhqhVhdoFAoyn4QCZsZ8c
Ta89/oNU/+mtl0Tw1TdwwXI1W8SPcKPAUFLh1vyqKN1jnThNCuDqbEVlkTxlGNiS
LlAiyqWeKaqjzhEohmClhxCiA9e8Z65Yf7Jtw6fyRMVMYEv5QTuJL4IxqehvYwgJ
jCyQQMKB5DjaXeeOmnVkLpPqWpMRju/4OWIzNHY8Yk2JKxmp86vieF+cYbPu1J49
NJG+BxCRb1+KXn5TXP0MKKduml+ByB34Z3V45FOiqm2gl8vJtfCxf3R+uIKO9HOe
Cw4Ov6iC5t0VRvW5ufyeUWtDRInHshj7EgabMHu0EiEy1/zvG9It41auFe0wtziN
OXQscLRfE8soSnWxzzZzOjdYzuXNxu/QqnOSVPHKdWZh1nHCFX42xjwEAsYdURP4
pxchMB/e20PFKD/iEXJJBsFrHEdkoAOoxwjRvDZ28QrKr/bXN1fEGt244fk3H43/
xCCM8Fl8DnN6QEnTWwzCAyb10DbM1R9fjlG/ncXFGxe2NeO3xhwXWImsmKAGdghS
yIWeGcSYMc5VrHoQyOJ+C7PcPyQUz1X3zCJd+1/lIkFoNsgMahmLIEMMQbIZatYD
AwVWLyRKGpcdVVQkoRQDlANfUjCuYKZJsAyOVGGWg3i5Fd89mNvVaYyeVm4/c+Ch
P5xPdmEM6xyfSEHMJ0HxhjYkW74ceYOKa75s4JMgKT7e+nWl+bR4BwXaQgzg2Em1
IhnaeSpja3bGT9YIYxwjQhKNHn2sYzOilNUjeoMqPyWJCCfxn1MUxkzZvP6RO/uJ
bng9zQ49iBZwfhfLek7jJ1nkM9lwIaxzVm1JHkdRDZXMhnofpIpg67SsByBAQTDi
9W+Ko1PocVdP9PVoGMQnWZXesR0nokRya/DwJ6iQhRGtPMMDws2bLzJN3YY0cjw8
ePay0epW/X8I11m9CzTYqX22voWF34f+hBk00wNF48Gj7ZxnJSQ6weM5Iwv4E7gu
3+yK+7ecQbmZjVYnHqWbwV/au7kg2LiDR14RSch+imn5Uc6cLALLBNi9PyTwSIOP
vweIylBS30a6XyWKXxJy+UVA+u+vU5YQIjKwvvZJoOsgcfNh5PXg5rKqbDbw/QQU
YCZS+Ry2zbcyQUJz0D3WSWvrxWOyk0eAHjqC1lWDt/b/4EBGlFy+Qly3qwCPUN0J
JTzV/4w4plmHT9oBZRjvdv6hUhiJ4Amtzq7WBCQ9Zs36nNsVR/oKm59kX5t39CtH
vDq1U+6qFvdxL38mK7spzpG61VL0h4ZFPoHC6Yfj3QNqU+ptQoXVykZfLJj1agWN
OCBde+cbJKvWRIw72LFt25eI6HsmdIbPn4alWNNZcDXWB5+6DVm6U8sDZUHNrx8Y
dZwirm/dIaClPduxyMzMmxhOT4ADk+HnyHqQCfUyVxVmCIAOfVHNR8GNU8bCZI5m
Nh4k+U0GVrjn8rsMC2yuOOnIASElMI4xnOufdJWBhSN8Nxcr74iryvZOOm/y/RmU
ikWlWY6ukohDshAQMiHB0KtDD5O0U37nna0UgtUDvFfbZQCqWPe94vvahZV1nR6P
EGbG3FO1YLUBB77jq/7wYHW+Z3zmlss7ZkKZnhw6Rox0cmYGlXAwjxrDvntnfZXN
PA9PfvqXHkX+OtTQilGqiN5f3F8Bt3kqCJY9naeSzEGtCamvIENxC5oDqccCDrN0
FuX31OeO91oXuDbfjldWdFTgw/Ml+OG4Z3q2+ZOa2GYEy5Q1CdYO8mzjOQaDDYcX
T0naHZsVv4oIqXXgcvOdGYmw/q7G3TGXEXoB8kx8C1AJUsynfNplPSb7lXVGB0zR
jQhQGsRZnLclyijl+aZgIoYHtwYbPjvOyRXwILOhjMRzybJ/09mfOXCQUvPUZwkd
xjIkRcXEDMo0DYKHxJRY6frwz1Sjxv6mzSwz7RUljNHrtFsYhYy6UOLlwAkwTIb2
xpXkOXDt0sGqv3nCWRmCMFIZmm3kE2Sw5oQogM4D6JHiczOsdHOvRU20XhHUeA8B
T5xYbsOn6y49ZFGqhWlNEcgkhEehdVgJ+iY63xOl5lYohl6IHdBbYcBXgv/Wbruj
pqMBjMZ2XymZgnHd9+gzMiRNjRbEFLL8clJOQBCxCiTZow6enLvtgGOnl3mGbd3j
gDy0w4pSwHEN2VSpGNmyHwrdIi6RNPhIA5btME3Xw05XxLWJSBdzBYFJXXvYyYma
a1Ojs+0xdWhJSFkDzXcHl6X6t2qNumQH9KwhojaWiDipmUdQf6GFyZD6MihRblGT
DQh5LYC4+fYKPhqicUtB1/pkT7DUEjXjBpOTnDo4Y5W9ow+tQu8aLFE8McCX2agU
OBA6GWMAxmpgTbzi/Ss1TnqclMLqd0ze45VBfwAT4f9dUEhb3plQs82AxySeYUKD
00rVfO0r3J/DxPBSLPjY2TapsgQLaRAoI/QLxXd5kFKgrsJJzyY2HMeqCl5vIPtb
WWnHN7gsJHmJPrQnvmCB+2lOibzvLM7UF54a97VgG84NaWKeOqNnGacfLFokk89S
12rS07UMMFGSGF/XKPl93HlC3gSRqgsys7rcvCGVD6ojvDwcIdoh2Km/mw3vVg7B
EGyRT95XakUbR9xVNv7iIstu6PksrmcZ6NtjLA4WUqpXGcjLmedL1QE5nbxzcuI9
vfXz3pvcSnJ4r1SG/vFgoE/BGJNHc5WLfTjHH9wtVDE2ftrVSY/WLjANmv1/Oz7I
gJK6yuF/MM0AzCQ9h2QMZsw0fvIWYFOknE+VvJ0VjkN6XJHahBsIbMVIl7eM+uQj
xmMeV6gCNzXExcmali3Uc0nn+1IG3MiglkwrLsLHXFC30SMLkQB/Q7QZz+Kqljdd
2hq8P+M4bCdljdXplpfM+lODjlxxxSbR9VdF1i2nS8quQgCTAwedibhJS5Q7Z2eK
Q99FI17OWOx8WAL+qJ2F/EExBch/adBrjrQO11JbIls+XXXNWxX8FugKcusx+oHs
K6mhhAzOefu9TCXVNV408gibmZMbGCWEfYmI1i0ujPlBW/3GLhln4SMEE9lIsWO2
mb7hvCtVHp05Irt1kzVgJH/ADf6D9HZFRSWlbw3YBro/zfdQQiF3TXZdqIpKCZqa
2OTcNcuC+sGGC9rNpqGftzXgKIzUwjb5KJsU8wwngKXgbkC93Sl1uYexQzkue2SA
zy7wCdAsu9jxcUQ19SgFA3hPUvj3zSvy3Hs0RsSGE8FMakpM50lTJXkBUYowZ8sc
aNjJQGTUXrDy3p3P9ZPlGVL508FSA4MJp3zLNtS0QOkjBx4dAByKwqcsklmdzhsQ
mvlUW+KK6ItmgYo/FBK9YjOa3a7eSvQZfVz5DreRcX9yvtWh1qsvOdBbTzAbSAxj
H0sBETH4uURwq83P7FwVoG+IMoo23+75Y84DgdRpxGOCyMvhCHhPe9GrLhP7skI9
IzEGht6g6QwIQVofR9WYaIJJzGahPqENH4b4035kf6OZbIHAx9hAq6UoYiQeKH0i
h3/mu7wr1zfQayPZmU7p7XaTuE0nck7XxXnNQStu9IaO2JkfVPQTk/4BMr1i2sB3
BqfvT3u9M98Jv9ni+seMAGa6bXv2ccQskvzzicjEKCTvoqMGyb/dp6dVEPs4N+nI
mcPGPz3n0ZLDV4Yapislp474FwLUOdsaAMqubSTzDtIgZPdpusKiUTIFmkFx7prm
EhLEqIisBGBjRPG8W9lgbTpxRsQ5ST5RRueivQX0qy7KXfH7k2N5IPo9QibyV4gx
3U0tKecT6mmWSSHZzeqGlD0JmwXt9+YqENKRvN88vOnoeEnpknvQ17dZe9KbIrbj
J9UN4d2aO0IAJg++yuoBzNfSaR7j0pFBJnvmJ8s6cPJu7yaYzPpHDPGi4Mm9/LHC
Dzbia4Wh7h2o6plyI4Xd/VSMyyYVwG7FL1avgosNHTXkHRDIU7uiTa+PbVKcC4xl
j83V2hEvwgFbsIxTGTV7dx0h2PQfZmnvezueGrZ8LDiV2eJQaI96wyHmxRlu/UKS
NHYm9ifYhim/r4KR2CkK7AHVa+5Op3F5+l1AkATjz6egLD35D+zPCfLPxoBN9Wju
vbVlVmxtQxX5IePDrj5rVp+tyg9evG/WuUip+vfWRCV1D6SCTZQ/qI5lgkNAd2jl
W3kQFuRtIDMCcXMUvfafG3uTlQLCQBW4S5Wov5fCgh4F5E7jhTphRxTLHs9xtmja
n0gojAqzFXGWabXWZaXVAQHhBUdITXOWJEe2M61VzAao1mup0TjGgVKe/hrSYBLF
LNUe+BNkOp4akkmu8aAmKfgewMuq8/B3ynGfP5cYSYwTmi2kHqyURlnJSMhTNhBJ
JHpwbSsgPCGqsQCzAFKSg4B4/lV/3VYOs87RmsWfnXtZn+RuAouQXnAPtQEBPbaM
iMFh520I4QVDiIhYj2JHNAb1e2T/P3Q90rUoKX8Gh8qdQz3DH9vYOSrVwSpjjtsG
kbsG0X7KJ63XZx2/XbNAi5fD5+QShKrUcjVnFM/KwOHkHMX+5mOQHuOp3YXBVI+2
kcPbz7UkSGL6BPRj9NPiVOGgnTDpY55/4EG3oPsl9rWnWvRTlIs5KEVrtAA3XCot
/lH7cK5o5qwmAXkYQMpXoD+PJsxtE9zd6eB+0t75y29bgY+OWl6C4/ZvR6XpOpW4
Oi2VHRGK9HtE3+ux/pZm1/CpI8/0BAsMRyBkZnEum+6yAThSw5akR5Reepyi3J4y
+I6m5QXezo9yGjKoG1cHq7c4tu4+NH69eahXZJbznadbfUwTHusNQWyx4YdSVJ6N
eoiBJuQQRyXLsMMWMvfUQn9fzsQ2sQQicYiP6oAb+Dl96vXvy5y24wKxPe+AmTrx
Mdf2IG8GfRcBOuADx12H8AWorL60WmKk6fjF5ZXmqeF9gNL3L8vHDnnE5/XyPyo9
N6qKjYJjWMYgBusgn1CymB5fiOhaAD85yF/94qyzz08MNn05V54aAr2w9kPCtxZ9
2XqJFT7ow8sWYyIuD4069txynW2GQwt4hHsKtJ5clw/udKLH1Zu/IKdRyVv+oLcM
Ol2uQWPA5l5R6CKSeF9zTrZMy2IYY/gQ52268+Pa7A2X1bsTb25DCI5B9z5nfJMr
0Q5e91d7oJMZKF85sEQIA4ksUnmGMOoudxrW9oQRU7EIRQv/a3WDezBspTHvLVu1
/gYPMHkIZfCfvK2laKfWszqrQN6jQ4IOdHYB2Vw0Vaum33Gn/D+yk8W7NdPG6aP1
kAQV5SptdtTvi1qnT9RFpiV74QyWBNDSy0KHJRTsmoh2qYUvfqayIUPLyvX9qV65
P+S3ejy914mBnOfihGAMlY4rOp4iEjuyKB9GlvhVbZUxNXSxS7d7ck9qIsE73bXf
hGr0jRWGVcn41xkDz0Bab+Xc/rVr1oM09fU5duAMeVF7TbXDQHrA+LDRI3uVlFcq
IBoibOVtPsfF+y09Nw8SEE319zi2tiHQTQKiycr4Dg4pKCpeQ0lOuzFAWrKW4fvc
0uADedig4SQqi8V1gFoiVtvUgjCXyC28YpSpzqIg99IQxLHSyo1MSRlR9L3a1sRe
eo6/79lZ4OeQqJrbpaSMF6waDiRam4usNLq90iNQnqUvJBWqsd5UfVSeK+SBt3ac
+ns+34V+98cRxRL4tvHLJnUqK9mDzHHrl2Bgg8ztBXngn5ZfDKheUAHOqOoSBvIO
3enyR7YA0YO62wWG8gdRSado7YZ4PkBJrFvaPdPDTJ/dAzc/JzxG1X32kx88umEG
Gc8vvBMWgTFnqzIIGNA08Lyr0dnwQH3Gv1Bm9pPOTpLO3KAyUmtWJQqUvU1s8SU8
+LEqs3xoh7hthIz9yFunOodOVlwAZInQwF5TZD/vLhjti3W/cEvZjXVfCKjoE+Ov
aS6xadc+8AOkqJCeKMqTPbd6+iVXBA/096130Kfc99DoY9K/ETCZVpWUOTia/82e
JnEvtjJeRR8Y86jvvpRV9Hf7XzqYAULRqkymzrhCdPjmQfPS5z/+GvS5mj+8pL/j
TD0zvSx2xpWrQisphwJPH4OGViKZbwiFuXn3074NX5mRJ0YADfBrm8FGfb0jk5VZ
qqMz473uAIXQ5tpApLdv4FpL53bl1sgmlYAf+6wbxZ17qtLyl3+RrCM6+kClQN5l
`protect end_protected