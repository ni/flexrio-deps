`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325sjWpFWZVqfqawtQjhOV9Ti
xjsylaiqHnTulnIowKyUkoyU6J/E3BHocHBw1HLmpZELKO/XkVV5+qC/Okl0Nt6p
sL55m5vHl5G8JtbNpJDh8GdyLods05RwSew7j8ZFq64fppRjMO3gR7FsxFi6hnn/
I/mFXhYsAl1s9wogsqF1aYh/k5NnqL9W/WGqhPwr/uxfwmJhTX4jOrVP5skEQ27N
HaDmAKO/FZzaXVTFwXxWiOxBvdYGyXtJgWs+PK8adaiu2vV3bmWQJ3Psz+p1Y51/
fLLqkTWISKW1B2KmT6Yfyd9NTQiFbHQwoCd5F1gDAg07Ogz/HSwPor5rWNCZV+Kd
SMNNFLwWpWWwTmw0DSjIOrL0BufotBm8QGh0I6cT2v1U6B5RNvxL3An0J239TpLM
nE+okX1072T2ZQiYpFTk5a7YLJEPNyv+ESd5xwyyv7voWqmWFsulXsGC50kaG2f0
Y4zWBHIK3fuh0sLplWu0J+ZVgvtXCWfCSclCHIIKAXX/i5eSlSFc6JBzJkA4zgOp
mQwWB/rY0O4R7ECJea+TbGMcXkDdhBxmfnMOUbElsvg+9fv1oJAQc6gws9jp4+Pn
LnzI0pJZ24GDCNHMDLHl7fhjy3uxHwcbf4LWLsfrv2k4wRThpVF8GlRj1g/YsH9u
Vr4SEyiWopm1A6BEqlb8b8ZyciCotk3WgZA1hFMZXXkJdUOS5H/kQQgHAsihEWs0
WUutRlvyU1DOP5nAGaxBzR6qo5El0kDuOphfhp27VF40ye+0cwKNzbz1MOTuGkNo
o0pdJ8bcSJ9B2Fosjll2v505go7Ks7XFbxN3V4J0eNW9e8kpPgCGuLcFdITF3cwi
oT5/o+vMc8uPRBRb4rsCInhzfq/XSPK/JivBvSu2qTmGh55qw2u60Ir8rDewBXGE
c1Watk+6L3an+FgPqKQyfCyDYHlj+JxkrD1Mu8rVwK0TX/5VyWijZYOmeSEBEAUk
QaRdUfLCaiFR9L1wEt69Lv9oTt3mzUwYkwABIvls2b8rT2p0MiI1JEw6lKCTWT4b
5Y0H57Jm81EBmvLl8OnjRwnF3016Jc/XHEEa68PrrrwtipRZEkKAm1KdmWqHjKhe
Vm4uq0BSnipTn1qU1ZPC4/f8NKt5MdfJLKWHRku2CFTTH1OV5DrbN6bXt/zAGdpa
uflIiLj4vSJocIzVPqe0gIJFOJlccnMfPD3+lnJXQRWwml1t/0Y88jMZYR8lksSi
rFkmKO0Jks3OGqKgBFSQMdifjT9FSPIjCLneFJd7Oxjd8E27FeIqUUZObK7FMOTR
PfrUDxvgYC3tNJYPRJYoQ6qi3MKWi7f5SxaN5b5lpTkyA+TXinV9W9QYrInIgree
RnMBd16epnUyssYyhos+cy6yFlB90Fzm8anE412i4K46OjOQo0Nf+NEtXXjo7Vn5
QBCdvUV4olE7A7JvR+tv7lxw/lftqI74+Cccm17RneO9YM4gF6rcPHYDEd/0qNuU
NYKAaV+kx6ZNmM9Rk8YOjsssjgsGzctoORiJSnA09VS0yNraYKYIL9bg2whKP6i+
KHgxtv7BJtq6v/RGJfdpPqvN8Ca9fftTCpzpCUtf9TdCzJ7i9RVwt6nrXI3s2hLc
xjZP1HksJJZzNY95Smvf3LAn75sgWWICs7fESF6DiBotLcmhoNFu6IHn8whK+f6z
8mDVj4E+FOsfdPAhZGFOwNmf9GCzd1Dk550uZPyM2hGRnNl6gRMNUZiOiw1PdKPb
r9oM94iy500dLOtlQ/eCBfng77UmjZ59VnPdY3AHMNPWTCQPmVxFnOHYn9ayGVSI
kKUrLPOXytMut5ZaghJi2ikIl37L2PhFo+JpKmzKKBPL8JMJpRwW8SoMEHaO1SHJ
QPJl/B5yn8xtVpS1rflOsFkg0+6wEateuG6gZ/MGXdkYFkL/9/eG1Ft/Q8xEbDfc
MfBIXGZK44i7FZqvFMkD3cC2MLSPbKYHBouhxnhf71p+C4JBOb76pM7KXUjOZYss
t3aAa0OBtNEcyXdsjUMmQ9AW4w5N4LekjySIAkjE8m+Eo+0TvwAETbQ0JH1IidRm
rYfyUptJAMNhNbVfy0OaT8OCq6KxlXY4IRHDW14tL2k2/2kctnwl7MXOLpSwZKOi
lXjfcDTlMCR/rgWrsDL4vR2NMgNzWuh3Wyay7IhGtuhkk7HOW5W00PJdHE1boMM9
ffobYnX9pqOvbDwyq56s2+cm4cz4frCE+Lp561Es0886jxWkSp4f4oGB755ls6/c
nslfAEL+pnyOxj88HVMtf/RYweCSFNqiPfspONwiqA8x31so751fza58S3+aAVdq
E1DHJVRAv4HVPRFWO+N+WWYQ3lmJXrtLmWlIaIr5EEtY/c4ivztMaqm1gGreM6DS
HMoS/IQi8dq3QaI5LPFzxWV/B31OgG/A+Jpxa1gty4COGCWnmW9Egqqe5P6LqwWe
giOOyzsV3D09AWYP3fSXB8XANfW2trzdSSuEXXE6Z2oq551ZHYIDsZKQH92f5eib
3Ep+whI+/abpar2UZTFUFhKPX1X6ATdOOSCsNCo2qkvjuxPuFqRw3TiMdYrYkTdJ
Kj/QOXC4bytMj7lS7JunzKv9Rljpeqfq2O2/sH94Hu+uLz7Qwu7uCyIkWJTen2EX
sWuHWdbMAicYnrkjzZ5eS3O2kWlqaqJQqcAMF94CjNdI9d3eylT/gUtl6gdOBBUM
4EQdmXEh6U/sJh2xbc+G4+ktRDpzE3o3VARPoX96sjJutqarhSW3X1ZgEyzsGExM
DJfDtFQq6fnlglmCSkcEciN8N+mOsFNrYaD3WFEZek21n15McwHWivjtZodBWtFE
C0uXWGHr8YYItZABGljwhyWuvDwQvWvjej/FybTcTbSL+Obu0x3KGVUP97RDedxG
eF3cXO/TNANBwcFueHqzPQKk0+CfGLpeu0NU64AD4+hqMpLjbiGaQlW37+jkjolc
qRvEaLd9GHa3sjIR49GGnDtVoYI58PlKw6x9fV3HBurzqyISAPX0n4dH/1wMxygu
6DfoUOUGkt8h7tsPjLO9oI0jlRr59YPPdLoE/oHZIF0OnxijFmDlgsJ0juzdohoV
Ggj2DclYNQj9BOtQt1s22lVkohAGHHadIO41JongR5cBofamc6tik7eWeSgzr42x
0ztPj5gzNUIGL5vacrglhSQ6GkGzsnw9rlhnPtYdEMHYEfKQaOiIQ5uTsGOLQZYJ
v/PKFw9JmhWVaNToXm+1n/wUagoSoeMq4Azr9CiBWTChiuyevEbA6rnnTl/3M5V6
wZe6V/uijN9DafTaxzqxoC1B4nwVIN3zCvKHdVNUfjLWL+qO7rXG6L9yfkEuXuco
6CHX5rptcmH+LPT9WuceINzUGVwHGsEM8abf0Uc2mugodZD2r7oSHPFLR4xOR2Lr
4dEWbMbMj/5tMUVKnK50XEhvqHXFavMCc1JDwxKfqBsmLlShlNgYJznn9irgCuEd
/CRbgTklX7DYnaCft4TtLgGvXdd0HzENhabL8sSEIEMyL+MQ0yhitRhIEqVSwkzK
ky+j1+zm9yiQdHJjGmwQva6Fxt+jG4GyGVBevZa6VVO7NyQ+/jzNqgIXVg7awbFx
2ANkdPa+3zFnB6/rL6Lh4r+A/8D9QKZSR9SdT6czafWoLRZ2oeVAlztdzzGPSLKv
f+jb3qz5BNbcanakoKULnCz7C4z6aoMOsn9fu44We/H6iUvcEFqhBYHLys3f93wD
e9K7tGczLuNsk2gOBjRVvXpulrFKnhycW6cr8vLTmQ0+WjtJY0i63dIsVNt4Dc9G
lvAnQz/c2PAwsbE4Qg5oEYutbVHvwcu+lRnWblZVC5oWWhFoSJzojVryTJmLsK65
z9FgomVz7foCpsUj8ISUxOfnx/MmdxR5SMYU2KAX7AtucBldxrqgucbrUjOjZD1T
xT+meG0l6y9UKovM5fgbMkaAUaDcsclx2oJD+/E27cOHiYxxOxwhCbMArGz+ia00
sfrXS5yueThVMb6M9VSjpmGBEyac9/BtOrFI7dDFykm4bkFOGfsH7YtEeoOlpfuy
sH9TpiFeMEdOzvrDxZOYXNvxDvb5aWRLK9Ik91R656LcsIQ+KjfJD0tMakMQH+xL
BhuAV2Jx3bhrkuhsveP7jwl3UFaYVf9tGZ5EPj49LoV+GNhjszu20Edf9G6f0XFj
mWTsY8AT8izE49YXqI78w6kz2bPXfQFqM++GfqgGnLg1D5tFqk6PMNq4UDIOkJfF
UgA/Nj2YOPQWVspUBwW/1oLaUMpvg3naTPdalAlPcBtIEtGEupB+ugoxcI3jdCpG
BTyEvzTFYZPaj5PbUkPTRisRccoCX52U0ws/oCeyfUjKuLiuCRLs6oo5U5v8VrJo
lOL5DZE7GEq1M//IRFMOO+bt98qDYoqFm3QSi0mfEYDIQa/Xxv/PrzHxUwIINojy
U2jYY4SjCsLEi8gB5dCNVPLSZmpQkfwpfnPkoaaqeVg0rryTprzX8bFiHSXaAb13
IL4DxB0cleJq93FsnfDv31C6v9kT3AYFMdEsjkQkNBIRbhb0rLqG6qn2h+p7p9e/
z+dDX/9lMLbILl9VDZWekF0QRrYPFZHwp9X6Xc0KmatUPw7GU5IEjKqwDCWfwLpI
7yYfGFJEFliFONPAxcrF8I6Lvomu/wm03z43RDOjP/pGK4yXv3fJA4XsRUy0dCcR
4BEkjyNWOpHijhlqpLR6bYkaA/v/wSJHieGFg4U334ithGN3nXEyNSugTwDURPKD
ZvzFA5YCC0L4MHjj5TeRN++y4bkmDHJgYtqI8LPwZeVC8ywos6btD4RITYqkhQPn
jf0+9/EMu9qPGj3qDmH+7p0+lWutrgK3x32SIegXw5jeqH3G/+tZ+qa9mgKdUsXn
Ug6R/LkABXG8XUwwE+9zD/vcPGr3QWjQAcBiRg5x52K56luOUFMtJs63kFhSlkLm
dX18iCp6LOaiGWJXkEi7EWewR0+8AdKgShBqBs7K9apXHB2A4Yd15ii7oPRGKl3z
C9vXZrSV3u/R5fUjhBw7UBo39/V3fvCvXU81Bn6dgbVbkmZFBHG4BkyIbuyCeIrP
9nQ/b11rTOnx8QYoxuCoZoISSrBMVmr8pm5Jr5vCfv5l/DyEjJ/5o+730Zdi8zSC
U3SlXpvgEMXakq0uLGDMmd/PY2g77lZ0uMeMrOY6xSprWtb/twWKZL3Afa1BOQ6C
K4gKOfcNGrX8RSUQC/CRxtP4FhDqIMp/drwj1r72/sk9gyI8CEU1m1g+MjdQw85V
quNDwtediBg4Cc5trJrxhEJPMq2ck1LfAHZdnf8rUUgAAtCI4GD/khLpTS+8AKr3
mZ7tXijs64Yh++RT+hsuY3ZZQyjYhqrf2q6FE77I3LClIzoWFuIP7uQ6H9boewiI
C1BEKH7l8f33kn2JspnOMUbLNxh9PN4YKs7wZO2UmQLP57t29XcJ2lHCkDXyfsH4
k0TP0Hf6prjSwn/Upx+XD5gLuU52m74Todfk1UQzS5II8Uag01Z2IJbbk76/fLvZ
XY7lVUVVgn1EzcuX91hodUA2mWdsVC5TkC9JcGcMdkS8QeCPZ0XDt3U5K1XfizEI
NhBz4O03nnyjFe4Q0g2rvTSgEQpdqI/WuxGlrbdfx0mF+t/+MPVOLCh40Hll06a+
ZWKtwi98iF4VpMb+xvR/gNv9bwxpqfgwjq5xoL38dP5yehCcvLJyh/SluCjYOBJj
w/biVfpYNvFfTUJRbFxVRJ291FC1nIBVb/zk2q9/00NbY9QcbvDVlB6JjUZizwtg
LrNQmQBRYA08MKI0ajbHoYsvz5R8Pu0V/4/7ywuzn5jrQlYOGBoee7J+wLka8JHH
urF6rRKoFpasH+TOluI69WC3Ot8fz/HIaFOgR5yDkXAcjncpVrpAW1GDKinVVY+p
uR8PJ4r/Q2pzT5cWD/SKPiHeYui0MkRON7oY7aFY0n/7vwbmrn7DlAzZU+9lN/Ml
yf8YS90V8kdW4jreHrM3/FV9ZTghKN1waREgHLTxrgJURp1/hXyb8IpPBa+GW5N7
rf+ogaGWvJjYkTQhEuSxkf58Tr9fSSs8H4ucYsYTjPIe30+6lkgoH15aNUpMLCFm
xzyD1kkHetSNtdN0MrvuvXIgd3yI1DIh8eLZv6OqYWzNSbsKFphc09FytaUhydxH
uwAQkzqh0kwJohIi7F4so/WjFSziEfnA6E7v8FKYgHWy6qivYQp72bcp10sjJGNP
ZU+nUK76BIjBCMvXtNDY2HcNLX4VQvscDv99BfgXJi3RsivAfU5jg7cCYqr6mXFz
q8c7E2QRfI8ITsIkBT0bW3y8MZmT6GsGgSGZtQNDLT0zjcvm3xbFXoW0q4GZ0D3E
s08T9rno/K2tYkY1kiU4/3KKH9tfJ+Lih4LppqJTKOdOSTHmGIHnR3GoSolStXMs
cJWJ6lb8Fy+gUm0USV9KZOLXrPdOrX6UuCtJ4ECSOghRXsqHcpjKQFYx17RPNOaO
PE28fO6pft3VCiNmAwoY8H3+HdWlMqL0Zj1P0XSC/cQ4VPiJw4UWwXSGMCpHIj4d
0cJFKdWvTqSmqewIGOnjPgW3Gll5/GKw5FdiSH2lEKN+VDCQ5LSRGoLj7oke0IUi
299PJWG/2hyZaD+IWU5qxmQY0pT8yS5/+CcOXTd2aXLsU5068Mc2v/pS9onildXp
rgsZMeyNDjiBuv2LCvvLIgW2WyIPiAn4t+VAo9tOgQ69Rvb0mNRwjYAOddfAyPtx
w9nRnhrTpKMvdzdz/GO6TCxS9LRjfNbdo0sS9Q+tDeDUrxSx9iGas7ZDj8+einBO
i8w1mxM2/2DBYrqvjxg/SL9mvokzPIx6YBEU6sS4by5WpR735x/46p8WqNtmW2WW
bUzc4ugWXCsjtY68PIZ/RZnCedE30RFwIv08TzmuRpN6wU8h4hOIDgpP/sf5tdU+
Yy+icdkUjxt5bw2HINo54g312mgcchm0qhDXWqVKs3IGTZDbf/Zh8FAF5CAwCdKE
snpQ2vUfIIUGvl0Ip7VgJagHORd9j3tuEqWh2VYyIDIkTImkl9few7H2CtJ7Rf1G
3FhpT0chD0+cBNY8vcGRAhPXoGofYv5LZuWDpCaVqYQrE+LC8W7C1GyL2yh0YwKA
IvtlLj+6495+/j07F6FvzVcHm/8UgcUReWv9RSlKmohlUvaPJEtfz+eTn8ANKmMa
7NB183oa/1xpJSJ1/PQCxRTf6oWNXjPq6H5P7bLnPa1bZNDuhHs02jGuU6u1FCCM
9r2QArHyhGM5Awoc/3W4t4kq34RisvcFsHw91jzGjj0CuctWKy+u1fsgnWgMCic/
JEt+4D0gWj368PXEpf1oNPIzsGJrvkrwS6IGmOCZX4iOr6GHxr2QiUROfzPyTNHR
HRfq0o+zJe+fj3Z17XTN+O43cy40reqcyXkvsQ4Fc2FxTLw5/En5JFwBtEv0eG6n
MWA4qnrb/VCyhUcvWIX6I3TgTF6qeKllAeCeaQSnkOqc1/EIDTfZb+Yv96EYD2PA
OhIvzZni82ggWaM2oh+8jTdFNfTpcjWiCZ2O802QTEFiCnWWlNRxk9D5N++47gxV
nDM/ztqC79fCEWYW/jwvlD2Bt+OQi2VKpwXW11OhDNBJ7k1hLxMiaH2ILjL02lSE
ceXpwHgBazCZlOJefeB0g7lOjMgco4ntq1/s2Zr8T+V8wNryP6wYFSsUOe+zlglM
aEerPJ/gYSkX3R2341sAxmlSRctL6YQaKLx/ZAX7dEugbDeXiW7xZDT7+MPUsSH0
YN2uY9+1aytB4DVWNVsvIpexcO0BV7dFp99V/wNCtmXmoJFr2eJJkj3IWmqCXyuA
2EwLiGcQTxQZ6RyoWJ4FrVKKjDLETZFECRlZgTRV+yEm7AB2goDVkxSkj+ipP6Iq
CRS3sZBWhaDJ0ADoclloRrQYR00xDbv5Gu+/2prZO1FWyngydmPTayfEb3dUyg0U
yLWRbuYoS3isereIItQaYc8Ms11OWMhQS4JxVRxYtMl3X3LdamWlXWTnHqHzs/gI
wzmxKCPV9wn00hxbTvUeIhzWgO11AV+ByLytu8+iOppc4f3sNHw49VK0Y1V/wANp
khRW6e8hqagiKadVmLUN6T2cNKg/v8V9ao03TqIY3kVMJ0nme5YHJhyOkmgELyFP
vbJdcbuOtixEPih7ec7NjHgcNBRMAHGmjmp3sbJDD2/P6jkYJTT5TPmaGqvOvX1u
/B+f2yl/vm3KOy8KcZCvL8ORTwDr+qBUfvAhiloR+Ur8IenovG5zvLQT8yMQF6XN
HS6HQHabZdJ4oGSPvmNFi7Yr4TPb9U5wMW9eVHBHBZZkWicT964GCTcBaRnF2vKJ
R7gaPeywXlgEOoLYPNjQJRn+x+AZRlIEYYxRT5C9FGHWf5LWOb7W0eEk3klleRoM
ciSKkZHLNiHco6Xj9AFJNdiZw/4uDRa51dKj12qS2qPFI6MB3rJnD8ywbFVAh6a+
+M1DGukb2nzu9aU5Om9y7I34UBADI6d6NxSAMRXLeKUXGT0JX0kTgXKZ4aY0OO5r
TbhVBS2QI/CPLIg8Ti+x6w64OqIMO1igWMW0SZdsnNZkzdRE2FXxWLqFhOOXaLYi
kEOiHL3P6VpEhtbmSryMsrRSzwJ5lgHNlnd3pdZJHq9PnGX2jLhGUglzj20Gvl3K
Wsu6K7TyaCtihhEfaGjnXPSH6FKaO3z6oAMw1W7/S+LFRenWIjrT9JeXHX0wcRIR
j1Xq8nu2nlkA/X1Bg6McK0+vltj5GR42iyZYOX+BXuEKI9loMLcThaaxD7PFMiAc
vvHTixzXG0LcIdDJNV0FcCuDGqBFoQdtX1VD4sFcEKLhd9qA4FFyOG09WA9W+5Pr
cV4IrI/39obIAX9ktoPrCbcYY20KsUkt3ZNAbepfIQNqsb+QCT3G9uUD94QEBKTO
CjKF0xaF8pX1lABXdKyDtHFhCw6qnrd0hXAQ7uK59LILZpesAv5grKsV4Q2nWEWh
xLBP4HdGf3gZGjhY4SwuVUebHlET93r3JSsB8Am457J8XezMjPFBcIv6O7SC1/wj
+LFFqZoHwBQoqSTIWaLNMOya+0yocef2rgAr0jQmMHlpLrXkYudqTTvOA2rVc1tR
03d5fOqnew6JJfqsGkEEdT6w5jGQQVSEm1xcms/OmUD8AGmVK9tPCAKkR9H8Twwn
UPNC6uNJ+JaHL/NvXpUHfqPukyrBNs592dA6KlzXyNCsNgqyasUUzHzZPIZ+gU9c
ICwFAB0EXP6BH687e0kYdD91oQvuWkdzhFf83k+ppN/7n/I/9m8AMjtDvfzzOflD
vI+XewwBCz5kuxVDsp/ReJPDr0BB73kfa5vPNCMLPI+3rD4sqhgArMglJ5nrQPJx
sJ72nWAV+GHYR97uvEfIA7Q9eautWE5kTOJAiwz+I0EfbcjOKsGSQlr/3pbLL778
0ABSFgUqQMPApr9L3Q2mNWYN8EA9f/Xmpnb6GqOiigpC1Yq8nh3ANtUNkoC8v7Zr
fU7FYugoxy9xGiexK1zqM3pKcAVHcMZh78D7Tsirjlfz2NcsZtg08FMcMbkDjaEn
VWhfUvpmkiz0WeLZrlnnA/o8DeXJOzdOdQK5xpc+aW/Ke9Syfz8fNKzpae4DOWgl
Dte1W1zoU7WZVuHL4Ni0tsngB/cv69VyZ7Qd7p5Y+eoK9II33Qv5J/rARbFKCxDq
eGCLKLgIc/osSTcBlBakfdcdpSqIricVJsolh+EDQC5IKDX6tYxPgqPuIBLMZDWO
QZwl+9GPLXAcvaDyfWjeXNMpeBGSvB5bx2ertYbSiuxXjObVLp/FY/DYy7Ln/woe
rIRlByI36Bja0M6hW+18Ma6Iqw02LAwFHymeiiHXp2v3xtrHUYnAlYKs4JRvs5B5
ukr8wliBShNscnB0VsfEsReY8oPAB2jVn2d0ziEScrqeEwss7JMzCxHh4w5/l4jq
aStcbeTkZ5RxNO+xBKWIPV6z+FxIJ/J+GeaUfzIgkXoF5r1LawN6430ZdH+o9/yT
PiOU/yd0uGorvsRKWTKENkVjMAI8Sc50H+QN8kQKbfdu9ycUi8YAMZzGjm33lGrl
Bxb9LqHxALfzIcXXaA1pC0o4SIYgA+tnDPsy1WB0SvCVwbCz5FGVmVnMSxFj7XG9
zKtpK300DnC+OsMGF3EhnnXdjUe5Yi5OnVNt0YSPxSqhG5SrZ6Rkafqvqeh4tbfX
lJJXMMu00gjcheiYpFaa3g/NcoNbHp30f1m33LsMKkQCtyruVpJeoz7yKuRuE7/Q
Z2CjjG/oiUc/OkR/nzLvtjEXsUEaozTr9cNJAkV4ZGUHhDj3XbNjetcVtOZL7feb
a2DM2lGz+04kQavufO2EQB1WhQWqZe1VZMncPGY2LJV0hSY+s2pEIKlH/5iBiQfF
4816KVF3R6SuIWePE79tXeFcgwWCXJdWwDoXp7yJ5TCiVOWXU1GPkoGide19uVea
rh5oSYYXKSth/uLopLmHerNSaZ4uu9XX7nA5BR/dEyr7J9eybuQYPZrLy2rZ0pFw
F5TZGvH4yjGQ8vevFbUfvhN2SKBeuIQCpMFTdmcmadNQEQtXE1hulMZoUR4/HxZI
j+f6OWm75SbEpaJDmJBL3P1zR8ijJchauHfozTrchqx6syHDtZvhd9uEwp4GXNIc
yKFVeC7fIKk6HIxmT8jTS51MK+DP5YtLT++TBvGQq3yGM3d4fPqeqimBCpcmJmu/
qwLZkXwJRRfQRYRrZSRgIkcD0DoWXodoTrq2vRtfWLLYh01fm3iKbwWtwXgR8/rh
yHwa2q3sjJtYEsi2F78pC4NiwjTat4I5lIYj96ogTS1QHeyWwUceASvjawLveDSU
q20t4Xwb34EK6vfXF4Y385mbgrFIXlx3LmZ/fwdjIZPlemDTRDLHDMJyEmhhFxke
ChD/l/nN2qAwfQjCiiTSCcmw2nouLKXRIekBwRdd110vHkePfV70i08g6D5v7PKp
2hn3rZyQIUB02aTgLQk5DyTI3i94m00uNtplRQNUqSIkXi+E3tN/pWVhOUu+7JDK
DrV3DLxrdxTUzXwXwlc/JacaIfazk123WEgWU+FCv/QKv9X5GbHWAqPyYtYU1yqF
vy1G3R/AbGVGcmOad9hCbM3p2tzkdbz9Y3sqCuN4rBYRJx0XQsYIfH5bvz6y1PSf
UmYz9ajTWxLLh4JFbh5PhUN/PclubOAoEyzPTUZttjCzICDcrNsPYmwfdYQBawqc
ot/zqUTzeCdHkL44YSUr9tcX+EXcD3qF7p0vy330z/PHWu8YRH+YPQ2Xf3T5ROYd
fmlF8mNSTfGh20OjoRiacFSjVxwmIvhWXo88wTU03sBkFIdHuEJj8OdcUcU3Zl3B
7NBJ6+sawU2hrEZ9fQmMAPpD5ti67qWgbcu7EpO8n1yI5QzjHwjWEKyP6EZl7xMj
e3i78YeO3wkL1jZg1EtZy+7kpaJONQwI1+Hick2iIx6yVkm18m1SqJbidk7+CvV9
0oDeiF4g1gaarpQljdLtkVtgGIbIf1i8Fd/bP1AYImUZ4sMs9zM6WGy6UIL5hqOW
L/ZJS5Pb8kv2rdi5kn5Cv2ZkT4WlQpPmox8DJEhsyq3bz+T3yPH2OG4Zm2d+bU5/
n5J6vAu9N6BzuQQqUL3fz6uYQQc274C50qQffhxocz8vZ3wa3aP3iDsrqsKzd9+c
Q56zbZD8flE/a+OJtWYahcvpvrh1oDfi/CPlDF5GlTOyzbxCeYWH5zutabvNppOM
/16+I0nQHUhH3l/Yep/LlstbCPwZtY3O3NpZRpNjCfuS1upEfsGkoK+PwfcE6Ojb
WMxkV4Ocd1vUBEm5oC89Qvvx8By2vAv3LtfvyqJ4mvMV2pDZ5+RoqSyjHpQ4smHR
kAI0Tn1xJm/8D07O03JhxgkxEvWRk4a8YOkTWklKUuvRVcGlUKfdHLi6Yy33xEi6
+gp/IJca9TjrL+x65Dn7ErupgcJNmCJPwf8iWtanEoQr7XRX6FCskQd+t/ydra3m
thcbaCAc6YKQetEAmivEgma8zQj3zmascblBrRgvI1XlUPkycJaZEqvToFWDnXgp
Xs8AYFFSMmO7DQhbN7eYm8TS/T3hGNxDYuagEGj15kw26Epn1gCWDjOeKxWPAP7f
5iifkmTcZve7IGznXsBNFJejFy/ODTs3SE1+5/SB6cUGhiJJI53bpDAkRpr+gdrl
1kGRIVV3m/GPWHeObkO4QZJpFfKC3Ff9wwzOv51om6m4Sw4mXwAECq0llDpvN7e8
Wjv6gUqk/mKi/ouPs5LoMOSCSjX63ReXzm9TLsTZbj2Hpqqu3JoYeQaCnC5OhgrJ
aOWKOg+Hql8oK6zqhThWMFhu+cRC4WiQUwSUZDfGpJy8Xfp8wyEEt2y6UszO7+UI
iyXGP8mEWQ/EWujz9iXwfTV1yZ2z1YepySWzGqA4lfjdr+HQ5Hr4cooS3Nvp+3GF
d8VPPOerXCf0vtTxIYE/i1zIBf/XYPBCaVmM5TS9tbqWnQCnizoO44/zKQogb3fv
INvfZdKh/OI4n+uUnOImtRFYgSj62pU4LdszErL8LaLzwwoNuNKoCOloIG/JFVHH
jQOS/TKMz200r3e15zkhwoFAnTi4y0lOrJ+jhb2wOZLFaiuEoM165NQWs/AiuW0T
0eudBMwcJ58XWE/Zmya1UUrlK2HipoCOsqtr85OANEzM46+X4x257yISLFH3zeQy
gYfh4rqPnZHU72uxuECNMjhdas4MMCtjICq6ebCb+ZHkozH495W9OWELVDa04+iq
UE0ykiC5UgcP0BzQPGGhWzeyF1/JTkT4/gjwpZXpXcxo3tkhvun4xkuvyeb3dbUM
d5yO4m7JVZoFeCWCtNmUlUGveYXs/+XJ5fAQOfn2F3J8jb1YCOfOPwpE1brbSW/M
nTNtOLMmc9hxEKvp/yt1/nWNQMoS3cEOnBb6fP/Cl2iHkZ1yFWbCTAmXcJk4MhVF
V2BYwRYEgeflTudq/QPvlCjeJvNSxmmaMJUp0f64KEFVwZdL8sewbHhtw3sDZxpk
6E96YGFRFPhi0DlVOj8Oq7GG0Jg/ulx+h1y2ofwzwp7iGj5E3YdnnXxcLHR9ciLc
YVXU7RQ7ogvvO0azpoQyeggMfrg8Qummh5Hvq8jQmkAj1ans/qFWudjSe/ZGO5ql
Rasm/dJrhyW5brdzcdTA1b7gyOaH6vBCSuQa+AtKoMg12sBONUNvOH5LiQl3xfI8
sy2mPC/U3z6e0N2Iv8/mFoO7p0PCr+amLZxCPDq45eUVfKRMo6Mvqvw19e8JaiEP
zdMjzO+5YBjpMIbPXWsmcDlaONkkIr5Ic0N0lqp0qZEMlcKOdn+3TkRsUGJ2ln1c
WuFqoIONQNriALKaB7ikWF2eqXMdd+mYa8CDL4+ylDvyblK4YXjyVdw5O/P5Yria
88p54OhmsVgaCpIEn3fyVKj4Ie1OThCwv/9uHaa0/fpq/eLP2kucomLJpLVKAyEK
/NLQDuSXQ4PhxtzCyov9BSj4M2alF6co820LrEK6Jo59qfrY1iEi8HvT1PEeztnJ
RNH8QnacuYVgPvpvuBsWgeoPbOI02o+YKDVDvvR2NN7oToyy2DiatQQtgljRtvi/
y8V/SULch9VFJRBFepCeBCOt+5wy4zhbvLG2l3Eb3pzBIair8GBITMpg2J7hsBDa
+nEkzWvEg7ZqIOvK5dU3mg2mmvCB7wq+KgUsKSI33htCs/NUMFzYoIF1a+tPoMuA
wcTGVAfYoVKbjSKoZpBqC1uStryoiwGoT67rjVcJ+u+2MYrAqpQ9nNGXKTt6z7cq
A+Fv2edpWRcPRYr7fvTCahkCCmN5hMKwMIgmRrOeukodbs4mHvNnpxTNE3pzhh3L
wtoIZWO1CMVIIHyADpCdHJmbrrsCMwqn3XJlViHbUVOK6rir7K1/YQ39BtscHOTI
I1R8Zh51rZypGs2ntPRunYconGFZmx3rL7tvi1iLH9p5fNWuAxBUItMWby27cX7N
rkp2wU48UmII/RQ1Taw/evoL9BeruPz8/Xqkf5iPYXeCnqXLGN7GqD6KhKul+fCN
AqpBHO5xWWg3kaYiDkWj3m/NsAVIQ1610B8mBqFYmoZrlf0NhG8izi3sVE/L6dJW
TvoZ+8jXD22J0aPmBSpG2ACflHaWDmXmqDtDh/HEZxtjJtdH7OTAfIqiQWD3pOi6
uLmjNtDDL4BoD14IOZKjHuB7fG7N586PGfnxDmghCDiLn0ff4XKpMlX9nUeIdm6p
1pnEhKDeDyxkBRfpxlNRFSjebxXyr+0nbc3xItNeTKY9dGaUKRIhuqpix78faWyo
ukYR7XQHNA8aEuXOUb2eLagHPEax4muGQmex7NPv1c2JrxPX32M/B1RyLPsfcpfz
ewDG/UUUAJoIEucj76qyvka7hYdXvbowPSfzDC6UsX2UaVX/R68XqFhNQnp+e/gS
jQg9VgwnG7TdHcZQfB+Rn545OFq39EuN0UHDQ9pMQgk7I4qX/GemdIS13S00Nh/K
ZnPahd6uoqVZ9DFZ1HZh/nhsuX+YwrUSYmjmlYxsjNuqfL8BW54QuYI1ARZG3Ytn
zid7bJPn+XQhyQB2GPPneybgUwiuxmfuh7ehatbFUlxoJiuelq24Dn+rxcFsJbc2
GELJQUbSuHU87XPP5O6mhi/GAQRhZ/BP9oW7B6dx+uXomY5MPQB7jQU3hC9Gptq/
fdb3e2ZMXrbxVCfbfbgzj2PRq8TSmXH/e7c8uwvCaHcmUtupagYh1CEyENxVEC4b
e9VMxaceE0G57xLWnAWXQZCgBuUUYWXFSiwbVZuiQKiJUD+d+COrr5was4uFJ1Ns
OC05jeQAfU4c4WlbC6QBE8pNLYgzC0dKnGEjNf1eQykdrJwYFQB5bIoxjpV6lnNx
jTKMIhyMg7GhLNy3ZdhWVz/AGHsBy6vZgC/M9z6xYK3kxpnOVZfpauwEW61ZtbsY
JkGM23zGQmPRns2706DO1+Y8/c3RhU8GscsolbA+r/CWnGQ0+9d3Js22Uq3AAXPS
eam6h7Zv2ENNL/Ro7+B5YGG60/XiLpteFMUsTs8crzycrAMMZ1cfa3JR9GAfk7HD
YqMXdhDor6pCqKOzbKhqMCckMj7oOp0RYjuV1HyA84uus2XBTUKlWKA2T4Lr3pcZ
yX9ogH38koBQYgkfJBU5arP5NZthOSZL1j9aiGGNR80i7Jkr3bpUvfBd78LC/dfO
oAciLMdr60oasVxwqcs5uUgjz2aDzBHyIPlyTlQnpGbCalikriI7pnuxhQo2hgtg
z7URPvTt2HEkYbsjBKsHLPuE32ZIA5ZXCsrpSMG/wiaMbVY5CSkAFzS9+IeePHjH
FKmrmU6O6HE4w4qzF6lXJ3TvpSHyc4hA1u1kTdVfJDrcpMMQO98o9IqEIlx7HhUq
leIpScc3poAEhCjE2EPY9IcPT5awPWFaEahba9Ft+yb/G+SbUccl1yHK56o/nJ4f
lvTCD7PyNuONT67KO/9bySEe4EZilQXTfyUSckujBxZE7thqABhJeRPraUeJZpbN
xE5B1ehWJSEssGskG3pnD3MbBrnTAcX3RYca8lD0EjWs2Gt1tGBxwtbGmenDdVqg
ucYa/oX+WgtEIbGW0do30ERTbz37amqtWjiS08zT45Bm9lFZXSJE7Yg4uFiLzLiF
NnqBA5lDjQI1847+5ydXkkuRrG+7uop3f9p/G8fmLShb8/ZdKWIXQ7AzYZeouI91
oxAApOb9VEv5SZ6Wz2C/1vTwpnzDVe/hsIizUTSIhcbmqxMsjkPgO92p8VQOx7+K
ZdVpN0OEDl7J9huVtanebYVgw1Mm2BBj6hbD+PHJUA4fvym/XgIBjQRL4rnKzyP+
e71wirmdvZbmec7HiqMDJLD36gcW0I4CtL3XoHJ/ZfPlM61hcTpUhLnLk/k+bvoX
sEsM8ZVxNra/g4zs2vwKm+X3PSCqloy6dcWurlb4w8TD+UJmsSRSOOdJbG8A7hFW
4PBOqS1Oj2zlet+yj4BY3P8+v/kaM7KPBUvmGSOdZ1L209z8lF8ZcpQjQngCzuto
eUQVA1kooiYsrlI74lYHERDOKb0xytTdhledww+ENJceM9wurhmom+FuELDGL37l
sHTFV2lZBet4qU/JeygD/K2jxSb5Oi95rAqdvwio+mlUhSco8mmwuXATCzQ+Qdwe
FW7lDcE9fF/stwTCgOZA+nEI7bzEAKp0dEepxK0GILBSzFY/bHcQuXkrvHSMaDeV
JlF4aKS2UMsKHrtZYm+5/v8UymOmCStL0HKigGxSlJX/wJrPQkBZjTJ0LIC3w5Oc
OTd8LhQZqwIpWdlhEFQcBfvfBgJJvNPym2t4SbhAud7+iSFgQH7+hvcRDIeUAWWn
QBMfpgWcFPYBf/3JexOJkn+TifU/xJsuF8IGkwJhvMkFwEHVr8wGGuEezCQ1dBMk
kmjEhNx9tVkgtj9W0AGn4ghZZLbClbwRXXofUU+pk2Mo3rQRElKJLwiGJ278taov
I4M6EAfpVWVEyIbUUa1htgqospPy0qnUJnzsi61Qg8UYYXu/UbvGtkotWDAloGpc
z01p/fEemfbjlyzlwmKfCGBi4kXK4WaFwmeRWGmaS4Z5f5BJAX7e8LAXt1JKNhsT
Z/RA60Hy5y02HGw7Y6HCW1UsY3ywMG2K/nGqQFM6DGCCRhzbAgiufbHC9fTUhJaS
84txPcP/Qhdk209zRO6boIlPrNKRYNegU4RiIOqH1Om/WHhUwTxp5tqaaJvopGNN
cZdW4Vf1wVIsjiyNUjaGh3pAnUwKVcSULImG3VOEDoaPk+XWSCgi7YTvIkqVvQnc
UCccBmDGRItzYzeU4kz3ARAaMfRsweGazVyo1VYPj4rAVC8yYsAnDHflmfXmRgj1
EFLwpZP7MeHTC2ZD6YDA4NTrAmpWgkADZAd/rQbf6Aw47w8sFjj7pvXV31ibIz9J
OiKT9qhLPS79cAJPr1+oxKc182vHV1h7ZmDqVolOmHSy24ITUXj+kzcb0I+P1piQ
vax2mC9DX9RQPwa3gpuo4RCtmTjIc97D1ihwqW8/cfSDs13+FzKhTQabofU7xB8h
/t0J6pPKHye/KPWo28li0LYdoiu7cA+vMN+iII2W5hCvw1ahcJryF8vnaQr4RXv1
w0/eHsM6DqdIG/D4qbtefGVGcoAMTTcUhf0VVMvLa4vMV8HxO883eywYHEz3AaIF
uAmelGdOjbvIYB0ESfVbP0iQVMsj3AZ2O/xgu391/44d8lYBRVKCIyJvIg3xqo97
fanQAtS+5wairvk+uZVjRX5G6Tl3GQtbtMkE5Ota3inxMnOocddpdOG0jROlsfrl
g4nMQ2kRTGuWqngdI7gOMkkd+kXWPQz5hYRvd8X7cCRXh8CBentQk+yVzKRwCtWx
rXUDowMr5q1/0+SdGJ9FaVKKdBUAizD0YUyFEYRRnGVJKth+Sz2o5HefBcDldDKl
RE/EDrSLd5E2vb30AoI6KAItNFGaCGDshTqXoxKeMypPgjEp3RAtQRt1JTcGeH7u
fqoIyHhJU1PEVdLJqaVK6GKlsHqt6XmWFHszSSfHnmGt87ZjJLCmETUzDYWavpJi
CiLQEKZy5q7xcGojqvjNpl4j5CBYaTqYRvYRxRtUnRvfeWv6fOdxeNGT9SNedUBn
wjcgzlJCSZZMBRmu0VN7S9OB1an5hA0IZOlLZmYxW5wr3xZq3Qwkna+YT9tim4ra
S4+9yuVKaHaSjMRhAQrqcH6r6nmQxkIv4/HKHe4uGgoeqVX64K1TkRQUFypFst4s
qUAjdzjX6lQ5xuHdb7U2dQPQhUVLhAm9VUFFAtY44dQ9ChUNgRsa0QWS6l2TB/vL
vHbMmO9+F91kzTKXCCc+/YHb+U7Rg/qCs4JpaG2VVjSWhG9N7x/H2vyjVis++osc
sXz6fBd8x6y8UrymVEDGbGInMXMzu9ruichDnEaZoYsHR9zPjIdFaRiOEg6mO79e
B7KwqMdFdvINSidfk2cKCGDKYPexk8zyc+23pjDwUt5kcu3A3hZTLwk2g74dAI8p
96oiQbaS5Dl1ZFi7Bxu7GQOqH8YXeQ3jVlQtoYNEcTJjSLQ/C8WGN1E+oK+KfVuB
XDdo0q5oKWDYzNKlpvMWHwkxzBDewSGL+MYqTkLtZV8CreRCzuS6rq7pDRcc0AW7
yVqPceKRk+bvkkwaKexVipT2YGg7JvmDXtyG4zwxaDUJlWdJgNF185RG+dHfmE2R
rgBuXCjOZXb7WkmoWY75Y1IeAVDBeFP8HnULQ8xgVfyM3YWsbeIozq4oaT1Cscio
VtxilCggI6OZIrB9Ufbm4X+XtFZOP2oivWc8Q06+pfH2Fa681Ii1sCXTGFK1GPhO
94qfixwGOTOI5Bh1SjzA09Lq01rczdrQhDZ7cxmx7GpFTp5DSoxseznXHNI4vCWg
XDzvY1XvxXOaqwpTp76zKE7X8jDZgweSzVb2edMFTTOwmQdYsNGEHnU6soJU8on+
Ygfp+lIl97ZGdhVEBpLTVvFE05J62XDghPnYMC9dqmNs1N+ncsp84ZNJd8CU0IEi
RKM0VqLjfWMd++2FAwh5r3AgwgtywIig9lf/wPxy7BLCwJxOtf/OdkL7SjFNzN3b
S6lrs9hHW2h0XhEQFlHS+AdyWZIstY01lEnNDWAW/L+Li5xz4zY663T8Plqph4wY
0i7w7uQupXTzQMP3tbWliuFGYBIynquTWfVgCIjzFP5/nt9VZAag537ckn9Lfcpb
47fsyoL/HYjYIF9PhnxWXg33GkN2uvWBgiHQU00keaNFDdlIs+f5r84/3O76px2f
Mk/znfkV/yGp6/0y/HaaTuiAZSc17XyiZyuVkXur0ENEWUQtnfYfA3Rmn0Dz4dZI
bw7768KNaWf1U0xfAW+4srhWdXp5y4R2OoY0GOzCiAxXyv5G1AfdyRBub30b1WOr
mhXo7I6oG+q3Y7jQWPPSSW7vqeo+LwRHl5SGNZjgtP6DNNGCJ5neFvzlzofbGm7i
giyJ3f17ChsSmewW/IpgWTB5XBYQ/raknQklsDnXpxiMCujhX8oGE0LArQZbOc5J
+0xtbZq7g/S/4/7V1tZgJa9YvKY7BNUS6B5p+PCjorkI6SprQC39RtIYicZNu6qF
ObrMmU6FGAOUXvdc5MvssMfTWTp0X9L4G13THp2Uo3Clm31KgSxH89wE5FDTLhOV
dm15hImzg4e6pdKsNWF+xec4LIeWvTUzshRYlkgkg20hvwJfuRbFY0kxOD4f7Rrc
C0PqjknlkduzDPNXfs+CUH2H9z3IuxfQZjjw9qlIJrexQELtumj1I2V8V8sN9F9e
YP8rbshk5h++tMnbsA8wBfihKa73gureLCbcBMfLvrKzi5uLTE8Yw1sD6VawTd/2
qqdX4TpsSzprtzGQqp1rzr35sLzBXzPTlxcltR6Gp2e4R7Nl009gcq+3gKilk2XK
V0ULCCULx8Jc9gK8voVZl+d7zLe1ZtN5ch1DLAtUlDVnv8nypIvYWUg7UYrWdM47
ABp2xacxOBAFveZyUdfNKe8ucfyT7McgxEWYd58v71EbuEOCN2X1Og4iAIJ3a0ju
XCemtRBP2OeT72+YHZ+kLP0DW1Pbo9AjJTdkkjiW+wrov5AKEyN5qk4mCGIXfN84
3vMTXAxCLGNsXYrPnpQIKBYl4kVW4+AsAKnkr10ybj3xg2mhInjvfjPArVHZ3FhU
eoUSGm19U2mzNAAfgPAsXiNUtAndUymN4KshQK1axK9wg0fKFxNWibnALrwOCgCB
rpG0q61moyLYMamtNmcwCzvTjDKtTxXsbkOG9+gonn0zrGlt/SHrlVtnxXiw/rCz
xYYNrfHMq7k/cUTohbX7BOThEUh3Bf8symgFATOMIrEnlJo9Rw6SDyhc3DswQYB/
K3I4syEkSxMK4zg/1iNnRJQ0l/cL2665TMim6r31d5sfCXxkedTs2juzgNFeCOZ/
wuGjQK9X6P4UWhFPsn7O63KZ+xkwhQ4bEd0gVcMERqKdt1+QpYPKGIQSmoe6qNrx
i3JGx6qFd+oHxxMFpjYNj3FLn2J1PB3TVsb814WTVbJ8CbJN0BQFoe839Uz3fX6n
PqdRqQoaqvT5mdtCtZsbHluZ5720K4Yy0sDHAPZrbq9HqAfZsb/0BpKO5ucuSx9I
9U7nNXgLHlZOpiReca+zWreMtDGFFgw3JXoIag1DV9zv8bK3ChnL69NL5aNWRreF
D1sF1SwGUObNrOaJx26URf3++BztllQWuqULnDWDUhA63QSguFPPTOxSW+mjiRhc
J/3BbduB4W7mdICYVb1qiNkmKk4oqBw9OW3HK/PO900Ei5FYulbm7FCm5C9hKQ5k
DK1r9SXdj6is+7wVoxp9AIN4CfnjCBYm5q6oKjxuxehaekHU5aXet4oOFbfDW/bg
HK/fMBaYrnNY9SA+5zYW5TGI45SA9lgTQbqJrOWxA1JuM/egwwGHAEtiD0hd8ytw
x376js8kUPd3MJMYUhu/AMFvDFsBkL8OBYhRkA41I/L7hRLfg2zDNXMC1n4Z/g0k
/OGkxegm/+aTdBkDcWV7bB0oqsHRxdDZG7kzIWdr6WhRrCKnItwkrPgvTczKMaGX
vSgZklnbVwTdsUfvAG7ietf5KR18YWyusQ/pN3+uzhIvQ2bIMewRnn0Yq3XzeSQ8
wry6kO4iT6lQOfI3mAwC66YZ0XLjmtQ1BiEzKVAqmUFZ08A90frDWKpoVDZQwVQj
jRlQJak97QjH48twUnkXOSvn++LS3vBA6sM+BL6fhcHZ6GxqmpnNI6AsllkeJNRp
pTS7BpEWWOpSEQEBPl7+dT51JfB7IIp6Q2uOM0xoDLH1kj/YY2R8gQIKRPs9zVfu
XtluE03U/+/8aYfMopDIuxaIsuM1a998LwdWCJT1yHjZzWVqssue7g4XT1iHzQtG
7t5jtnpBnd4fLIURlFnwR7iiyvCo18L0y/jCJ+OCFT47IfaUoo1h0bn7BmMJ4d9A
vwFmT9j5boB32YBbL01WtSob9J/nE/46zNwfPLicFKMfFXui1V5/kS10A+pOKyV6
X3hTCVuZw9VEJR3CrqsXQkFY/GT+izzbiRn11wkBku3zzewoRc9uWuQMhjEm0IJZ
ijWM9ToLbchvOwSEcgxEdYPiFCrcXwCeBjx/XA7KTnKPg54Zjgm3FXrLf8+SAtTa
GNjEu+N5iCUmC/UQIt5kkGdl/5+eAWSYn7GIucGw2F5hOGLiI6yUukTj6qZ/wuIp
Pvme45m0lgBunASIaogjkAo6phPdjXPxUjM0sC+aRj4YER2Kf2krEu5TJ5HQLs0d
X5Urud4OCCd737KgOccjkkBI1FfYImy3i7BJFjmVIhjipqU+y9OHK9832gSO71nO
8FqiaX86DdyFxo9gBORCiULA/3DinthHstJbXOXYQzhnd97AVBL8yuNkZA+mdDZc
okd6BybDUnWCHfRCrtg6ObJELljTTPx35JbXe7S8kU66gYjTIEVa3yLp4RAowGSh
2uy3W2j9JUNyoJpqHWlAalRNmhjck2dntKPQ0FHP5tqeJ9qysIlNGgBFX+jqXczj
ULGnq1/zX+Zb2KEVz2MFpoeXv0yAMJwI0fJM4j9uJcNkpF/0pwMMfqI9IZKsgLZQ
Q90/eNpjtTrkJUIGccUJ+mCLcMfgHWaHbSf8cLv4u6QwMsDoztJEW1Rx9a2/PNCr
PmtPPXIKtTQbtRyfDtXpV2jg5I09bXAWjovNZxfl/iG35rMyJQuF1HHY83oAiNXo
U9HbK0ji7FecQkRgPSMW4H/A17Rivwe0hqvV6egoabHA8nZaKvR70R8W0bLOk12B
w0lwYwTlw3SPJ1XC16ad1kbamQAJtpfZ4hNVg6LIa8ZLf7vbR5GgU2mRCGsyJIot
/CSGD4E2b/3l6sEfJEo1GABTalx0UOcWhgJ+b9tzdJs8hcexfyYdTvxzg8La9mu6
d2iouKiYLMH6krykFrbwk0AXBqkLdY1VOnuGtlbgUDazjIJjavU6jCc9VoPwbh9o
4H6FhXd9f88UYYHdODjlfg8J+7+Mk+qKCpJHcYOK1tPBuekqq8DU9YJt1Ci7t/xT
bFJrJ/E9VLEwF8uTvR0rPwrMlyQJv5MEcTkK4ecmxosX+KBn5fvCXv4Bbg4nhNBW
ZGSYMpw9RZNwUxJfyogkayzOWwIQVCfdZ/ZbrYVwBbfdHi84+yEiMpd47l5quatV
wLvxHWSNsQQ+/szK4AJsopJ1qnjqfpiY09T623fhRHlU2iNjGTrN3U37RQRGMxls
MLz47Fks0qOmc2BbH6tGtpue731I+zNLMtYdvuonrJtRKYJR6Su76qMlL8rPDoPN
AXt7CSMzLJNnaIXor7UexpQLHFtHH6ZeXMXmQGzYnrQpSxK2Bv9Ko3xAqMzJ5ZJ3
u+tlRfqoX4PKuncOsvMiFsM7oXWTshBlgKMAi/2Mi9Rxgxs1PArZkGhNUBQWJWEf
q2GxdxZbFSPlM2Y4tjtRP5DrsM6mqbimyQV9XXe5tkXomVgl72i24gJHY1P96EDb
oAuuTsGf5lop6F8dn9GEKEnntClqICki42WD97vQOlZ15iqNLVC26m8xE58eEhwl
oi0Upty90Q/gYLbfdHzGaX4KTuG44iDT5vbsVSceY98AjjndKfe6xaCmvKLRkyzY
iHm085JFx9HsUDXiD2C0VBkK02pCL7R+IGTEcF6XIVBDXPd/mJB0tC/mlOsB6zH7
kQxpRe2fOtGk0Ek5T0VuUf6KOo0TdQJYHuzNI87ek1FP8vGdSpemMWszn09b+bD4
7lKz3lalR3DaEVKC9+DFJ7Pck8gTGI1jgUy96ncZKmDG0mXRs/KOil/zeIfRZbk3
ObjXiSKyT2i6H4LuCplxCaj3vDMWPE6reD6ZqGtejsdUBhwK9O3vJRwFSHPRIbnz
0S9k1qUstqF4YCGswJBeOvvBnvNLRzKC3yh9YPkRprMjYuC+cwfr/R+GG7Gf7mI/
YM0Zq9k4NcC+17oTZ9DZE81bykVtVEMaLbwJ2Mmz//p0TnawwW7lFZFWCLNDuuVw
WYxuP1KOLPpNhyWwSLnLh0zKvOfVogGU1eQug6HO9YhFUxUgavxx+GwdiddQ8UQf
Bt5FdvxEegTqrdn1dEfGMvFc9/OblFhzmyt0o0+wAh+jTooaddAKAoyP0GH65rVo
VdG2Wj3akWLVNNlcKusZUYv0mgPAna+Y5In+8oB6ojsMOTUU9tBCvRlqj3BWrVil
WkWe1XCK+aI7Gj2ARhp0YLJxvwBzFRFyNgcA13LcVrbHN2sycmqPTWq7xswclzAo
Lr3/lc2qHtxdxZNkXbrCxyD7JGG9hXUM5Nlkk/IA5tHnNidCdmvH5cX0T0ef0TQO
0KA+cc5zeBfkfpi7GvJwXBCzo6Q6zzWW6/BkergFB7oRLXjw0VZPoGTEYr6mavwM
+jstHZbsmSn7f9akrA4IgHiGZFj/B21KPy8nFS0kicqNa9OSuRUsRHQEa8KK0V6L
oIitf7RbXO+ITae42cSRvMlm/Rt6/v0qY0/48gWKT3wK6bxHzrYhqM5cOJN9N4iV
O9ODNdpvBDwVsOVGhN9Ygk0i2vbVlihfpLymSOBOyF3vAhGF+5u6WC6iaxnuoKuZ
OwM1Xifo5CUkHEgRtrKW43VYUL7/HJTXJ2iskQ+3PX8EAdu8r9scMBjyycWTdnED
7OBvBPHL8cfRHmPZstDPhEHzgwSDi0bKggCBD4kw/1Wgy+tPsucwc4vBanJzeQIk
XzryU+4i+6LtI4jUjicwTsyHn7RhOMbeMuL9NXR/ZFk18ev5QJDCDZVSmS4VNqya
SMOpAB9HhNzijLXUD6EWTPHlPsIRn5/J/fp7OVr0Xt7lpp3iiYtTUJG8k62eLc9L
2GPTFRHs03MUlLUJT/KFDfi1siX3i+VNhO2xpJn+cqmqg4PSVw3RFjb8xckoFwyZ
vUjVR3UVKLuDwyLtXGj0j14e4FQ39zuqMX82zgOxb0bXvpAcA6cSLwZdSCRElQXa
XVeIEqAjafRQtfrRvrPAs3TktO8Re3u3dy8p1NwYg8Uk5oC5v3pLpNrnHMQuM4D9
8QpXSfOWcV1yMOnFIlI7cWS8tP4y9MR9EeQOKEcHOkefN8yf9ainZn0+tzqgsXRu
2iAtWjVjpyERvFhDss6hoaegl6R01bnFQ/qefSp2J5eOCi597elj/j3MRkj/SLlL
asOjYJJ/YDcZujPWdI5OKxCC0Am8Xir/pqeftH9b62NVdI7iEFSinbCmPwqEk07m
/X0o90zIpHAuEVNUccXnG3CQjHRNbLbj5gJAFAwvWFHypyD+ObM3CbtuiA89G2St
HNJ6dCL3zuZUGLZapHZOXt1E/E0aIUoSuh+8OYDtzS/z9AId1OXP1CM8lYpb3Cde
178JPdOd513yTGym43KRxaboqCC545RqAz4bC5l/YhBxLyV4/zqL3bnD7YpY0+dz
UIWG3JZnAA9KFLJJg6dysC9KW0bIN7quX0nmiqoHIpUUr5q71ZIvjKA84ZPnL3l+
NULtyxNtEAuz5G7ITSMpVJjap0qeCLgIa4zHUN32N5oboEbV3q914it2DgnoLQd6
fzj2pmax7UeItXffAE9m8gVpaaFJRC34Uf21IRB+mhv3ZGyjepQtip0x8FXRmvYb
LapilMKjLXgJ8pND29tevNja/+ezkiohiD4QIRUbBrHHa9PKTLHYoZY7faiOOQq4
M6s0Va+CcjB8ldrzlVu/i4n8pFi86Lo5pIuNLFDTG8J0mbpoFHmoqN4+dkdVNZGn
ae2O/B6ES0XqoOu5K+AshAuBVHVcpBuBVknFqCyDaLByRXURdWV/zKqD19FknSCm
DG442ScUWUKzp+kGsH3YZu7Z7T00AQYtlazlzomm83edZmAVpYtXO9FOne5dIIbs
CVMlKWb3xA5qROP5jM5Lv91jJGP2uOoVBHz80liK9fjrohyNi8TZz99PwoZKkUNu
nAGNue3JAHWcnpc7wWVEgjDQTzJ7ImEvJU2pAffcNC+yT6OvOR4GzfnvlE0MoLnm
lZ5A2nLuaZ7cd0PFHgOmnx6blJZGRG8x+J3Vy/5SXlLqsPV/xxfrvDUMqTyiVzjm
gj2xxs73rAym3v0gdCyFO/niwJ8TSctaFLoLUYJQmFsF5IQtGZBiksrmhUM7t/+W
iK7n8aS3lUgC/zFR5Cl3AbEvBiEKhkbua56R+rM+BWzEIKXJ9ENK1VQiHFKvVGKq
LNXGpU3XoV/5QgpVsZIQS7bxAOqd9RAnJ96mycuO9ZsU7pNPCrACZW1C1AxXO0Aq
bLxCh34x6u/WCZOUpj8tTAAENzG35Kt+4+GmdTP0ERowY1BNNdrt8ogFae3YZA1u
PxBbSdea701y/baDVJHBMUMOiBzGDF66OHAsLZ4WdGjm64mmjqt2vtWfEe8p9pPx
5jSpLUOEo0RSFJP0lzKiUW8EhtBIFTaPJoEVU3woBQZK0Bzfo9BTqka+aFU/OfOE
mapVXbv24vWQA5v3sZ7Lh8IZVNJVv3K4V6O384Mxdi4rohkFSlHgU6Oa6SVUBWzi
erL41Zj+fXaio2tTPTJCIoI8SuMKK5qz8ogNIx9e7PhrguHGpOnhOOu1kZl4Lng1
zP5wNInrMupaQf1KRRHELtJ+9LA16TgkJ0QP/ff2u6Ntf4OOzUoBp4QkEAomq3Qr
RYNldtW1o3KCKRDeDEJNQLJNyFcqKo23K2aa2Eba+d14j2SU9L3X6yAyzG4j5VYT
gCQW3+nFyliQRqqYqjwF8v3wBw4UV3aSvrSUckRE4VOGf5GHT3dITkBLQPCUSwnv
0ljW+WXvYbmdXQjrG9ig2cMh4+roZSkJ685sJtpNsbwdKLIZCnuOt8g825LMe/a9
UZO0l+vM51RwNQKIHdGF0IOhzvpwsPull4Yx1V8jc0R+1xw3aqj7vPBFiVsgd2OY
/p2awzVgCX6ri+gFSStCln5FNABQgIDikQtd0GWQ3CL45MJpxooBRkKjXm7VrAPE
pWIjB8N6I48MN3/Syh4FFgAa8AMZz3m/sTrmfCf9YLTLvN9audfObCyx5h7jF3jl
nIH0/urt23qwhbv1+Za3yxN8TQbNK41lxmBbA3TjxwINZ80BEv+1DO+7ZStPKwsM
QwcCECP8hhwJvZyOS+TKzKapmSTdStZOsxKy0ntzhTOCAQu4xquanc7Pe30CfoMR
3e0LRqe0CNasefLt7LDl6ctbxRwkJJZz7xJRusCLk5Q4cuCNtc055s4bQmsXj6mb
NLxJH6b12SKj3NaDL5WoglzbkZNCgii7AlYs7pEDiQy4IwHdFfFqV+eiiinxgEnq
sQZYC6WVO+o9hI6kpe84xRr2fykVaIDGMEzNE8xq1QgD0KBGLVSa7HhsbwNCb5o6
jqOumjWCr/eB0T952kop5xS0nrZ5mv5Hunp5tWRm+ip66dcYnL4WAvuPVV/7xOyw
uDsxplrxp7UQV3Olx9UOiMHnJCe5rxwTPIDpFORb8S8Aig58CZ8PFhgjREVnBHQb
pU9NjxJtTzNcn54+hllJ3ASZpDmk4Y54ko7ImH4oztDl8zDdNiDC2bu1QgstbAQ8
IUWF2Gh9SHjHpuVJl20cQ8y080iPUsnCoPPkaQVCLuI+o66qT4Y1lNznSlajlgES
Pn2IjRrE6L02pdviNxxUXnCLmfI6pM0ML6C5KvLNtM4yQUzTaJvPF7TLu82pBwdc
qX/pOOzuQ/VNPSVu/Ft9VCBxqg0MWlfa60kX0Yvsg2kCKJPiF003qaJToJ270obs
E6xF/t4oLb08K1SExE4+JFluaa9733waf41XbQ/Em6siNmqQ176sNYh2Je1y7OrS
Yab7AJG5g74vPB2dVktp7wO4IkZqx4DpERV5MDEZQPg7zFNVT8in7MXYUBDPdaXw
oQpQ3j/QYg3cqnn7xbX6OZTg1HfWASqw78ytOwnVoEFtTIwCj/vBgrrJSvOMJ/hz
wf1fHlhbDpsXAcsAhZTsTsfyAXvVmAEzFVybLjtDHYROOIzwHwTiuHhVaorO/oYK
FKfwLwyY5f5R2fpAj+K6yhoD+3TotAOG2t7hbISJ7ngZQL1/sulE8r6/TB2xQQeO
QtCbgSvUfhZbMwz7kCRzIfWaW78lmvVgAeKRgGqxP3+0O8QE09O9/IZvH/w7eSnH
a8xbKBZLpQf4E5uzmawLTV3icMZocjRHvB2v7+AMwviFDoSHTDhf3PJADT57iIdN
rjP226m7OsisSd5eHZF+WL3Hfzubs3JeI/SIpwzRfOfYv5wtgy//BmJzkNpWxuKl
ubTJPhOFqZiaYFDB/U48KC8lLPZkaQWsJ5qprBf0I2u4qHLrkjwqeo0LsXA2OV1s
H8sIUKVLzplHmwxtBXXtDgZjrlYkJy4X79+ImxEfXrMPr82f0KBjg2P4MwKRSedO
pVHRi2+r50ctUa0Cy3HCB5efc9uTbekkH7rgcuGy+GUO1KqQHaVi8EeKq3AJAbcI
LQF6bxst35OdIHyltgWovEOQvkny2iRtzu70mm9dvgG84Cz/G/v2QQbxaHWHrRNB
Cu0y8WlmMlARWvrscPHO0TOghY1TnOjZBh/RsKekAjLle90uDu2V4QxzL6NxIkv/
3OVrJi4UtyNQj5uoqZCSu7fnC4wC8t2jkxekxhrmuzWftXzHZampt8LHHFwDuar8
Gq4x2svXiCgZN6/vS1KZEx5eSCxPaGtkj8dwmmPW7zk5fE2lHs1lLDVfrOatFM0M
O4w+phSM8+TUyTXP7LEZs75Is0t74c1u8iqGKlcUvuaKsvrHyNyTyErDRGKaQ68F
9Xs/fhztEJe9PXuo81zOCBL3ETqzvGljrai6kurbnAXT1gsKDDA/nwiIbL2acAVs
wgZdhsZ5tiH4fFLtt2JDe9kfZkxDdLoP1aPA3THIBYcMwYGEr0cX9EwGwvhFpewE
Z+IH5wb6NMrZviVHpgT29hE/kO/7N/uZfGEyX0xnubrBGqIn9nwapUPy5TUcIwXN
mS+Ioqx4NFLzYQs522f7f2XplfTecBLGBXd9RqGJ/kEVTwLMxZDAHCzRTkXvbwg4
sBXfkx6fP+JrtUvUsdIUNt/r7UCnnh9cSl1ku5kv1TG5AtavV2JsKByh9h6eh2lT
CWCBsJHSus9sddVLM2plYg4qVSt24VfCDsVqFbdKupHQZ7eQgxUB4axFGVGdMhEf
4z4RNMSjmS+2V/UtzmOO7tPe/GeMo3wTSHd9YeqELi3no+AYX5NEihbAkPEghrvR
mYXO4BpI2QWHm+5u/QdU0z1VpgZjiBYsKMRToDF4rA+C/39WrPgk6kIax2h/Qfb1
975TkK3uMP4lD7d3z/eQW0QRwM2dK+dZwJUDXsyDgM/1r7UAwdZiCM2yhSY/nCj3
lIAU9w66SYuYPACTkOVPfA==
`protect end_protected