`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
LZdeNM1yImgoPyGqSPgENLiwrt/khFQO9lK0s0uGtO9g5e5ZG/HMsZ5x4gJuM3cY
ImteSp+tOnTl5rwIaX9EXyAMiJz3uOoWTxQy/0jWzEU2344uL6ZGK6dbVNl0b063
PSRdYbUXCbOuGofYga8kICe98jmIvbuO0T0bw7TEYYN+LJRqI8aMaJWnyg+/KO1Y
hyUTgtOeFF5OdqMDB2lcA7kW1P0sqlij6w0evAFbyvT32DeNAxza/oLTXMa9ZYnt
JiYDhFcuQ+Fw1UhRkS0QuWEjNvj51gd5AtU/1y1iq88BfpRJwIrnYen7/ayUUSEw
T5ORcFI+FTJK+CHJZBFwx+5xhB5qIjF4dtBiYG+NcZ8HmEd4YFRG0kCt/hDsELzh
3nav7mpp6/ktRHMoC6ywN0XfB2Yg5/KvaAFdQqqUN/aMNtC6Tqx09kALo7aKwm+V
KdE1A1cf6DStFh6Y3d1D43+Aa3/LPuZl/K7U6y93lxYi2xHYHBwW0uaHHhCBbtSp
+vFpcaQoUfjDld2zIM/AHZn5q8xvfvDR9ywJNJA2sdPVLYsVU/VCzeSvbfHdzn7l
V+LYBg709WOnqe6H13WujoajYPfC+OJ7gdYPYv+CBcY/bVR2AFMDVgyFDFp6SNoh
VvA1mBIN+4OV5shzqg9iyKYIVwo3CVvlpP7ZlKfzjZgIUn/VytMAxoJXz74xL1/y
aWiEOhzh5RYZA11kaXtPi4nE8cqN4msj1fIC0bHZZuebrDIQoHL9bI5eorIrzj1I
MtjXK0t2DZxS36Gkwvf+mPQfkTQfkyIMUbkFl1z5NXRGJ0VqrBN40fCgV/ycccPN
ALCGFvXsd62zcll6OcIYUlUgCvjcFXrUDKpjjWTv353YrLdjtAfzUPHmkhQSVf7L
T8eDu//vaTn3MxY4BbTOqHg25+cr0OeuG67t8TgNbMuTU/d5g8brHXaUTbQRxoEp
XcC2uALkAwwSh1dCYFHZGJy9aiJwhR9YNpknqykPiXWgft96xXCBCRSSNXpZQPDl
K6o+B1Hj1/QfHEf6kvHmBwACw8L8pAGZg75gJd9ZZyfD1yj5LpbxQiSzKOYtoxUH
rUMjvah68hEmPiUQGqMg3Z6NF6yV5BG9mZdEJn/m91iNwbgmjSnssG1oR1UdwkRe
fIRwP8wdRt2fQZnpvkApidgVwY5d0YSq2REsIGxOqKiGuRUkItt/yx40Jir+zEvx
7kSY+A1mGCq5j5tXq39PRZD3qPZSngDzBx8EMX+5Riq/2kAIDBd2xKp7c5Lq+bM7
evzWtsclPh5cm7KnGxBJDbQZhs0JUb9yp1r7i8eGzYOyTtVaMcGHFkJVCZa4tLCG
zaArX5tLFZMAMcykFOIaqqxgEoifubhGgvWx+GI1HL/Kj2IyQysUSTKlkhSFSIa9
Re19e62QUTf6oOSq9PjmNKhcvAzi+NdZCkKFTM6gzc39hHl4KYNNb1wLkvNP9Pyb
kJk3PHfodjBetvAp9iXn8Mif/yZ/2pvOGn9q90nxr8SspjOYKl9lq2epSzr61T8i
/SSpE5jjjC6mvZVSP7t0Orm+aGCkY06BNhCD1PlFI4r6wg/xSHk5hXRNJMn+maPS
81snh1xvmlPasXIsFgskiNTTA6X0orRqh8xoRn/xcEre2X6715JdpZ49sQ7z6tzI
NJ/+zZYbfhvz0IfY7dtXOo41PVB8vCgwDchwZpeH5BSJ0IfNTXVCbWntPrmBopbs
HnM2Ke0pqT7RbfkIAwE8lAIBvpx1yXmzs0GfYlDibKCqWn5+VuozfI6iZZraiOpS
EKIw1oCKjHZzxuZO5a6/UPLbVGIXjHPFCDBZiWv8q76mXfuAP9uowRhMLjdk3tD/
XnVMKdkCwUJlOMJXO8JG/uzQ8lNCrLqu5HkkfxnRhvhGcgzCVc0v0RUNVfIWiECU
/5GYekv2KiNOYZbrJOvMQWkiD/Mg9/h6N5v0fUiL5tzd69U3+iMrbo44wI4Ghv/C
elPQFm7ufxAGB2ghQhUwR0RVoIeq1C6hX8hNJZ8KTDsoIXvZ1DB3mcqVzVS1ocAa
jZKUIibcZ+EDJEda2Em62TTjd+TgZo3L3QJ0ySbWHxjDzThfhZ1cLymgwJDL/KRn
P6mSa3OqO3oWwotYa9aI4UyKqhRSZ61+YlN2wb6C4Ko=
`protect end_protected