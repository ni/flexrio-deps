`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzltuEBGe4K5uPEdMunCWo0hNpTx4o6dmVJO6BhlOuody
ezAs8INFZAQcpfQ0z/ir9uzpW3axe64gpDgIVh98F+K/wFFK/hsaWBe9/Dz94EE3
m1CJeVtIkYIuoSlK6P1hxcJHexGSSJlINnvxKToXKxD6IOOcw6ZlQyKgDtFsLOGS
qh2rhXyYbYgCKHD+MP5g9WFMEB+g1/gZIp4qiwVsn3bqRgMmUV9Ty4dGXNCavajw
PFnhl3t+Dd38Mll1EWfb8DgUoeBTp/zPMvWDBexEsIIKnS4S4PasYZxySEzeuNtO
9bcW94Ebz7T9s5brXgReh3YExIRN9X+ftfvtdyLaOFG0JB4E8a34FPSPdM4R8bzE
1MhsmiY0SVXsBHWNE0NCyLXGw19EsyIbI1hgfJyBdiTc46te9K5Tl+1Nz8uTNJTD
YsEP9QPVZT1aCfunQOLCQSjHRCJi7Z5m9+pkfvMbA3cwXG43nUh59ZctO/jBBGlx
iM9iyNcrV1iebuwcXwqTueDP7xZOUB8DenUn5ylHh6Lkq/eSD/txldX7T4SDp24w
FYvrife6OtbuwhY7NT2fiAO/76MjkO0XUtXp93LjFZ6CpMJMquZGpIYxm0lXqwPa
TT7MVSGGFJWJ3cgRez9JUaOeUo/eEphdZyfH/AsPTQTG1tAN2HbqFbS84olPf8Ca
6/tuSB64OKbVqpze4Fx/KyfKrWA4bI38AsK7IpWxqp30pjpM1gacQQR61LTxObsM
feUfFFCdfXsPTvRIIavdYV0kOA9nwM0u8pXd3Ulvdq3/GC9zMN053voSBWkMIMXd
MS9zmcFiZkgXw8fqlmpIio2YPi+tSzLyIyDosp0s4br+wlQVZnQ03pKJxH2Cv5Vy
UeE1jvhlPQOCKqPDitfmikcFZl96w2eK1l674bCto8voVcjEnDSlJOK5gRnJTatQ
TiL3DO/oCEtRtg/1lZ/XDDMILvy0A6q9qG9HnhVQiZAnAY+4SMXjRWoFng+VZw6a
0STOFE54etVJHV0l2VplQGFNKS2Jhe5JD3+15Umjz46mVtDoWXI+YdrxEurW8MAj
HzLziwdBoEVEc/MoCW+37DoVozccbxWzvvxfjtBb/EPcK38A/yEt3cFEGZNtuVtb
sJm0RMQAAQhEzLHuwoyYombDxm+fdZVtO+99l9P1mQS7u8fIa74gbM8PD7gUY0wQ
yftjkXdtS2S+zIOXARKEWIj88jhlgPwJtrn/BXAUSDpilbS6L6iRTZDvNbZwXY3b
mW+mFVpjCxZVi6mTmMGlJ3US+whbF6Hu+g5Bp9VOxTgmA87I2BYJDJDH8Z2x3+97
XHBITJHmTur8ON3qeZr7WccDye/71YAZNCz/v3jKDEVNyR0ugo4G8+etjnAOuYpO
CNsGwFnBnLNkPzzBfy0xeZvctNwDlUm/nFKGsRY1Ozrr4BgSeZ+nNdqvAz0Wi3dZ
HhIAXEiQ3gPoBAVpngY5dMJ3isSeFwk3LiVXZYaUmNSC42Icc3ONBdh5hFFe0XKr
FKOhFvJZGXJtBxrKEo3DMkXEEQLrII+GcBlCMW9NGOB/UUJYwK4MddLiRGFEqio/
reOgOCSRreEhxvYMmw0elnNYmE5320q3Kcn0BwaIUwu0djkO1w5yejRH3Z0m+QSZ
AaPlpdE0YQhDoLo7JWEM2FnVUZRmFX4DuQrP1buSyWQGSkSuggY0uPUtv/JWwgia
Ppg6rbVt2qviEURP6c21wHsHf/88bzrQZurzCBvprgTNxaNrmF/k+/SL1U3OlPUj
Yg4KzJKn/+aenHYf1orBlp4FcG2TccTAP6F4IvekRtPLoyPy8/Od1jrnxpqo1a4n
50FQGlfRyu+h+w9tFDlYYh7FyVmNtHvFXuvGxXJHC4/xxdH/+nlGukZqca4jN8wK
Xkatpp/JqCaqu4P51fqLYYi1iD6Gh0lLRkkrscXTuhenrUsSqfrsyZF6f+NaXioY
nxlhvs8B9pZxDIP7nDaZkSV0nTOfS4sV7tKD+b2WN/E425kIcWHyZNfj0M45Gjtr
JYrDcLy+yKdUHQ7h/tmHgm4WUPqrtE2ETwF0L4xukv934Cq2pd+eVtGzx5bCPVaB
vSd0LGfc3mA22QLGNNHdBy31VzU51aCNG8/K5q6XE8VGcyhqmiaScRexhKvVTYr9
/jW/GItwhTpgBZSMZadTKybCkPo4Go0AzulonehMTvxERN6MnuFnMeiGAAqvMP7v
AuCJQEUbLLp1KvIlrTHk+tiRZUo0qvfTqdl1nSkeyPhvtMNTEKQ+95upuYHqV5h/
NcI1gb8NEVMil35uDmKXtNpGkwjvPtI8iyCBMfUtqdFlhOLi12DoCYu8poSgi6VL
AkKueBafgBoc28eHJfb1GPGcr6yAF58kZK9SQJWN5tgzI5o82cWiUqJFMQBLop2w
3UvnHR+5fxdK+YfuRLFyYNc5G3Ej4bcArdd7G3G4lycjgTReWwumcVRkHC0JPpk+
UmTyVfeFng5X2JNHNzSgGdoOhcyVooM+TPKCQWI/+cFiT0q6PHQ4fIK6hWpyD/cI
rGtrmNfUXF/B8vm5m057wbERb4ErinswAWdjFRN5582yHGI2RYrjkC7hbdUoDNLw
yLCOYlLF8XN4TvWwHc+HSzlt6l3aDahCNOun8876fBN6tZSnx/ul0HmkTy29sT8l
PqSrjx60kEubecfu4BmpQvsXMxWDDvb/HX8Hda1Wz6oH02YPtYfSjNmZFQCODn4q
CMXgeZM3XT+tv/9IrL7haEj6AhqslzFnyyEljLguzeSF33rXMyZLiGsFtT9qRK+F
/eyXJh7GXK+7uvHGp5cpuZKde8Dl9wmX65uhc1FeOmregQVocxshS6zbLxVMy5fq
5Tt477plt8VjW7NfnYN2+DzuikDqael65y3s+4VGbPvxB4wQvfvU+lEcJVNN3NTo
OhOrI+Yd/QCP9/UJpALmFF4TDTRKBdXT/YFqsr/+H1BHU+TPFo8jH9Y4Jho4f7If
+FRIJstZRrCzMTLU3kVxXOyZbNjokFMQRakS3weEYIH5dUD+Pfx4C2m5Qt2Fl7a3
UUbwSZAINAlXahUJzvR+WOlztvHU9cB9cCuBXUDw5GtzRqBqsS8Xuqe+Xx20e1xp
oGlwLSVBTrd5R4xD4QdzCh/mRgRy81olGyDyW4OZsN1nY8jGYC7NHb9CUymrtn0J
JGNOf5IXEYCmOWrw00tx6SI7kfi9AtNTf0RpTepuFajThlUvERUVmZNna0blN/KP
zieJ5y/DX8Awvjh2QAAXzfnwTBImW78qIkzwZ1OkHIiiZ1eSCo3I8E2K8QVLVSBS
b/tSds0RawX82H2m9TZ+bgmd8+325nurWpD2QvfnNujmGqn+q3fVLDNudb9UKHPk
7owtVm+qqsoqzxmi4r2gkxZ+c9fjEqHEMcROdLiEzdaacH7Y+lwE9q2bTaWRPRFy
S0J5mrac0SKrmhdSUH9Qru4cVu/3/4Ti9thUhvMCO0rzXodLvoA5t9tKKWvIRjwE
YIAMOT8sQtEcm29heDDXhPSHuoIcGhpDEd6iAChGBnIyiA5sIYCzEZ791FUbLGFe
SEMsyn9KDLAYhC6H+M+DG6kKw1LpJ6Ig/rYS8nyKgf7av+A3Ld+GurlshT8WA0j0
53zF1rXz9CNjs/6zrl//IfdT5Vk/KlLhQqpMyYjjCdfxo0FtBS5iSWjruTpgVsIC
m44Q8Cu8p12u/l4xsV+BupiLZGz2dyInpcBUgemzbFMaWecElAhV+bZGMP6J+Zc/
LNqFVsj4pIxkdVQBFXd1GfvRAYkRyxLKuaFkfKCEsT7VqdVzEfWM3UkJM92SrMh/
7zBzkQrFUSH/bPX48j7HGxH5EACJ1QlVTyDFQYL4qQtE1i6fbjSO9PoPsOfJA9if
2D3kggrstU8xERAg/ZtO9Ub2AXRgj/TGJlwBRCk/U0HyE5hTWhzGWAkBui9Zlr0H
UmqFCO5i5KCbxkKraL3ev+FInOyxvI+1sCBFM29NDF1nA+F+q50AFEWVCU9y2Ugc
1uRvZzU/FCxErZMSEU77kXlqPHd7omsVxsyNKdHqdBRrlKzEuazOH7poAE70YP3x
anf4sZ5xga3hrC0MhuycyECPO1pmTLDhAgPmprrAOcYCWdxtdfFRWLajqYJIFZPU
utwizKXXFVMASv8pvE8QGKiQBR6ObgFYJ8Fq8cgqFOTa6BPOiQ2Q5CvlXxE9t4NX
cUD3gnWW/AndferqchW+e6yWy5uza9epZdlrAXow/9WPr3lWBptN8Y/VXMf26h41
zixPGP98hjR+MxremaRqr2AX5eDjKChYXcsKqiqP8mG6CtZTkmfV663Lsrv+PPfs
Lgl+IGTLeNv3WAuQXon+KjUbQZlco9mDEAPGeRFhi3qGgO6qxkvV+XIxFMYIMZnr
CxSBn0iLWV7VzUfDa8Y6UIK+wTGoe+d4Iv7IVOYlo8edjA1Mo01P0ncqB073+/dd
DCCwk+/5iMDXAemhoISHULeubpVB7A8NSwJKuC+GaZHptyj6bt5Pm80tJhEbBJhg
UpE8rlnMTBvvqu1JndCWdNBUNOmQuTSyR5j2Gv/O1c4xHi57XrbnheZfaQg3abgG
OlLrXUUlwgSqlyQObxZhiheRuHhHeywbGKaTHAR90yZJcLSkAqB7zqV1s2j23Fu9
DAGJE5CABzmf9SusH9TfWhITjdo8iZc7t4x3DbGD3XG92bCjFM52xKK1TkspHi5r
eGL5zm3aMAIe88zBUaCG/4ZovSDHmksKrwfMpYohIFPmaLLkuV/scrdPhFbo0PyO
i5s8rRbDg7MNAtViureRwR2gCvPAnhD+3SZ8/ImB+YHK9N4g8Pi+okNQKTgQjJT9
xp3tRd3QgbG63sMMyZt1TQmiavnSY45RoiNbWf0ClVpTRmQv3pCwKb/AVVEfcKKq
5hx7GzaFKxvZZOvRMPr91sKJeCDGP1nJk0sKgY1rt5ceyqT/5LfDuZJAxTJXyEEs
afkUDhJx79XarkaV+ua8cj5NUcYToVNzWLSnseLcdlnbpk4PJwhsjXDvYxsgFUrP
YLRNpLhleUjqCHvDOpAe9VpVsIV26QTAUULqk6oK9o4VFMuD4tiPs0rCjmqUUMLv
dTl4kkKwl+Ble6vmxhYA6aHXPVYEqgRH359cRejFz36F2F2wvsG7nzOnMxEbjVaW
+q7GjgZzNE7qoSKwTolLFhqo/17PqBFvMbqpy9s99MrorJyEjbWV6hB8AA34chit
qvlOL5L8lh9Xuzef8/z7twaxWfy9en59wdZqrWbs8pCdDmzlDJsrtd7gEyPpAlGs
qAClLdi1b39snADY67/HQf7A6JopsFqgsHwfQ9ZalpKYJZoFC1SwCdOW+IMLpywL
VyO+GVRnK2aiGIlVwDrCQiQMysZL/mOucjSBq2Y3cE0Ed6DZyjdj7pwcl+FbxqN7
WJ+zSoYi19pIPkBR4tgiv4Q45IsxcgLHfT6w9AgMG72bYqU71Bx/JQKc6Yesd4Ed
M1YFm+KvFvYDeTwIsBop9PVNX5FrHW6XzwXcqfHuO1UebfWF5q9DFG0+r12ckj3/
ECLyLVeQgmnCEGkpttohIsVUMBcotOAI/wabhSGnQ1734Vd+qDGtb63BfxDd8oNY
ZO5Tx7ur2G4+Kfs539qsGHxwN4mcyGxj/LA0NoYfPNOMCruVCYAr7J+jG+c4Ptzd
ZxFY+mno8pZG1RDi2A/qCdrWbrxjjtZ3e+Hav1HKaOvfxKiW3fojOaV2WYMslnb3
OLUuhSKhtXz1xNI9t8fxdK0bJMRwbYBRSO82Qz/b9rQAUzBLVd+tIysVkjjG6lRp
8s6slOhRv/DdokZFfomU+VOsjyuRZ97q6xT1LIiaRXgi1HuMtUNGhtlSsHfI18ni
APoJciIg7aSLsfyIZXfEI8GWcLvE283qfU3VmwPvslLR4DQtz3PIIX1ZJMSibRZb
6ZaGH9vIfhYTOY2qMKExc+i6VQ5+5iEvby2quuXgMPC7r/ONkwuEX2du3ofhwTOc
PTrZLSS4orbrTGZ0hH3J+EMxMFnl+lkoS9LuIUrjw2Y1KJViSm+BQxx5VjK1BBiQ
K+azkGcGVQZv2oLTT9gFqNyNkLFbe8EAwboefgeWT74tbGJNeS7NYRbR93CzRaxB
9kyK4kMys7wA1YGhfZp7Dbd1PSsigQbPp2Z+P+PbzWHDaNrjQnWmEUx/5tAI4c4g
nUaydEwDkkvLt0qTpKw3HSM5aPYDufKoixOikpNesTkrTmqhF3XL3Dms32cVPmgF
0Ewwe+jN+ZO2USiLt/VfIAtQJxB0HY/Bxyvy8ycPuITeZhXXWq1Uejs2/F4q1bQk
rgvrW6zmKFYPExUKlOVZe2qT95whzT3Fnr/6HsiWcC4xVXVQwjOiZwCXgdBukwuB
1GYUMJPzrAVZ/SS28ynz/E/0QeBj53ZUtIrVyN3cgZyfx9twmLxCWxuEZYKfVeDe
pIdugboXNGBbVxHAe91N5Efz+J81JY/z4gkaeXffoB8njhywSmJQrqesOI5aGVkH
S5w60/2fwcdV5hBODSIKznaRpnLXuvZ994aCpjw9HlPM/JKQ3/Frysl3HywEOx1p
kesZBcuV2sfbaGVHNQWSTuLDUrqidNNNyz7SHnLBhY7apmM4exzY7lNa+f9tmDqo
KrpU7d3Kd5UpvZzefdR3v+cLq2b99rUkYjZtnEMHGpX6qZO5E066S7xLiP3X17h7
yCxp7Vmkjg0j+wIfVRLDXzeNpeDGHKub9KV2xHCESLK5gFGMKvEyGoQQv7UANcak
dFPainngGXEp87/FJYrA8nhRb8cJurSyBn7to/oNUcXGT4kPRoGnjBfMCLEWZDoE
twgnQPsjodMICSDYk8S8f9vsmEtSAuohdChCBYYNjIt8vYVsXs86FimpbkuJY4Zi
FiN5YodzFv1btN/nNClVT5NqaQqfNKKJdb72oMektulqh35vLRhIJiOqF3M00Bdg
q2188ksUhrxLv5hLgG9308kI/jecgRQY78Od6Gf8Q34Tm1kQmccwnqn5BagyPypj
5vC58v+VEWiNfPiXZsLXK/KMbLs9Op4KOfzXN7ly74uYwWSZd3CMVCHbrZywjwRM
TMviT7NGFpNvGIcp9zp3RB3ks5uIALt4MdPKb+tsC2DuoueUntnnIM4L5YR8ZLuv
rzldi1E+3VIpwWcdaQpdtAExRW6PCDbB3mGHrceEpvBXtNiebm1ByhXaGXGyMA3S
yu9MSBRTjT3yNS/CLDldWHN9ZJYw0NhSU2U+T3Nd3AzETM60U2miNVRldKr/vdSx
8qrwnFX4nWXjLfOkRXHVzUdFh1cpD6fQf8GHG7Llcs1RzCkzdgBxi7W7VcCZPUPT
uyPQjmSr/aj5RLMiWNkk1I9Cw/xdVTA3jcIumX4tdT8SXYchJKC8safB8Wlzm++p
YB3+xVG41PLLHte1cvPqXuR3cv2rShq/tLYmTM5WYAPmxZb2aTb4gchdrzaR75UX
jQcbtEZ0TrYXQWs1Kt8iS4bSUk4VPuDwliPd6ehxQDd+BUAx8PCJd6hTnOLUVplO
0kuYgz6wtQSyamvT7kt0H6QUQpn83iZiv0Sp+LOmEdmmb5GenYJ8aj/zojSX25eL
qWBdXpF08Vy72HTGd3zxZ8ix2OobuvqlQcTYc/cECB2ysrKqPlew92eGqMqzM9Zb
F8mPMJQHZZ/WgaUApO/O2Yh8ToRHvybQ7TKMCeXktrhh02rBoTq33x/OIH6qhsR7
HM0FkcydBU5qDTleWthfNGjnlE6tjol/v+9/MuSgjSmLotLuE7WmRkufQW39GDW2
QsXbRvQalqzDsp+a3M8+as7z578WBo6fPghdaXPin9mwZwqtA215BVWezyUu0jnj
Xo8fFVrxbgaKnYeR+R+etawHhfEc8bSvER93EwPT2tVBlGhPGJQR3hVYBkybV34t
5UJ48W4JBXUUFOWuOVffvgO9uyaeXqeVIhEV8BZuajjoebpfm3wwkXdiJdhDZjPG
TNWp1f1mDicJNwHgVZwyXoBq2MiEjDu8BaS9RaTwYm13N0WwZrd8pCSNNa8mD/fQ
JgI06f7xD6e24o9JN6/nt0DVpCODgKyoaHu5jz2zEnup3hthTr0sUn5BLgSCjAsh
m0Pi6i2rdE6ohDk8xm0NGKBQDMPyg7N71t2SYdjCJY3DuTTRT2JO0a3NFZbudj/h
YIZpXN2kneNyx9rYoQjY13/xCQDo94RQQu3KWbNlbOzNiLgzpT0bbaKTyi3xsrJT
nXuFoo5jCCQxXFFnEB5PDL4FQu/fbwGp78rYtWWol5VzS2TEUIcPLzMG2hLvBXe4
VS4e1GH0SfinKUjdHFvomZO9AyKT2s2yoxr0jGeErb8c/hHM0vYE1h4/AEfdno9N
ayfqBdGOxcn7sJXewvzBzoiyJyjaox5rSgIuDn58GsES9pvYePvFqvRuN30syccW
DjisZsVipfeuV3tjTboI+IJIdZ1oJFTTv+ge8+MCxJofoMEAaxcC3GUJZ14ifa+1
nU/BH0dJwQqi2OyYZ3Rd9rPB0PQE/49k/I1bd+nXPZ7O7OUNkRWTEmPHciiNSnjY
FN3juB59H5u2vOQOT6CK1l8/uNl2aDUZP/AHxtcZi6CZxIigvtBNk/xp/4DSsvsb
aCfxuNWh+BwS7o9UaYrjhQh/FkqLGBXfyjvqt9sFylFw69/N8Pk5lZ4EROidOZPx
JE/QZqKxwKcgaU/w7ZzZiO2Wm0wD1h7rioFaZEbFYBzu6ETdHJoYUnFU2npUlsrg
cI3cx62S+XPqoVjRlcTJ7BB+ezWt4k2kk4H4JSGhF6UuwjvZ7Trkb3fa384Pg4LX
Uawki1eyzwSZ8S3Z+Fr6Mqtjag24YCHpKHewsoJU4MrlAKMZJjlQLcBwh36kwdpW
4jqkCtwOmaSSy0AF62zM2alKmKtBzQILoy9xufKT5mjaWSRuyRrH+qOx6UePizIJ
rRTKtrI7vMnfPVJIiiy78CYc5bFN1CGn7lVN8q7eL4gIJ1MLLF7417eH9NV1qp09
xrKt4aRrbXQO6Cx6EXimLkKsgZvreUBxOBO4nRBrnKsOnJqgnhmPBLDaEQbi71D1
aPjs+1LjCoO5p1rOEdQoxOs2Ifho8aDwBnErdLtQBlGMm6wdyYQ4JY/F0NZBWHd4
OSgZnkWmM0Wr7t3HexiGCgCGmhOSQmMx/Uxbx6RwqT2LwZaV8hk9PzSA+RsvXy3p
IXqynBKpWHqZIgbEaUdljHJEywJidV39Esw+KT3leYHxIMIVWHwHRz5C8uADvVdl
8t7UprXbusuLjZSBCWZsInsjSiDTwdQ7BUnOifyiMyMFwZg+MoRocQj+1ICGgMZQ
YXPP5c6pqD+CdwPazwO/aUhNyIW7JSEjN/pHZV3zzMyWB6/FedG5t1tWvJPGmplL
oIRGEpX3vCdp0BOAaFSJJq0EGCmPH2vgoa+CX61QqoXuPU1xAJonC49vStwEsdCG
wD3tBaM3kSOonhIqVsXFmVhNS8Cfd+xZiP/zApdBPVLvx1bO6nYIWKJJ0MiO/iI9
b95jm0zA9G0f+UmvqdKnyweG6XR3ugfyyK0nuxG3fW2HAdP9+UiXO5wetzjM2SAZ
GoniATBFcwyhlPqQ+dHxl3QVjKfl9ivG7CqPrTigxSCSZfr7QsfpseXuzn551fbf
LzGldjzc+Zx2/uyxH1PwkaYG4qjH7NG1GxYl9Q26wWE0yindOzjRNBw+yMuzPqFJ
moMWLDsCzX3p0xLOFDl1wEYyqtQnxYsWIPlb9z2dO17v/hDV3bd2mjrqasgyoWoW
C8f6tpibm9GNeLXW9I9riGA9oePaJdSoTk1Y/c7MJ88qwcgGRnmKLPQqP0pFXvpP
zffTyaur2ok1kNwVNWbbqlXtSPN9Mifw6yCDD+Yc4WTAHGEHsL/fsaE95dBU4+jf
YdHzTLlsMD3ISWREPk7iw4KrEBKZ7gc2jWruHJackU4LoN6rdpOCGz5tcQxLc/ar
VR1vCKWu1dNXBb5mHK0lgHPhYb8NEM7+FfF563tmWZsJ+WnmurhUncEdOfup3XC9
9PZiw9d1WMxTE2yuwCAQ6YScJBYVxyWTTIJY7pp1UdhxvWOgotRcwPQ2+MWED8oU
U5ClTB0HnL50SfPT+oydH0/sxyXv2bX8+9RDqyX8e83kl6LSGdWMZIDmJHYKYahR
OgYH6OZXBXX8XdnmJgpQoTL2gcTafvxgIuWSziFuZYNosESSKl10omkJhGGYdfRM
968hF46vEqT5lkpHclgNKYD6hWqqSDEAlwP1/Vs1Cv/WL6CnQ9iPxx7saovIIgSS
V95J3iOhILJBtPNMBeBg005jR5OPd0JWJe8pjOnqXVKoKNQkq1ZpW05xlm43zE5D
4l4LJT9Eg6dd7lNAbrci5Ka6q0mltvilKZoaKCzmLNERvsxvmoa8Fg48BcIxBoSJ
ZcthmryMEsRRacZr1s9ileR49frq/uhtMVomzXXTG2HavckRW1BgtZ2gl9+9Q4ls
NvTdleGgjqOjGLer5eQZ0ANO2qyMKIPCdIWa9ckCtp+caf/aWDp/HN2Dvfhp1B4D
G+tGTNtwPW5fZwN8guXgKCPEtatSC5hXe5seWqdJi6VCK2eiHRccKMaYLqkvVLpV
8okxKUKjC+xIIl0a0kRKb+NV5nLm6Dr37GEDh/Y+WNf6hVruRC9e6qxIN/LMsyHk
iiXg/RRN+7K1o7haJpMb/i7YllQ9VGyW2PUStERHKpH+iZ7xow+y+tMvtlUiFF3O
YifeJjXMj+44hOXRevXTz/yKbWFEkfuimyiKqrHkCQwj1wbOJQfrXwUvaSX+j/80
2UnWqXzzJCNuv+eYAMVyvJ62utU0hkSnluNf3oemZD11K1if9fZBgklYfqQ0RpmQ
DbBkmEz2eDQN37q6jc7UuHpz9JWnDNzyBteIhj7eeaVr3gY+veHGI4ud7HxL+7RW
W3cCNNOE33z6Wgx9xBmvE80yCgiVFh53xJP8ax2EHbynIq/6LyyvcwDYvIEiLoCV
EDEdjDzAVhrLZkrzvnHUFr8mkvexRBZz5CNAifdtv81V9Z8lEtUVyVbHoxhSpx79
ukj/O6q3KkRL+qP7Nsm8q0Kg5Pg4bE0ydhmvOF5PepBBGytnQMnG7yErGuGjCWpf
rbBn8F/GNe5bmkOrUVdKrvYHBw5uM3CeitPZ6fz5UXtcCAUWot+1mZ/eY5t7pbj8
`protect end_protected