`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemH0BOd9aNOKo6c/iV/1ruwDqbNRNdFIYNVh2sz5HB55L
+xHQP/0f8pnR/wHWfSnpnQTdDA1FLz2lXgsAn9glw7IGpfkxLEPa8Sbur8CBljnE
Kz2nA4fZMOBVkRVu+w5oFA5PYDxoGQnIv8y8Hwa9xYp5FcilMZ0Y0kha3YcRbhSu
EB6TK1txgd8Q+he5oEZmfHAb0O212vVXFRPBul7gtw23BkzpGINC1Uut2dNjZBRG
PYopONT+NFWjBmUBKHynNRVs5KY7cza1CZTTqOXWtug/v+sD62+kL4nBDt+t+w39
ZibzNsgmppPFiGb5PdJsCsODb+m6iJziUMSM3p1qIgqMhigKXxf7CdRlh5a96QRZ
FZWxxcqX14+zov1cR+Q6oJf1CFAvs9hXUGI4KbTTDcMzL9p4pwrXl+egIaHCkqqH
R32hC0U/+Sm8b1XeFqft63dg+hLxTTqB5vUTMFkP2VXD+oi3dKqd70kJVLuRS7H9
4mr361CAJvRrIxtoDHdMCuhaqEoOMTuZ4G9D7evW1is9PScxsMIR8qgQuhaFRObM
lHSJCjNYJk4oHUgLLoEDUTw4p08YaDsA31QpYhWOp4jsFYEy/xBYqQ908KPAQdry
7OEl2hoP6jP/dpaEojECRrnrWqSzEdEMwMcjhhwyAO70R1K6oaS1AkouME1NBiVH
KgXr1kSB944wxt68CyFPPXIoKTwAqEZ2tIRJhBPt2qOCl0aErrvAsuC7uTBuA84T
idJq3KLq2ptgN2ZgCzfXHl+d1rZHM0F/B30rku1okfwyVfOUx2CE9osWAqBgWpGf
LrpSKbodE0rTj6fKsGZg5nKoNz62WW+aHvUkhiUse+kWrzV8Cuq9s87Tlg+b3GjS
btFL2JQxqvBSKUvf0J9Bb/8VPkrHTC2NJ6pLkVgzjfUhAJAYsOlrYqW+O0GmGWqB
555ChrvVy5z+xcG5oWc58YjDNczVneVtJCIYOc/7Rb0tZeE7JPp3LbZWMWrHEp7T
Yt19vkimKFM7jfzhmt4TZFSkZRiuiQ1dqJTs0TlBxqDRdb+eoHonai1hO0SFBfsb
y0iMotBz0V31V53PLVnrNznYF/TzE21KE97yk45W6SBvG0z1IPL4rOz2CgCUWD+r
hbwxQhPPASEbtMWOntrGg5cz1YABS07iaIgSD7VXnq+GdzulAmW0YL6PnVfGNJ9G
zKkeqYNDsG/tBQuJ3uvFGAAjCnyg3M2IpvMfbqji1a9zsmW+slD+G0Cq8NntKJam
0FG+MyUyfcf8kbcjvSAXLC1m5kVEC5LsvinzFt3tReZyvjHqmSgKFuo3TQbhLGoX
/PggcuvMKJTwHJASTLKH0ZaSGzNhGJuDb3GlX5eXbO4pafzIPyHCK6+6M6FnC6Xd
yVtdjcbY3SwCorJZOr+ZkiimCFFFPBVz1KuMPhHdZlC+j1VCGS1T0OElelyRbhT6
a9N6V1faEYo/iJIXFxk5GWRRdGMpT9aAQpPS+Q+LwlK9WskguoG4Gj7ofc0g+NNT
Zi9BMHL9xFplYGU+NJ4qh1zWrYQfikgYOziCNTn4LnsXJ/OCJvXDb0ifR647P04T
2VfnSunpvvj/qBz04SJdBx2vtGr8rMNLNyRT+XBGt19c4FvERTojiwGpLIF38ARR
8SSTqSNaQfSYb98C5Ggl4DrqI0rFluX3QccbdNr50ZvNk4EwdVho552BT6KW34mK
JXh8lKVwZhfBlfvaYlKCos3dn6ik48JVXEy7wq8c/A+OZagSu14bEBd57xUL3AYd
q1TOzX275NrU/UOP7SuBfAAPwmpYOdSSaeqWVnDez9PRDPrKo7TNbm7cNKV516//
NeBJgAJZyGRgbnnAAwv0ZrF3BmHoi3KG40Eh9SP9EUH2rs507YVGFal98utstYil
60bgQ0RjXcszk3Bg1O0jq+Y5Xryb4P49FLsO7UJU3ii+/GvBon5VVlZQlEwYBw+T
n2Qgt4V4XTDHIkeCInSJ0wlNh8xfH4OrHjO5MmHJu4C/Gi/CBC1ZHI32+guteF2X
3RIOoK4JF54n2+D/5jLKeRXvRJt8GQnrPevcUCJ7WBstqyltECIkO17BuIAzN+Ox
7Yf4t//xYwsWr1qcBxtzE0FheKEDeVGyae6fo/4BJSwj6KH83bJUY2lTWu823z92
arbeEwuPPodzCJJ1s+rmrURT7hbnbbYY9YuhZLK/tuodfVb0x9CI8euLcUdJ/29/
54X+i/V9UQ29CpdXGOYWQqjyt12I0G7dz6ih3TxytQ+NsieoaLnSTxQrFq/bSTAu
pwElWGctCX6PmuCh+cwIR9C6Cb4FrKwzgswrrfxveTSyq1GnIq7bWyiRR0Vel2pt
O9V8+eU0cOy6LoUE49ku9LZnTiSYkkP1O8zQyjXJbZ+vv9y+2x4EcIliYpv0YP1n
twHKYF7A3Ick0mWO0XQ/tAJOCfR/EBc8LrrKhxr6/JysLEOOSwRRfix3XRv/pXuy
kltLpIOD7t3SJjQmfNJUPm/48ZE0tTf02GfKMBHhxS7y2jgin5IAzcQIkTXdYfpn
w2WT2ontmJrh8g2jXgULP/Y1G12tIsRLg1Qgmq/lvouURVBEmivIFcKJ1kY+qRPq
TWvkASCbODJwOB0sYrE+tTgIgdj4PR4iWUdyqeyEVtsd0l87uWCqEgsxWSr/pnyZ
owDEH/6blwhRXTeHKMo/9hJsbfDMbq/XpFwTSDiRiLrLjHYAn0z7VUxuGnVDh8p+
9tGcDiyWVGMlOHhrBZqSYy4C90TIGFG18tGaksLIL+ZY4yMPB/ijP66y7B/gU6s+
Wjj1YIzC+44VsSDFVMl5i/DxMY32Vk6cb1rRA84Fc0S1z5ZPhjtTUHtW6MjxxrJP
icX0IYvlK/Uohivo2NSxHZXRxhNQ23g4DwHn4AjCebIuwnnz7IlfZdbIzi7zg7zl
towrKFZPL5NgFBjPwC6EjHzKrghP9W9Qq72hPaBRzSQcG203Qe3lBI5mhDHYWWh+
469CjXE5b3rOov5qVF+pGWpBKTpQ9wvaLJKcyjZhzzJqqN76pJqUoiHOp9qoXUm3
gQNEdXdlDU2fl1PMuRCJ2xH45gQXhOr4ZO3CeI4HLjFIGi3cCgMJNCIVc+VKhOw5
EBdcPcZOcSVDuowPajUZiIfU0ahW5FMvJ5rp1k9ql9l9hG0RAWd/nCRyFSBn0ebx
xwgmEBp/N4x/NNdquddlkd62fjkZOGl3eSF71wvyvozXGxF8r7vh3tDGVsZP2UKG
UJILhyzuHMvTD/wg3YDUbDheA3vjlY9z7UiJoOYqfEvJm8OZFvfpye2jQ2byLQfC
ZUFAv7kE6PJco7Pk0icPac98Cv9rTdiL4t6kA4tcX8+8VXHOe2dxo8TQzDzrbeSN
ZJOzajKeLivsx2WkD/erDn5sbUP/Joji8lORx81Hkf9TAef86vwb+7vvm2AWovCA
tFBtLGsZaCmUYUc9KyaLjsltVwRj7tvVjGVuveidoEk0DKQvyYu2OmGphbpNJmW8
RfZ5j3sAa5uVwO15ana0Vbpu2VAfrXgB3Ca3ZjRMfHPVhEEbMjHZNOR8YkffgmNo
/UPs5JeoypdeGzu0IBcp0YMsMUOJlS0Hoo8fFVRgB1+g93tfZAImYPPtMg1eMcOX
3ldZug7ADTghbKLrDJqyrpoy2QzMnwnCf/U8COtygD63E6A7am4UGkuLY8CQcNUk
liTP/sK2SdtMmPrlCLLaDiumanPRGSQI5zpZuhyJLXJ/T51HH9aSKRCZfFJ9QpXD
j9bQBvcAITvqvgbyQcL4FfkXH/9IaiM4rAgqOqEDWVFQ2wNVUzsDJ+lR5J2RGXmj
fSxb0lC6xu5l26+f5Q8y+RgYUge6OLAvC3sFBWvMSfrmIs0aNwcDu82LHacwETGi
IGwUgl1aLIctreWanLOhCu9Ne+4YMyVjC1MclRvgFk49iYS/rMXdwkXfoYGoiL6u
3DpJzh3REJmY2F8pVdTjzjlySaUj5hjwvJSPjSp/oy3poZgmHT0tVeqpGaHAV895
sC4AgeE5KlnwUtEKc3BVe+1GbUoTCDvvdU/Jojr58Oc5v2V+SJG7REDPbxCrQPrW
Yuh3Mshz8ay/xoVo1QQ6PtTg0jHpaU4A9XVES6XF6+xZZSbrOQouZVcRcGUeoijf
0ROKRdF8qyT1YuYRUDMLIiMe4Mr8v4T4Fczca7iF3il8nu95Dz080w6H7HaffwIg
PR2aq1/Dg1ektaVsuSe3HNM/m/CfnfqET8MTvtZj46TYJsIozN2YMSQoYb617lHC
Mk/5LV7ojE/6rFP+X7GI7ywiR/QZUaTKwXObm646gK4lH8N+xhOwanDo605i5iXP
4ODBLww0fgHdcvEIxckYZpWlq5nR1gF386+AdyGUaZZkZAgnQxoQYq1jAPEpM5DH
hVodGPT/57KbTGKbP29ITSoOVjrPwHNn9/GOcwB8t9Px8VXnf5BylZ5Z8vh5eic8
OeS7Www6HL4eAk0UJJbouW1gqw6Xh0GgrEoW24j9ev8wQzt2xwj+saJddQ9WkxoP
qXf904dvMRq1iPBewO62nQLkZoAvhmp0he+rA0nwhKnwgvGevjtS/54ehc5npgNB
B65oVsLKFjt9cIwPPp+uoIjiaQ3TD7dLilIBDFqu42mma4Cog07HpY+wOUnnSPqV
EpuE8S4mvmyCedmVqFq9Y9tHapDHDMRVbSz6/7DW94tNAB273U3ppp5lP8Z0tnOg
aN6hXzYheB2Dj43Rzl09giGMx4P5UBdmocg+lNzdRAHuuHlWWjgooPBvUdsAfdMn
3uBu1X1xYI6WD2uY2CiSarjGmuU4cIgL5tfvZeqrAHci56HfWJ1junekIY/Luly4
O8aTLffs+5nZ2g16sYB+HuvB77YSyf3OFmQUeVLurMDUbhRn8z1rtz+OazWef7jA
iazmrX6fKXb/6CSqdU7eH/A8VN/dkQ18LKCZfrUjR1G9Zxfik6Nvh4+oiLwzkhLI
xsVVCp9TP8ym6fn7pYpcKuCaJg0rh+KaINeBsPid0Q3Ql1NnN75jF4RqnzF4lVPi
4WuBVun1vZ06oHAx0gAPIrjhhOb+2Mth6Kq+YDm27y0foinSEas2tRIKtlTTIYxb
PlrKzfOqBnQb2e/j6IRMOAhisnVbAEvp3Lr6j91KbMyWj7B93xxP1h5rn7yeJZMU
2frYHX8s8GgDM6QJXGhJGjnCCfgakFMMd40roaKY0nzrwJNCXJIAYRPPIVJYmBKH
hsog9Ez1tie0PrrsVWRrWKKZt1PsyC6yWACTz1DxB8lO13JKkp3GnHEeLyzBQyU4
0k9wjd/uF9+TvsPkyRXWown6I8q50aMgdXqJoh2To5xR3FIzI8fSxqCkQgfQMSXq
rrmRUqepiQkYedtqIcaF4siFYk/seKWtsPBnVNn+nQ682Gxk0LZ6PZGaRd+BDtcm
Mls2f8XMkUS1iOW4PX9wJcV6V4g12nRB2hktceUbAnRi+l6fpZVG745mqDF8dbYW
IFbcn9H1/Mlsz3i3KHuHa0QWMpjds6EXLtjA2Jd6kzDLu01zhJXbzppCwWege1ad
5So6Gwf2iGXqviP2vT1aY5/tVAMeCLlpk9elMV3/9/D0BUURecZ76S8L90ExEUtf
MP2qkIjnlGgEHmfe5PW1w7CdEXnVDM+mocNjKmc05RwIHUAMdx3LWcslDrQSvu8x
`protect end_protected