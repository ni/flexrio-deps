`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1adJXUyNzEKX18xw111ld7mUZWMUdPGS39zmQM7G1RKq0
22ZVOx6Hx2AxnYRsAMu01eiqz7k/94ewuafYUyTU6lZ52yaqwf/Vn1DVp5H/+2vf
4baviWfDyB9l65lbR7tyR97+iEQzsJb0FRMZniU8pd3zkxKYApigrnf6K9Z0jOOV
uRNm7ePQOrcvofGZG7pXR5tiiFDMgdoBUTU7Kh7BDnCJKprza8bLBTzFCtzWxa7v
nWZi3ZMJah9bk0zUgA+umkI44zPG/rAZtcM0gE1H2LjpPtNx7e5nqGOODxphbEK0
Qo9oi69yf677ccU3l8AvvnynVrj77tXGlLvgo85IZgabMfTAqdczkHcE/aW7Gvgf
Fz0/KY17F/f+JIAQPRI7dNy51fpmJOMcZRIx4TfgwAR8ROhsJWoOBPsXrY/I/drw
fIyoEgys+h+DeFWGYqBzqogBcA7kQje0KeesGi6H3FLayo32tQ4y1JHe34aWZBvP
uF8XTXTQWrQSPFUB71wMVbAjvMElV4ROWFjuJrGFq8jOyf8ClbX3UEuUaUN3Z134
2Uqu8RGGMrKwve4TAiHR0CzfTPkMuqe7WMdeRiUMuBPNkLwAac5/26PRI8hKBhzz
Nr1aIc+dTZYVVixlaUd/5oNsWeombytfk31gTlcXj6I5e1vYJFUNc+ufMYkJA8g6
3kHpp46UjHG6fGVSlZLNVP/pZrDEI+HmACigJeOlITAp/UWwXgkE/sknFLUdoUwR
r+gnE0rqWbgsL1BN45mDsNaawJ5yprifenvRzWCPjlYI2TGujea6i0oUETIUONWm
P6MJmR7uO+pxrL5elPgt3CWlV5evT/GvR57LQiXHRERYWc+/0sXnovn4hMcg5pU7
Y37cg0gQxXDf9k/cq5x/jpKz47JINw551aYF3rbCo8cVMnQjqqfk5HjJ3/YuCUp9
5sl62tu9kT5J9BQKHqzCktHsE/gaXX+QdijHssbhkeeLvPfX9reLE+IGm/xfpvcR
JYgZEpGoT4kxOpLZcErdZi8iwqOtq7yX84t/tApGdQ/u7bRDMNdIwP4k6oF+DhuM
vXX0drDhR1EjrFn+xiY/TcEvfegExTao/s3KUFIySRLMlR1U4fZ63XBsLuaHu7uw
EGMdo2sKB3Rx6ks07IXP1/hRskw+zUglSjJpFj9DkcAvUIQLjPjwhbEL1Oiclh4a
kAYhuZCt0UaY1lZTEY0GQEO5oLJ4DcR7E23Fx8rkHqQq3s507XgpZBk8rqW5avDz
MJxsxjPW0QH90gZxYBQFcmU2ifOACSVJ6you9weRQDEvmrn1fM7NPW9RP1UM1/3g
X25op1HH10K/RpiRYG1/J6CML4L9HNmIUUEPaF0jnLwGb0RojpvWRg1WHpGzW7I8
1Xgw6Esa9SiEzhtyzfMNDBsbPnfPTpoH2aYVajRTOsUzT/rDeBX7eXdiWosaZ7Up
MSfXcJIAxGp00CX1wzNIaYSD0e5chvx7B5EHbPdm+kdHYsyvpajyrwLoPHhCs8GV
mc6KfgSjibcq+0Y1K6Ry1UeRZpbxE96x0U9LdHjCop4yfIE/ho9Sy6i3inidIE0Y
j+4cbe5+ajckKgLqkVGAQnrGTK1J8Y0+GlSmk/Zm8d2R93l8kkufclQjdLKq/Hy/
g6oryf34i2c9QTuI0XhWsG128am8TwQvjIfYOAGASst+QnQjij/+mNYkfiW8o5kO
Rot25U5O0DjIHSGN/IMGhzjeTbHd7v2BdWRzbu5n7o77freoGHgeQSreFoJQonUi
6mQQ85S1rQLGIV9887lJ3HAi+YaWROkYTLXK/ZebEHG0sVcpuLCUMJ9mfn5xQYRN
/jAEUB72eDj3YQDC0kWWQe76ker7ePVZ1+oVPIQMjI+rVwURuOt9tCWwuxG/h97h
j9HatkbQtwl13H8lYMLzfrc1Ieo/pdwRXMaAYtTkFTeexZwt9dOua1eWuATrla6I
+zsE52sxQi7C5d1tc2H8WarhVUqkat5EIV1b+w1KKjuOX6tzKx5hze31HqqkQErU
VqHR3MJNa1bBmHVKOqpLs0EUFy8ZNKflbES+BHLS9gXby89PFlaUGwRb0tAAs7pa
zUUW9jY57cpUTGBKzU/ahdDzyFTyn19HmlOSWrt1SCBhiIa7WZpqwmA7D2fIiQkG
CZDWeP/SdVntBQZ11NpHuLGGUSVBUbn9nMHWEhJrnaC3nuHslyHaQ20G8oAU0abx
/q+EExXVAcRnHFKo/oLa6KPRue+xKdEYI9AzVbdMo3/B02uzNcIwIb0n7VtvSPKI
4IoJtjdD134kArzpEt2eX4tmPv/NcaMsmH6LieENYEJL3V29etsiXWYsnzCBLeTR
DJ68ZRwdbqb8J4mBEvs6DH4qw8LEBlAqK4wx30D/KnljOJQ2UYPTX4cxBpG+D6C1
b2FWo/rqO5f+8z515/P4MR/kS3WXSjhT5suzlYJei1oaDPUWHClOPD43ywdNX1gh
XlCxMQDA70lnTXa+G28hdV/fw9vCWyIwD4e3RCub+8jby/6o/csQrHwR0jSz4wg7
d9wAOCYwbFy/03O3wJlM0/tfW+YrLQfO1VUqoycnjY7nI8ZgccrZzzruJuf7gnSW
hIMgXLRQE9NXMjsfUIVGMSf/UVxeyWWJECeEkD1hyG6JfRRUXnusHUKscnugOu+N
OlghPPjCH8OoAu8opWpyMNlA/OpYZv5E3xa1EovlQASut5UOf7sIpSZF3VzkSEWr
vaIP8dA34Pdy25o55xXM2TCukLXUOTKNm1BdryFNx1Tqs/YiJxNoS9Vek5D3b0Sg
4KpKiNAg7kLGEaEQ//rKq1EfyM+J71OgKqnXgRFg0tsUtnpmnAMbJq4GrrPPqyUR
PONfNBQUETJkPzcxFGUGOcr7I/9cDNTl5cfkihlLp8q8yhBVcNmSkGaZJgqlG8cA
dGy5hjLv+vyByaMbAR3M8fajcQnPbOoCijURiQ6dt7gLch9SdSiSzizbPOWCxDF9
WmIkg6hlQG3yfe94wWYC9Sb/qh1cZMhPZ5pToqO/KDRVFRgCbC5B4unL3zkNm/pg
ENIpuEX9xtUvcQX8EI/ODMrHMWmIX6dPChrnBmOilb/6T5+u+49AWueXBvPxAXJw
AiDot/u+p8jhpfZBY4HVLBihaHznNROq5P9OUpgX/44J4mFqXGiz2uwBC4VNH65a
k994LNCQhqQ8ZNtCPdrjwRc4asl7AL/wpWNH9I6NCOQRxpzDEtklSffDXxqC+UQJ
ONsaowF7Lg00oN3vNU8Ic0iEDTYgK26FpY4UcH9/hwMzE8lEqCJz9N7193Z+iKvw
J8vc5fUSK/LBlShIhqSCr0+I71tD+5lSNjQlM4nHoRkaO7rGIy0TKOGkPMuNRG4c
uGVoti86B0zM2bH7sa3qauypRbXMP09mm+g23f+DKGYQ5auft/JkXxnE6kliKoon
OnkMm87Gp9AKQOGcPLwPw2VvbILIlsRiEhYUO78hFSHsZTUmaqSO2CKfaEwNxJhP
SEKewu8j5/MSIII/13YPvXfZuOj7+X70F3GWzPb1AWvyQL/if7kfaCZYQs1FHctt
RKzVyrhO9IbeAc2VXdGO5gq1r7NBx3UgyGvskSRyJjppHOtACQ6w8ULtO6LqbDuJ
ZsAaKUDl2TNID2BIQftXzMgjFoE0We3L17xHfDC452I5z57xdO21VAGTPJ2wuCsA
C+INOf7hwE6Ab8E7SGEctnCd4LomOjpnw/g8EuvKNdfUm4mbzkG9O/FLti9Krzrp
M4CtUQQiGDuQeN0M3Isz7s76sYzZACq8T3ZsqIT1pmzrUIzxhPg+ClFq3CRlmq0U
SBVSMISeP+VshH65pdf0w2sDu+DKlslX4e/LQxfHbJ7v+XsJSDy+wtQOszveRbQ8
Rg+IgmGomPqdY3jjAatEa4zxzxyyW5nseiiHLDTQ2WZ/mxOP/trw64+mePZIxN6F
egeWGi8fCjgCIYZ5B36NIBs0W8lp03aQJlYUf79bC9sEQpF6qBHrbMbPrAQUauWL
+dNy+7R4+TJsiTHBQJFjkSvqknhn36QGlAUrY2JwDSX+8yaoHaJ7vaZl5jDXthIh
fGZbgmPt4eBbPjf029vVwjxwuu+zolznhgG/9EKp5JaBVfP9jHyiN5DAq3fbcsw4
cfWWv+WbAtfCs1/5UZvK3rMRMtz71i0ZA8kP7KAusgJ0pKdoQuaHbcSv+21e7dgd
wB8h7hlRh80rKxFw4XvcUWt3VEDUOPXxWwYcUR/ss2+oyaHYx58VsBF679Y45m88
IKz2bAY+sTmlDRMKOGbjMBb0DqgB5JegOQptJoZM2WzCVMiq2y5wl9CyHvY7t+hz
Qz6IA1EuhKOlFb6huXTjEp7dYXJD9DwIX2rEB5LJtT7pMmu7RHcIqtYPGLFMtOJE
mEWm3YEAiFhCSNvq7wsmdmhIJTb2rFnAGT2Vr3C++poA33/xb/Saa56jkdQlb5Fx
nZonWjE4f4RMoLPptnWswRrfp7nAAbjv7lZp+2JPu+R3ah/+zKpKWJkYlKCOoTOy
Oc/3MwGrov1JOPJKFwMB+rmSX+wEj7aqvn3ztJ+bB8JnMMfqRjDPNZjSBpiSb4U3
bi4T2BstDDAXlxiTmLDO2fqfu8yB1unUG97PKaryJ+uFfFhupoJRDs4a+1j/umGK
SARU6oOc94KcBH7uOc/8nECpA9p2xbecr90M68HmcTitkIVeUT+vZEwoHvaF6UbC
Z4NZ4VCAmQ041bWxSB8tW/h6n7hKEM+8msts59nSv9ZJgNzwKsuVMJT68wVwbGM1
KXNTN+zacbhL2RYqLIz5sgeK30Oaej3whI2ecKfcYTHDbauNiBhzfCTVjAxNMHFx
SXgFBGaygtTpZfeILtaPFMfXkM9iVnhCLyPc8LD5nk775z6SYVAKIwffW6IWAYR0
iDMbmvADuPVBfuAsig07MKYnxwoVD3k21EbgvpAdMowZUqrkGNSQ8lhJicTicIkL
AqefPNtPSA2SNVf/JNQeD3yDdziXuvczDPm7gmVFAiSlg07gpJhSHU/TZbfSviIr
4rkjBfc3Pk/X9cWcD0UuAhzLdHp7O0GmtFQJjfybXMa8d9hqcTRM15T+7GUcfsNV
6d6JlesGo0HE2fi3XF3yx5PHg9sXsFAfquL5YaTsg4b+lrSaVuuAMf2E0ajNGxeT
GW20ZSPjor5Iv2cJXLU4eNrjlvM7h4QkmAObApfcMKnKh6z/rmUe8R2H4Stdh5Kv
BUglFneeQl7Z4c4TcSK5qAaC3uBtG/E2ZjZF0wjTNqAi0USctZnumG8qdXgEXm60
M3tFvX+BmGxYNueorUwHYBvCy4lIQJKuNx4xhpj0iy6rDnNVkwVrB1Ni3kPZn21w
DB6vodDVrSVBHMaaXMUGa2DAFtPMvDe37xP6I2on8cwgfmZGEqYhd9Hv7DAMju6B
9/AZC+enyjBvsJa0AaI4sfi9rup6HE29Y6W1yFWhbe9375FGhbrakVKCLhA5LGF1
1djdCB+Y4BGcXGcODowzheLC5kRR5+NiHAcufCRdZp5AMRDtKRzTqxYKQ5PHbZha
6bzIAXoVsxFV6j2Pj5OvHV++ZRQrJV0EGaiTCgxKiFBQ9DJ1smBEdmuUkviZ6hvH
5CUSYLvxal+Yw9VNgDY0nd2d5gL6dH9y8ju74F2pJYh4Axn9JrIaxyLs7Bg/wWD9
iUI7+YeLFYATqJD5hhUo2uoDDHiUU7zOJHTfJueh37DbIx+IGYqzTtrEnKoAB2Gj
G/2OzxkjvqXOCMVpLlFkNaKBFec4wXcZf9m9zWzYw++6rDFjzHPjbmqbBnf0JLCj
U24uK8JvFIlxRkhXinWU/omcsZk7mCSZycF2c+oOms8MJxACfzEC/Ewqdy+OxXzQ
bkqqb8veAovh4sBglUI8Se+smcqMvinV/9XHsJzogNLX5yR+cgCXZWh7YuSHuRHd
nVvzakTk5HjBDTMmJ52wpVrQRQ80TTL3U7vob0b9NAfEgrNXVlRZt8fW6BAcGEuH
uWUd63FCjwqpjGWcUsIVGUhPGpwFsdQBqebmamR3LBo5d1Ef+6sklSQkIyoFvkHn
z87fEYo+LSgpfytYaozE5Ktab7/sLZ5yeRiEX2R8Jzlv68bm6Ja+Wa68bwv9iu9S
/v5QzmF80vLhHBRUH80wijIctkBAejQScS/J6ENUhyytJahyKIIbA9Uw1/bMwSBM
6SILK7Pya5GwQdhTbZMXg2MpeHpA96/b1gS9MmKfy2qidLdJ0dRgGS69Pg4ZfiW2
266GnJb8nOK/gMR1a9ePd4wEKYVW7kE9byVMcz3p5jiXb3xfdajUTFOY8BvloGFO
cc/47zQEsFskQ3XMIOCY5wS6Wo3f2SUzU7db4zsQ/J/a/kktH/DNkUXHpv6ejhY+
Qy9hZV86hskyTVz/uytlCGBVuR/wHlY6PGctkHRnxuPciErCKsFRufdmJ/sRmPR/
cAF+FkJCNQV7y2szZ5qlxNj0eFRLDnVETBfRdKlwYCGEPS25vr6PJHjHdjxllxDI
C+d2rbywbeZnjxnP/vA7XL74vgJulAZwAwUiwvTZ2TcJPkZInOHN2UqJ9GmLmunk
QfCYvdTO/gZlKI4zkCDpWhb9fGA+nU4faGq2BYwbNiANHGzOIT2RFEDdxwZP8jhA
+7Q0rgPHP57cLIimGg0L192QEBCRXzTP9k3u9NZ8SU/+55deZGLuZYVg+MxInHXV
qCz56l8n42p1Ot26d/A3Dp3tC9lyTp/ip4SFuheV3VqXb+YiuFNPb5XmGyzbKMmQ
MksDRMbrEF43GnUaVtfz4ML54hI+f7g5AsQFHRTs+vcl0j0G4oPPC5JUkT/8RGLd
qub9Q6M/kVOxqmh5TwDY0oNICmoXFFHBA6ZQbGNKGijzw8yIUqqE3m6C75FpcG1s
CzCCczNMS/vHGN4dYneOlDyfcKG8I+9piZWvs+1g4KxFrRDjpPcOPE1UskXU7Ahz
X1r7j99ebXiJBs70lajVnvZ2/KAB3S4qQAw2RC9+n4CP2izaNKhAA3jL3PG3CeUB
US8yr2uYqCkiDTYeRGgSg7LtD69dCgnfyHj4IisXyr8pNVXb37U5gfhc4tvP5ELo
fYKxL3zz667huGUXukFxFlm+t5bFyt1gZlc6jqptZg7rQfDSUUgmvQ8N8hisPriz
7i4l0dfGGwEuhDsFoT1g9DRD+xnSOXKK1ee+xC2HVHcDbod8q9JKuVtHe8gq0F76
IHabWRAUeDjmbDL1R7nWl2oTe6YUka5SyBW1S4sMrBueQ4YeYg2iGt6lxCIn4cSV
hO1eQl3y+2qyWwt/qwLl+hjySdQHBdA7rEiWmzVc3J1F9cV/ol4QA/g1w2zY8uls
YiaE+j9F8iLWHkih91ij7bhLMK8rWaXukWfkWUnnbYTNSefpETGiYGgQWnZfAlH5
1ijxKnSRDkT7CA2KNOZhKbWp+I899h6r/TVyWNzFxzOJqkccxTkj44WcoOpeG1/J
+gI3TCFhhIXhDk8laWNEG3wTY9KFo1kQWQ62kAyKh+Mp0AxX58ZjXg8ay5gdqUKd
CrNxVjbcMZBifR0tqLd8exulkdI1bwjo2FKdgFpCKwELl0P9OEmAC4XVUirMYO3a
bXiDDytDWKqVqpB+tQzo3CLmUVRvxUOi+a0h5RdShY0Fk89ZTVuhBNz8CTRV3vSC
jvd29as2Gw3feFXOY2RCRWIJw2L/FF7nbyX1BvlPY6uBbVNUuGWG8lcRsdzSxt0u
QbRnhevS5Xhbkh+eHI94K4lCl1nAbrkXmTk9QCZlGjwNdzzskZ4w5PmyraeAcnY4
Dg1O93yVNb8JFwzZVEmBpgCBADKrZnfhzSKBffGJHGWmMUkRz9eRrril7dWgdR8O
+6wzYglSk7xGfV7f7ZObM/hzzWuNSOmzXLDTLwF/WQimclQLePMOBu25Cb6Kwve0
R10POlATHKNaxnXL7sO9rR1Jw5HWkCYT7sAC5lSsaxpEdjjYK6M9zR8mxAsiW0V8
a+0CeU0OeoTeQDODENCnnLFwVAN+US0QFVxK61PCSPe3JSkZ9zLLgzfRFUdkJTfj
zdDIXVbCK63/MN0kp9DGz0nGJsDiK6skwsjyHw9LD4HySDAAYHb7uKV+ioEbuRow
L2rFNtL5SbDTzLh8K7iSmwdwK/aF8w8NShTKIdX9mVMTL6FzyLaRXMp6zUe7FCTx
A/q702OoRUFPD1xl7oyJ0BHp7iujVOB4XjVPv84KVVce3Io8LiAJOtp93A7X41Kr
u+P0WxBlhiuGny+mKdV/G2JBLu4DqLJNpgwNjpjPn0cOCpmlglYxTnpk9WamZXSA
+aVRWg+bexnRvVlhtDPLtFkqGNd8yobFITEqI+eoPPBJs0nKghKlVFNLNwr52Jdq
TxGXpotk81PMusqW8oVMfi8HTIvmtVMJ0PhxCblB0wxBdPer2ynghd4CzPkZnTMz
+a7I5s4YyeKa9f3Rz7m5FAaaVJCOpoUulhdiwVGEL2c0secI5Ky/X4ny5q3X++4S
nbmrRqsTzpRGi+5KR0DMTZlgHRvJh/mPyoNp8xJVzOKL841weUYlGBRjWTBs9Ylq
x5eNxLvCRDb1OiHFMsT1c9AAb3/8yrA5DXkLM2C1fyjDc8lqJRyaFAF9YPlY0fMQ
P0EkZNzEG3e1+Q5bblKLQ77m2fStcGs/Zj90V0gYShM7XclNIu/nCVrbKmZ50bO/
aZYGm2Wf3SP+XX5CMvVhMdPaVFSIX14VyFI2byiOf684j8GflTeD9mnBCdyQduwi
ghcacFNT/EM/7WixmYYf5khIFYMPs7BYuim0KT+3X4dLNXUhSjd8UkKqk39/ZjSu
PNoZk6mOpYNpJB4HUZMNY3+wg0XVaqGHATyuBpO7BJdp+GvCktel0/gaRA3yeMFe
Pj6B+ndXzrEKdjuhUv+o9e4ygvJhX+gh1ZupRKpWIJYvpZvEVwO7/fUpkt+Emswn
yAfWFLaSeQ23DZCBpruBNXv74O8MOO/bY+blx7VorUg0f2tW67EZQOY+WF7kfHzi
MziTdbT4zuY61cJLi82uzzLAPr+JxmYf/ol67M+92yplzi9pbk4BrZbDj/09QBvI
V6CToV3yKIunTzPlF8Unq2T3Veu84I78Pd8PwpYLzok7DNx2SjcjJfGNpE0/JbCM
MoOeDJs4TQuTVf018c/GKpye8xDcd0Hs45rS2xJHoFIXhgqpbQLwXw2VHq6uaVbL
c/QEbiDnz8IoI/Ocyn1DNGCAWsSd9ejk0T9q2N6VbWguqYZaBTB1FrlaBLD3IL4C
iZNHoHJNTzeR4Zf3IE4sXF9k3FXZdKRkU+a0Q9ecHspSKXPw2wGvMyapa1cb8gyl
tbyAVYDTbKfpUMIrEMmnNi5Z4FxolhKWQVw/jWnyRIhg/L2C9x6ph+DrbNF1PayI
lOaN7q4eKKfD4HBiv/acI266vfn5aoKmP6+EFU2tdF4ALHOGTu2JOYCj368ikfSO
vdMskvnd+USTGNPSOS0tcl7h/9SeCOmqUSQiswbtxdVTBqNl7lWItxR2q8NpDAE5
vWk/0arc6Eb/Q2NDmtYmiElheGWqH+nea83DiNe771rmjEVuQ9HCC26NEPBx9dTT
HDwGmX3OEHozXogAc/rUc+8dKmjWmFk/OPg/PR/XdEfz8RPskbyWrTDqq56VNSR5
/iQ+aty0Ww7/xNJUvVoroaY95OguZDm4CCTRKL4CSm3al6YTQWV+f9lFkKTNr9bS
RoWHCX71EIpBNh0X7h2MTWK2v7FV7nPqou2iGFLqueyGb5Qr5jHasWT9Lp6+e9Q7
UQ04dHO8rhc7kpAWFqYmrLorV5rmSOzODyuTkmSIoLpSvLLEh5PLgIRIxFi9Y0vG
Tq1IUzYGRXdR9DvX3EFVCPUrIdApnxLdBihIarJLqpxy6g9te2EBAfjM0slnjVML
yP6WhEHVnt1IlFYWC96E+dFbFuhOAf9HRKdU8zcBC77mXPY4ddcrEuSN9WDMuIuz
/Uap0D1WKOhot+WAMTsdKXJG2RsAk6QbTzRJ/ixkYadGfNp826R/W9113m84EQ/N
k/jeOg0WaAZxtAGFgqk5SU4FwFdkCuW11EEUkKktnAk0xTjNeDgBoWR1Tkuxhze7
3kN0jKuQXjtHxtFaKOWbcRgrzq65vCXqf98BBl4zO/trhqgakPDYu68VDOgZL8Ex
wODcLBm6uk69KIos53pjQdZVPuNdRtLnxLFWYgw4ba+1/NalFde5XvjI/MmCReM7
FfuTjRFlesavZvU5oLp2hOEZIfaJyzUzKhuA/SiI2LNnqmUzxtrQcBG/XjhYFvKz
K8IztVEzaYYhQBvZQX7ATgVng2Vqt7zkQW8794QSi6oXAWb0n4wViriAdjx8JSKb
5C9AJmLPZ/nyci4JTNuX4HHQQzDmfDm+qHWXG6XpP2Wk+PTIY2Y5iEgLqmnYMxDs
xQISTqBq57Ikn4H8iwmqO28cwTeIGJ7Z+TPATavZt2sWGNoR/dOISl8EANqrtfC7
EcLH6YbJsbgVuN8nieLfE+UNiFEt2mRE5S/cq1f/i0VwmVrP4oWwdVKcRmTKXq6T
sf1UcXPDwYL1PjqwWr1tXyOAsUVR7mh+iQC7NCwtSrKAnh2t16P2FDgjDauxCeiJ
WtMGO5RGuX7rj/K57BRK2FYAdFuHib/Hzs2edLrYODKltIPv89xsm/1IPVddNRrk
NnqfLvoOzSy73DBJgcEIICsXpiPYFIcwL7yhROLjGzqOtrz0QlTOZ8k4DxJowkgZ
zjRerBzix93PzchaYtm2JmNINd933+1LujKfQkCz1cyVCQANNGExJgfdyAPjZ7mo
w1A9lsgyeAOTHzYR3j5CQgfK+S5NUVEMjYAVE5INIXRPTCrcNLsU76esrG9x/wF6
xSma0DcE0zVYw1siNhlaI8nfmYsxaOMuNQ6IoqaNdhj9hVltSjekmBsagPnHI3x1
cML09Dwy5kr8z2S5jAwpgP9OSiIKRsO9dGxzYzgWLDEBl3qYnNaijqo+jevfs4JC
uBVtL+BmJXzVSgdPllyOFctyjs+QiOa6OM8ikJv1H6nGx9teygQJKH+Z9dcHIPW+
pMkXwad3gDNqxBut1J02jCVvJFBoGHOtiX2yk1S7PAsCxABepS4X5pvrZ0WXzhNF
Qo1MpMDzcyNtOOOlRYkVkoEgNmREnjI6aTCxeVG6b6I1bwBA+cqwfz3Lm1qmxM64
uiuNwixSwixib2t4bx0JsdgKBlpNCVSYooPe3fZYg/Ox14Rg1INt/rjCioC0Tvfa
CCO2P+v0fg1VBoGUE67J19s+KegGa29Qe3RnvBVgWTye179KYdvWUR3fdMko3v+7
yJM9Jts0W0c000Yo3/Hza65F++NKL1kwjHp2b6ygJ2qo/eQGwwtVeQzqeeWXho8O
AjaRGAGskABGD12MAld7xKr3Xg2SxplGHampbvn13r/EQsLxT4WWTihcBzVBEhp6
aZfWmhROsARt3K66Wyq8PYERIefICQST6PT8qyizdJxLHgafqdI9hS39apk3FaKd
ypNNzDWFmXjY2orr4sQ6QjO6JbXWOfr0pe7yDEYQohQUe2K3Hcmf4EwRANzbe76V
v9rjNwtC2Zzq11mg6j3X8FhwTfdHf3hhy+W02uiLhg6knZTXUWeeExIpEPmf4XB8
gQXorbpOjEyH1uMxfNrAHiilMeUi1Gvf9MQto7EuA49QMbpmBtvtoP8OnMm8udsO
ON8YQQBr0v3Z34QrHAl7avKp8uXqi5LtHcQcoIlxjudBiHaClvsPDVbJDJXSq7GG
xSSikb6qbHcqWt1Cg2t2sXpYD2wM/xJ7NHrFqjZnJZZJRMsqdUApun6b7FuwvjtB
e2P8uM0Weq0vAFcSVF8K/DFmG3zzwVekDWpGvO6pE4+lCEZwKzTiFnVgMhv+N/iP
Li8FfsNIW2fS+qp0cSUgkje/HW+Qgxe2aTGNAkh4jRB79f5YtVCbEDKyOTZL2MwG
glmvLtuRyT3DhmUYSkrOXp6o0gJUN+wUwjT7CohIuA2Ss8t1mcEO+6WQaGodp/0X
lLHs5l6CPIS6yXoWYlB6EOK4E9z+DV5hJhfMi+PKDRoXBelszmZ7Kd2CuhSI3D3M
DZSSR80ecSj5GaUXktWW8W3izCUYFXj5Dzu7RBQ4ZbYeH37k4RXdH1R/20jKjlKt
3+iXd37jjcQBmCvKcAl2wuj8+YN3eA68BY90bSzm+6A57jO5P8GHO0tv6AehgHzP
Nn2HtXKfXZqtUGqAc5PgEKiPKiMj598JSpmgYXhAWVmTgoBxd7QmNp5DDpzCG6xw
kf0ftiRmuhoO7GWjzZpQKIg0amf97DWxUtCQK6B4J1hhHR6Gt+vMPac902fb61s5
+pVQCfrvSVObul6TDRSq5RqEuh9wg1Ondi2Zz3GBDNw/e/FXr4qlULit8Ha36abq
KopA6ljsVPNVkBCAOlu5fjL6nqTv9XMQR91jZi4Er8kjS0NfXs3Qtl4gX9P9WbQR
OxrMsy04x6n2HikfaXyeDuSKkwJSTJhK5QrgAk2MGO3Ou0Tx21N1/38gh+wPeCOS
62hhVntLkz/ITnJw08y6xNqWKBaPvTur9+gZu9b6DSV/b8aNMXAuyDIM33dnTsYQ
i5/tSjuSVq9h1Di7ARh/0QyDN6RFKRoztxb11becAMZJxtAWKR5yNDkjX81PxZUZ
BXC+ixSD7FcE4P8R9gGC0o0ihP3cSUidwh4/PaldO9OSVmmbFY+Yis7RPuAl4NXL
ZTQTehsFiXJjgELnGGwNrR1N8BuGELKjHi5NoY9k4QRlc32ORQy4/P+FZY9/HBpi
aY4LHWrYZ5rXjVCkpICFUQepUNg38tGjFyB6QbxjmlyFvLUBEJparo7T0v2sXnXE
z0Y70FTY9SX99DZY/eHOrXpnNzoiMKDGhGB1eIXpfHTYdH5lhSx1TwUCwRb2Y3Bk
OJnswtdHFmNuQWfKgo73A27CRNrhgRhurHfNTpsu1II09WwuCakAA4N68b5/51b/
xWysBhv7f7Zsp2sgiKexq0wk3ct+jlXMoQgfvNSL6VkBoJ6cptjZMaj2QqxNVxy5
6D1UqZz2OeQ/jdvrMa/Dv4dbeR2jI/CmX1gdtU4NqdpO4/Rc+XztVEIGYzaA6pfN
Ec/kcunE9KC49jFYvbbnqzxQWBXzdJP5ELQHmMa3M/F/reqse911faI7zzwhCy20
Q7y2BhpjOJ2vgomUMwFS66iTEYlHdw6nA9LcyR0i5QeS3t4ji8nFaYdwUhvjc66x
az5qyfx3UU5wLfyiapi4e1YoIblOBl+p/njrGya8rVUPd+TKmrG/z8rV1auNfee7
vrumUGmbrKp20Dpzc2kCWV5KFO7G7tFkjZrav86wXBs7iHQig/K9h/t2poEZ5BGF
`protect end_protected