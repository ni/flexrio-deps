`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
0+LIRl85m3WFWTFxk3QeDfbWTXsDxyeu5ThbBIWC/5CO6Mj49PVjc3H927DrzxXf
dGUgm+ChJsI7KVZdpzcgnvZXibFeSEirQFEy6O7yZiHPeViZDrbm/gVVTF7VrtxZ
jfF1Eis+FVnFPEFsWw1omSX2cqodL1P0bK/5YhqxQOmkYqxIf7Owed+yjZOTs5PW
SoNI9pTA8pOZRQ0E08mylQyT+q8NtXG7Gnp6kDpXtIUmhqKAhyqmq0Xm89xXtT92
P+1Z7JZMqNxN8ofdOF9JL44gu3wrDuUtdOsRTSpkdmD/+8Aqdwj6mvUZSqynAXMo
nTleCGgelJVIr+Q0avXLW5bVr+SZCAd5XJ+E2031K7yjd0ZrDMTTq6053J5RZ51W
a24JFZahIA4ZWBXHKIJg21DhK2+mX7wOmFerY8p6cl095WZG5/B+HMsL06Tbvspx
87UwDqwt0h5KM5NieIx1Vy6I7Mt4QRS3hnhOZaJHqSHqEZuYOzlkGyzZZnLbQS5i
LY9VRbvqoXNyX+29stkOll5ETYu+DL8Pfep+IEQ5AUV5ndRDG7K6WiLbX9vIgUsT
c12s4q4iYkLZEvV07X0ymxcO3xcJXgWLzUESTBt9CTzcoYgkzuAW/2pbW0wilOe0
nTifjJYbchfMh/i6rrceivks/ptEVyIvxb1QGs797/ZSHB9umz7QCiG8fQ9Kc510
vv6p+QnOxGnWtQbLVM1V+Le/JJ0aF3u+9iw6/8FbgSiMGjlNIvVIP+almv1oWeOH
jU8BfJHWQqTwHSOTqefo4g3BlO/Zv08Wq3Mc3IMm4DqEE7OnoUfYHKbirPrqjaQg
K5F3VQuq3jX5ODhsXWGpra1btf8HNywaFgqn9zDTy1JIMLYOVsxyRXHO64LWY8RI
/8FFP4ZBVqB/ZG9L+9gSK6tnWdSjVpNxlOPUhncfxmnwwbyHC8gLM5XtxMX0N3af
5zNU/I5rhGOMRBI3jNhL507LQLYacedK14mAuCA7gw61SLjIymZ0IZXgMBNdNGKH
8JZMjSm/FMrXMu3rFmPaF6XAqvMPH9NcQO3G+taNnMrzATMBHv65h1YjTbdz3jdy
hcJ8EdJlQx4MuLDwZ4kvuf8uVqxlZcMOcwu5cpeDDq4mXKXvX+muT+911hbTvAfc
fGYeXD+LlOGgPbAElTSlKJO79JC0F3RpY6A4to0A4EHrD1kH2NrW7LbGCL8g3uUL
3eX4f9tHK7I8YDqRpZzw+onCDR/hKxdgjVjicN0nntnm2C/nJsb5m2gQUuLw0cdE
qUNceyEoOndhz9s1QwWQLaYoUHq/9b8FitmfmP+NNbREiWbvTdH07BCqraOQaz/H
ONqmZ1hM8HSRPOjpjeBL2izcb+j3+c8Zwn2ji6o3rM0vV4XohU3hUQXAhqBL6ScW
c7oDmfrwYtDwMoiHlTLa7p80ChDu6I7vIGYtWD+RUQlYkbiKLPufbJoNzV5uy/sU
3zo/0xdP3YzMq3im4i6aPahtG+Sk2+Wp94cm/OEY+BBL+5RXdssbpQ07vO8C4pfA
90cChXtvTUjto71xoCRxBayD+58oaZ4Yad1MCIxmxNEXnE8Yr61ysk9++/ek/V0r
yo8HcZAvNJDQ8kc0ZGkDmzsM0RHhcdsxLjs72CN77NGt6jt9mb2D2UnP8zZvqjIz
+ysAKUSPYvP6Tal7wpJgC8hIH0aB6I/pZuHT37StaM2NlEToMXM+04ytEdSutTsl
Q8qmDEl/yLM7RgE0dlyDPC/2UFK31YXL/TEjqHFWrEWOPTeJ8CaBEHfAsihN3irJ
MVSNiNzEQtmh+cWEAnC//Vth+Yr4IcgLZcXjqplP/twGAYovQRrEOT0ngf4W3ei8
uM8GSvh1HVa8F50P25nZIbDoEiBN1iTerAzebCJFX+GV122SvER4/CT6Zg9xmYS6
P186bI6TRu+AkCKOLbmxkFI7QvZJN1HELoyR/JAJHTHU5ehUTUusG5Tx6lT+CQz7
LEu7ITmFxTXioGtI6MA/q6ru+0/88HN2GMpyBI4pGznnrtLeIcFM/LK7Iul4+geJ
ZrxwPMVfN+erYC2b6KGdTK/cw0qqgfHEionHsJxZNFJGKPV8e+npjotm3caxDhM7
2VzSLcLv4I1JvpJHiPXuj5yEqEp0LQsq+KPgy75NvpiAzsj9t1bnNihigm677n3H
5ZEXqAiSIn06XFnIBBVKrn0AOvV7lY1POOzTQ1fC9upij8hRDbMqk3sh/v0mq7yz
QPAru86bnSz+A4iRmCya2r1RTwyuv2nn6G7EWPCei1FYPGKP/nx1QFOdKSgVdkaW
pfdolZ3jakA7nx9H1zoTwGg44IHyfQ2YLd0vXVM1y0MMbwD7HGVu2FAJ1TzaoAnW
rzNwsA1eDBXhAQyqg5X2EqQzIKUgkNCxpPoffAHf8K68c49cHSIzu5QPE3iKCpsD
SrPzSjqB3zeAUx+I4LJ6eNYAYbOYk1eau6j4BzSvJNMn5GHzaQY0qeVQPOrcxlbk
T+lbGQxwBMoJyM5MRUC0N4uSt9rGka8j+y4VIZ5l+PozlBfMaFJZasQPnY9pICHq
/L9jGh8Vjk2L08fmZUVrKyG0/LAGtfM1jGv9SqmXZ8vQmPeuYSMei1OYbwwbzHag
ZLGTm94U+kYjnJk3TJp+34k9vy79lFsIMsWVvRKH6KjQg3MHGyEK/KJPOnhJj9dC
a6L7Lym6qa/VmMldss0ERYQzPBGzfrxAO/o5BRXQiNo4ZKiarRzhBhf5zzqRxCZy
YqySJHw9h/lU50M8wKTUUpAsmXANYkH3eJJqmiVARAD/vZh88oB/1cB1eI3v/AP3
KkFaOVLzbSItJ1bjJd1zmqUE+RNKu5Y5xX7mBCEOfObrNIXsguNwE42lfMQw0tsZ
EAolQrC4it8UA+4mDks4Yid9CSro5jQlWuB28e3BJF2dyp7OOGO3pTEF1CWCc/+3
5SP4pihR6eGHTzI2lpc2lIa63n+Ib71iEBWvuKE+9TDHh303IZAmrGVHItnA6BZL
kpccwozpBahd1XqzXHAaYadXR8al0BmQKBJc3bVWbvS4yl9ShXdXju2mY+itbbc2
TTdCcrlg+wdVBX+frjd9Vljr3mDyFfflYraBTzhV5RGXSiT9QWuZyGtn1fcQzSq1
6y0D5cq/dkXjOXgo91WBynfGlv1lc1SR+1YKgmX5Z+rhcUP2NfZCp/LGO0a7Qzg3
DwWlKeiiP3WyZ7bzqXU4n1gfYzhzcuJmGBIx1J7+vuzLOO08OfPeRgaGlR+64QT0
EZcSfQ0pVT2v9T8TbiRSSP1Q+KbxoBTnZ9e2swPaV4HavmB5lz07Ugd4KPGxJdo5
M5g90ZeJGaFoB8/fp17uZSV2dmbYmZR+f6YlOUficGCrEgXyaRZHqgIxzoGAUi7T
noVec24T7AYaNxp5JA+IfcKAi3dCXnX4L/xYXrBZDIAkgZJmkx523r3lwtAVk5d8
4cqNnKOABUHrGEjKoUKt7eB49zOJ1Vt6G8Fi2KcKeagc/LWIKyguXRmN09/Smmgs
nHJt7ehdbmXKF7V0PhjZMAhtsT+p4UV7/bADEMnq8Atpmk16dLN7qxApf/Ac20/n
AIOBzRf5AzDLa//86kNPhL8lCn5xBMUWClb++Ou0oqKOXFTW0jQ6f0erXXq/zB8K
dMEhJl0rYPNxENA+fD0dgH/XKNfP7Tx7Vzwsak8WeEEzSj37GfmVl3v1cCXPKZSk
zGafi4sIQ2HqNUwi+5tjOYbxdXGoghC1g+4Bn5TCCqTRZmKVTC+l/bs8j5Y93F91
LavdNfVvFN0spuqwdH8ghhwtibnW5L6YUAJoIRV5adx7zxLmlzocioU/Qkt6bjBk
ggEqIjlLpofL78RyEPqEvTv1D2djDOYTPQVpJ6ItN+xtJ2n0ECAiCPdwyK3WgnCn
+MPH2XnkS0snpdY86PWxo+r5dtCNy0UPTDxa94305esZgOxNzIXh7kpjbxguCAdP
4ipptsX0N7ICWWMq/ADAjEPFYgnQdwHjlxh37EVkOFyPnDpmAWiOkIbc6V2TKky1
xKeNsOSbENnUFGUjHZb9eD8B1ijfyI1mQp7un8xDsLlTeEmIvZMCj+4FwXJs9Oqm
iD08rEIGLdRDwkXApFzlWXhLfDFaiveDVYDrbF5pEQB2Mk7NM8MpiLjgGHBOlmQ6
/s3QN9k/a7N+bIOIv+2iATVRZhmGl+vovs8VNLM3VoRdALuqPm0XQU0fubDAqG5D
56pB+6DKR7K2IqDfe6e1F4iKiv9sboR6Ofw4Akm0krZy7+H57GmNJhnzffE6U0Ey
s/bxq3Bvjafa6DqhR9vk3OLtW9OLUU0bgP6xdHP9sF7KnA+pUjz5omdXJ6VAWEhh
lYXll+cTsyJ02RxQ6cpuWL5ViQYFzutrVgD17om9Iqf7JzrbRWKGYfZRcy69+HQr
H/Znk4xHvo4Gxdjq57xM3I1R6c3U33/avkr2hrKNUhauwGsW2IHUUqBRG6FIadKN
c/y3bNyLQ5A+wM7fjJfsSGA+5/+DPNs23Fv7En9OfjGgZku8/HkxRCypLl2cvHxF
YAYz4cxz0A1wGVs/JP1VZyPZtMAaeR0AmBo4BQsH2T3q5tSrhGMFT9gAS86pDzrK
mRsxPrfGT74IiQW4HYDlSjq+0HItSK6C0Gkd5Lpk/ohd/6aXeW79KZ+O2p2Kww1c
GvAH6AqT16yd9BdlFUKLFizqKRXohfCwvbyrQKJNssi+ZCUjU8So4yEsDQMsYjS3
NkDDGa1INDEEAH6lga6/6cdQ+Sx/V86kFfOyKWVJQAoddZKcWEOeNq4YNV2FRYmg
+lRTKBH4J1BtdX3Un8LY7yXOh2oKZXl1+0FqE0CuMnxRQeVzkVKL80/6/Ggvl61j
ZT1YnJSoo/EG4fhMxWmt6Gkpzh4Gb7swuDiKWV0Drkkbam/0U8y54oRjaXh5R2O3
qCU4EK3988+W0kMrgcDZDJ0MLv5o8xCTeR3mYPqJmW6WAAlP/Nsk7meZzxcfie3f
3QYW7m3yNzDHp665Ksm8oOGFeITpzSLlnUw3+1WoBboAoSbYPPb0W0uWKb78fSQe
o0ZLVtagXZA1G+nfdqIlojxbEl9kk/AnLltAQDsR+dIiPv8S+p8Ikze6AeQagbxA
3otLdJEuJM5QVUDWNQ03CmXvdwBqTelJD3UDdMEDQ9A/NtpmjSKimeEKA65DhaJH
SF8CIrzdsXBZM80z9bN5nTXtHWM0JUUw5CBjgpCMmJAiqkG6nJfeSwG0adPc8hul
ARG8svW7dmf0T4+aBLimgQmoTy0y+BFfaLufCBvb/m75el6FHzMi7c5qXWDC7DXv
z4lNVWxNZE71p92rNCzZ1JQiDUN3LlD9LiEG97OF5XLKs3kKItfRd7n/0M+jUv3I
/si5SjYgjgQ0+r6BXwMdIe6o4cmkuUGKG+j5eJboXB4r7Kdh1HVzG1VYNnznprPL
6HS68UJ9X80UrY4LJw7uvdZIuD/rZKNo8uTbnUvQAi/+SY8Ph2u6Bx53m/ozejVo
2mCXfDmfPO7L4DW2tQboSN231TSwuXHNs25PJP0/KnInS36GeCbWAbCbINsOh9HZ
CpzOuAm6U35aBHSBD11MOEJJM2p2cllgXIOJcdUKPaCjLv8Z28iIywoGdmEGP5Tk
pwGmGk/x20ds/Bh+sUmWwId9YvYd+CsIvUkNGUCaHbF5CYBCZ43X9RDqMvmtc7dy
NTfrKWBIe5iesTtR+fCqwWVWOx+DqSieJpSYb3HGUmc+lg5bG7NFE1WdBVluWRZ7
K7KH6ugHZlT2F3x0shYLufNHu6JANFtciJmW8l+nu/e+gQMEzk/GItsuukJs9E1l
r7rI5KczyhR7xEXgPOvF72fzMW+p7iKgV7aS6c7o6GzwgZ0fwk2gx1tpvzoTZGjG
d+Fn1BWK/2TyAxjB95WCwwzpJdp+JSZ9PsIWNw9lcUGUlg5Zhy0UID2AueRGIUyA
CjJohBXXBvkgNJPkp2M9VCqslyq+SpbmPFf5oHBr/Df+iCkuVV9aYQINkfIPGbF9
8xA4VcdnCcM2b7mkMXNWG3mPN98HJjDxU3FZ66olJafaix1ZeeEbPkry5u9sLdjX
t7A393hjvKFJpbsueSMpwT9Ufy3yaYHgGvcxQDuBTz60W1REe6qXpG2qLIBc3y5W
rAmTr9fKkbjEzYhVjPs4Ju4DwzUU+2Ve6MC+28jnsBjxaDEoK+iQ4i9TtsdplOxl
9jWtS56r6fjNM5etiwmw7/WAjzp0+K8UMXVisHcLDmFXRNJUmAZzGKn4XNsQg02A
OOsDsjWpHASv/+S2k3Q5wd2nJafoWEkX3ALURp4hzyq3L4hi/IbqellCInLYwuku
VcuJlqmUsHB4TtRTqJq3HmjxzOqltSnJbjLu0hNdODOxxRPhqQgQ+83V9pwAZ9ai
Pq6HixdWNb54G/ZRWJEXY4nnlS0lHw1BdSwmY36JkpkNTf4NqS576BQhe7dAzkaf
2fsDiaR9zhu/vxmax/8FFcwVeuG3qyTElz7EQXAWrZFy6xQT43sEIirbDWru+ksj
txsBEZDqPyAxlAE4mDuNZ0SHUNz7qKzBh4AFd1qH9FvHPKNt6pIdUtMA4zddnWZ5
ZuqJgQAib+JYMZnJywkk7UXWFhz+Gg+4t4lRQ2ZoHYfQkK+U6Rw4uE04y8IgblwP
Wq5VWe48D+w6uwlB8D331Ezf3P2BgsOPAy8MkJccYBAF74RJasNjDfG+HEIKP0SQ
WrydFoOnyCJ6Z3+6P/LnLwP9wTVoSYO/hrsjNR9MZ2fAL/RJpGCKAak+lT8QHNiN
vr2AbaywUvL67rUckAX2EDC6KC7twc5zj0rGaBfkFh9SeM1BNnwtRop0tT/L2C9L
jGpfkMahZHyZQfiH22OlgHH2s/MbRVEmbeX3Ao/1nuLzdmzVytWKvGRMo28ge6Pl
t0ZoJllLhly97zS5QF/vSFqYw8byv8aVGVQO8gE0WAyWPV5joGqABb1F/pf2YYvz
+uAdd2H6R7OSE+dtD+CHqCZuzHhQrS9GLL0OdCwPfdJVZXt79HPgMF+4Z9XHjqDs
MNq2oqvvWZ0sP8T4PTHkmL27ByJ6bVqGHKtOLDuitOOD1HWpWWAbWmSdztTDRy7U
fgTJ+mavyrHquS6Hy+EUZ9mUwNgQwvKMj7mcxj637hY+XkiGRqWLbXfA8AwmtQKc
QFHI6rN2xjS1bVSch5yO6GVKOZ+CSW0TJ6Par/PpE1mMERiQxOdsYH0e4H/DtH30
yQ/7c0Ew8ZMUC26qg8utvUXtj/omi80z5fjwqLMiOJpuaPptXXwG7JHz5obLm8OS
svlNOdJe0faZR6jCXFmmyQ7xTU/i9m7vWtKxIstQAgnUaWyTZ4qk+iAkixcCdPtv
uUYZ9/7jbtqq8pWwmoFEVJ+ogIUpj9Gt5BeoK6zkBluSwDF1/UHiWgZbyeq3CHEu
+2aZ+jEYtmiqdzDGiqo2L8K0CEy8XMXNpUK22bUm76QzwAkIrbJOM2LnvsOFv9Os
9ghPkgEQDcU28Hyr7wcJFmgc1oqYdCot5GKD9fbGz6ZYKWXfBJGFVnACbf5DgIfo
bqXFlQZrC21jNUqOWuJ9bRXHlZBXFYnxBANZ6/+xeIXXx/ijgJdwjf+FRgEUsFO1
i7yfWttnPePOylJCF0sG/PweMlXwxKuXlLIZ3sN8ejzuBuNoLij2UKihJOPM/qCi
bE8B1RiMak6+lUVbIdJO8UABhdrih8i5iSAp5XxdMeEytWaWnxZvyKYjOGx7H+Qu
odz1mwRsK6RmvwdpDXgnDFPOCb4E0cam5D5WGPGqwHKgdUOTkJnUIlf21Lmso5JK
UeQp2QIaJc/uR71ahLcYlO9yH/GQARpLc6sNGx1qomE4MRTTQ7AR6neaJnQVv2wX
CrRP42x7jMf6VZ9yLnm54aUPgThuzTnR4rJXYCKh8RCm+fNI/K9QemE2vCv1WdJh
UuIqkyLeWfCfFQbdQvG2TWutIqc8Kc2LdkJ72gI5qfjGem6hBXZYujFOuxJrK947
VRiL8oSyRu6SE5Xwz9CTGZ3E0ae+FBAD1hVqjuG26MEc0KGylDHwI3QNOPBj1bpu
/SEdlJK59CzNkocPmTU9smq+OMr3Fq2ioLZCOWST6lq0TEOsnWq0HCHKHxSVq74O
5NnfUfaOTAjoDfBDf44Vi2NMlybyzLf/tszinz58PsL2xdKEEpfMuwbZSVli8iq5
3SlRq+vXBtDC0no0EYZ+nszZ7mox1T62fHJUAihTMcRIFyP6QLJf2VwIayUNsUWj
Mn5DMza3I1xNK8tNW190ec7z7aZP74l42WU32rWhylk3ED6651ZE0GasnjXtjJHO
IV7zzX2JtJ5n6Tj25JdEq7QtAefRhbNlJs6kFCAqTedQeXdysUmhWtqgFRP48fge
XZrCi7eY5a0xDW0QDYTcqLHBbzQbPwVX/PNCp0GxKnPVgusN0zShyP1vKsTqdCNE
AYFEFaO+UY6ZUxudPj+UjrziyiRlG/6T49bF6S+8Zlr89Wyo7wmTKkjAEnT2gEvA
XQTsDBLLDzxnCw5PbzxLfRGvnOJo0oORbvUKdpyQxoSYAZPoQPRrjO3CipGHkL4E
zebybFUygnu1sSBeiVzm9HSK8TTbl9j1DRAD88M9b/DFHH7f/e0qcomcfzDUoRTw
y4vib52XyZvPxtqvGlR+DK5fQbMcmD5bPSotv+Cf/rv0e4GItLk2Iir23qxK6FJY
cR+1eRUyZG1hVw2gqwAHfZp2tB8/JvebnaVJv/1mBHz4cOfoNX7YMcpYS1FWbbem
H31cx+V5zINuYlJWZ8WeeeU0TJFAm5mwkX+OojodKiRQCpQzpa/pjNXSQFh990xa
0mH4OyXcjaUOO6/Kwxf0pws288QS6Izcqi+1UrMKUiHAuggdQIXnfVeG7HTQfApO
3JGwRnFtbI2h2uHl6GN9++ejPvQdrwBsxB8pyupGIk3rXdEvu+InqExYtbmXYNBS
q78yr1jhbzLHkWwVKZ0tXiMGokZudJglbhkmmeqjnAuMvebT6Hjp+CU0vXZIRA0P
j9ZPjhMLmnmiSOC1e1TAfAl3FAjqgraPshUyvpph64TOceCcRuoFiJ0+VPmqf6Ne
iqgWjxsdok6bp0m7KZveMk3JTtIqMd8UNN2suC1ZmtUsmCAFwv5LCYAMngYZZtB/
8fqrJE9zlh6Mrf9crRf11F/FiP64dG2jco+2wIfuUsO6eqr6oYJO6U4jBAeT7O8F
QX3MnUId7itB+N0y1LLwNmpoi5TN68G/fBQFBiDJA3AWd4QWEe0A7USoxzS2pu4l
jEu1dUgPSZhZxpNH/ni7d/KZGHqjDtKt+mIhkXYOlRGvBIzaPcx0xCLOysA0r3us
B/rgJ3PFAfqKduUxbVp2jcVD+xe3tWNfaKWBOdb/BODLLA0vOIJ0IPE4Ps4vYRfI
iREYJmGrtaIYg5lswNn+WxNe/CDRBoAvmrSDVf4yu3wuzfO1f1aItyfn0t3ZspQP
TPz5FjR83s0FSPKfFaDyXRgzHdCeRSeevrBdYGrkVGVuyQ6Ara+y+ybZJeIfaB/U
CtLKtomhzrahsIqFcjv9qao1qvpCbZJ0CM7ggveCkBonZYgWpuPcwuO8xQUNpM4e
aRJTZmR3N1vKSexefEpHbh2Sa1FacPq4HT4fCzACiw0KGTqGSTYELHrB7jlKYNwU
nV6UkEdizc0wMjFhM4LQt1V0MXV6gqAcIxD0GDMGcgDh8hFx1fUCFbnTcX+prRqD
5Upzbvxlu65aK4lOinMAl2pZ/g9zzknvHyYOP8XO9kSt9pkgC37UP6aq87mzySeE
mFXBCgWnOr8b0oiRQGGUAgVGOZUuBfKF71Xiolzl3zj05+5Em1m2sUTZz3kWnEQQ
Fg0+e5Q4SPNE+9bRP/CKos8WaL4Snw81cPtAM5v5+Xq/qYX7WN1kmjZLKoxCcfD/
HhoHgBMYTy9+/zVWD2jKYJ1jMfhtck9RLzW6/6UFmRdwq3QgASkh9Kn2cnFm+imt
ffmaFEJMpDznXwHep5NKIHVwSTKE4OHA9DGuCr6cepLBPZdg7fKjhMjnK9pDBjW8
RJ6ALWVY8165rK1tPaBd8wtEEv7hHzHkWQCWhM7mA6tkZPi2iUK4D/S6JsqFahXP
zyInDEY3ZaP/bA5eEaM8H6XPDBEu00cBmGYIvk/f43VBpXT1xKIUBNuvpp/jLkqU
QkOX0SFxd9fdJ826tlreiPwsA2nyZywd1x2XPBrb4XU/FFC2uor9HhBQfirFymuC
IRheK+V2dc2dtKY/2MEdPh/Iv9IXu8laoHvQRfi2yNXY7QOOqkrwlXoqERvqk593
atuAyd91ZdAbBD8ItyP+V4L6LLoVXcWxwLQ2Wq9BekdkLZmPqIIEHXC4CXC84c29
56ENgExIZCyB+9d68X85iXZl0DzYgYCn8PCoPLdvIqjvdcZcZPwGscYWo6taGLPM
LekIAy4dkpfQMrvCqn72W5jgVU2XryoWI01UhiYixkQzGHnIBajRdEngUCHAHyVw
B8ciulPdiCrsZ8u++Wlt9aKpLGOIKIsxjZV+JNzPh9qO6a7O9yOU8n5cgZoEW2Rh
1KsSL15ohcXNvOaKIWYsvr3pMoh5iE+41MlKp00yv0JjhUzFj+TCJDn5Is6JIvf5
sraNIund5CcmMwA0GbEBFRBEF6FW2vkqNxWaK/BNPQGD+KGFnpnX7Q3EAkrXXZB4
oEltJhCcBKNtu1NzU69nexzcdzqwr9s6rtXFHWD+3CFonbKx2ukw+qknE3nUdmsM
6UpDCQfKaHXRyaLyMSRvS/gUt4gglN/sSwv5edtg+6MvF288K8B/TNRIxrm4naNo
OOrGgsvxxG9JXxQt5gtKUgfKyrovZsGhGZHxQB7CUTOUZ8cvDTSVmChHj17nLbS/
F6uJUzBdMHxGVX9YSLAauJK84i8gS/w5kMUnFVzFIk7vcY5ebQXur6+5ED6Uc/Pp
76Ke0MujqWClxnmiO7u3ZNQkQ16XCHypnqbAUouOrWJmwM0t280wCqi6tiP8P4rD
W+PtxUGA0HL0weNG96RtXD+uUY+w2r6l71vl7ww+KpvnW6FYUHphMjnfx82hP5l+
DQHJK1nTP9Ep8T2Geh9ospdKHSELq5cxeEWfJpJh9d4LnpKAlf1gUW2l37vfFiAL
2vy/UkMblbLfSd0HVnsSVGKNNBXIl33mA+yuNch2GmMpM6SDsFEGomf/BfkGlP23
SEX6rmQqMq4hFVJKyXO/4cJzhQDOdvNpyxUNgzGvm7cpf6Ez15hKmLyA1Ia8Ajvf
6YtjsibZQxujZd1grlIxnhKFFiCrKvKGhzWKknkweRJtkMgGDtD0NtHadIl9mJXI
DdlypbXoSvnj4rs7fkE8v9ny1pMExxCKIKX6UXB0WW02xfHP8mRlSPWqWwYv1BhD
SFgFOXe9u5w5HcywJd2h1vTUGfdlnpP0XqlIGrcA16Bhjr0Tra1uLKharHBrJjD8
+o3267kw2RlaGVL62+Xj7BWMMOo/DBWcQb7FKkaJU3nKAE4XiFfx7CSSNXtoLBRi
z2Xkdc7JTJhySgO1pX4GJkaKjsjSTMzOJv78ogP9nyPvUAYfFEk+wVvw+jehxn7d
E5Xl3AoNA2+jcFiFSKqhJf6ue+mbJSGitueUWADQmkRYxPlmdXgz38I+Gtamm/AC
oYyGdYlp6RoXRGm9RjZyvBsEsVfG0qgKEQpJ+ciwTW08MQRiZbnv0O8Gj3jD3+YQ
xyn1/RgXg52wnTgmamnXq/KNiMVRFvuaiCBzp2op9fi2xfq7rrfm9/TJ/DDFiK5l
ktmtCxsemfKLQmZmrFVZjgOnPricZNo9U+cu+rq01cQeHwJApVYVT4ILWYErw7dM
f6TEQSoWgMfoAbXcyGKY2DBlvcTgGBp0o52Hbpgf1fZ+PaAhNUqzymKNAAOcTSVr
rSEglvjQKOUl4ua6yCKTqdLEUD8DthdcZ2xp2J769uxEWxpQV4ZenBKSzZ7eJOcn
edhB1g4Swk5BANdd1NUWzJ0p6hW5eDq+8Q68kq5c7P/4YA+T6x0Cl6DBb7rPdYHA
FG59ogEKcCKzy9Giwve9znYL1PyoIQDiv7Jz13WAGbr4APSm/gIQP+WK8caNrjdE
47TEYLg7rvpvE0LoH/Tiv63eZppbEThAcyKfUAQ66o4ec+Rh7sVkv5ulAyNXVvao
Ls9E5Dh2QF3NgAmzxq/A8ky8dfHd9Y9dpAdZtCA2q7Sn4reMf4/Y9wklSrbvrw5w
P4Oc+dqETX5UBZnkt2SpV+rr7pP1wrTPo4TgP7nan7PNxA44augCPloLMmCb3kBD
CSyu3U1stsj8LWsvyMSWVZLYKLon1uI4YjA0+cilmLYo5MeWtj/L+JIWVluEAjkM
hvlVYWz5i8eItKkXMkZKcL7Wx4Ww3YBaMPntp8z1X9WrjUL+IFKtMVlhhQ1gMRmi
z+Sf2xRHOzhGL+SpfAfbH7BgLMb0S6kVwBsmSNDwKJhI00KS8H9O7YG87Jd1Q4Ts
mBBh8RM8j0l5rHHqXJlmw8Gv3I69Zy9xQOpPbLiFZtkzH73jIMAoe74NeJjil0mf
16M6b9GuDVRcFOaRaty348Qgs5i15+hqgSBoFspQFRUaDWf1GX+CINnwCtFbyDq8
rYpo91QdcNWAStJCX4FqQ74EMyaxIH7l2hHJ2hVtInOjBjOiq3KLW4AqvUOcJbTm
++JIANJFWsZ1MolGIt3bt8cPDOeQWCBqGv4GB4NsWNUTAwTsBA2r8F8LCZd13QB8
zN4pEYT1jACBIiyJh9NS2q/UDNIMxqk9bwrRVNyyBf/ndfKztXaRbmeFxuEREBcB
0367Oq8fzPrTOsUwzTZyon1OCwBvaOmLNzudMsz9WMXsaCTD7BjFfCv3A7BBa9V+
jtNjWICj3+6fxo8WoLwQDMagNfJAeMsEkAmRN2mE36yogjJhb0AVNvUMiISkNjhJ
GFrZ4tlm19nbcG1hBHwDJJDMBGvIZov4xTVO2xDtKj4/LHxj2RINxE6H1UfqjVJ8
mtoAZOQDGFYVukMNq3WPtiaWyf5YwgUwz0rnxm7Z19YP5ZG1AfgKQRBePEOTr5w/
kcLbR/p2ESSWAVEliLsrmfVls4PA17llqD/YUZ+U0SzMNrObQp55Aq+WDBfcTPiO
GFH0M4Xea0TtHWo55bZmzjHlvDpNnAcxX5KpZIkUgudP0yIekr67zcqZEHABQMK5
P/R3f+48nrI+sIBL+WdZA8Jq2Bui55gMuu0focBNJV0UqAGZpf77oWmXVRRlZk2K
oiAyUqET2ZjDTy48C/adPea4DtWv9smDGAdeKl0c1/alvuRT+0qJ5wY3fSfYt65t
xELPHG5m4989OMa11eeaZLhx7nOF7AZzIwzHw3sHx6t9HiT5DJywFwJJTkI+fiVt
lZBSsPrh7OqnLSyOok+vH1DNSY/iQhuiyI/Yq84ugVyFk/LmhrblGvusqxoXjpfE
Q1SiNuIYijcmx1tcK+jxVMCFkHldy5LYkFbP0L2k+x2ZMDEjqNUfQzDpwA5Q7zlN
4U5e4JO/QfYgGvSWTiv1FwfLJgpl1F5HPgSivqZHbnKc11Ioi8Exj526T6Zho593
b6gcd5vMy/kPEIQW/+EPROyOh6GdX9GtB+YWlYiJhpxyPZFrz6NFMiBlRsA0Za7f
kv9IU+PNzIxdoDej/KMjB2SzMOsVCNS5owllpCTUnYODpAvumf33OhN/O0QGvKh7
HhIE5LDN12uDzwfUL/radq1lfhHjLtI8POvpM4SitaKmJD6rKDYLzUpc1eHoSYSf
JdCLeHWiet79VO4f77MsaLTyOKD3kt0CoWX9sF9fCy2gyVruQjrbsvil1LIGikz+
u6Awffsk4UhiqX8L/dd+KIQJLjHFdT2NEuZ6JO+vUBplXDfNk20voNrFE6Uk6RlZ
2/udWUqpve+C+pOZtGPA1GvrL8qPcu7VkjgXLvgPb38WpPHr7fl56BMdo+dGVkXp
qxC/X/oaAdL1ao5nPIffPBVbKKkaHdqtRsDc6XnVdYOo8wrxtpKkC4fMUCMNvph8
id09IQlj4t7ts1VYxMSgzU/eaQMqrkbFG3uoIIAwwFvxbWTnqjDOfLaJJri6al7n
YVSdKzNQU/AOQ3jmEpG3veCV7GGGzTkngvxuXAo6HB+DDk1Fgelqwd8UqlAsHOam
dogqzagNfUkFI0DcJc1eUiSz5RyBNJJ7m3sFqF81n3lReVx/iUpQYb8RocKoVwMQ
TgeAyBUcxewX6I9nuS/f5K/d/ds63JU2zwgtQqkFWQ4CTjPlU5EnZ+QiYOgQljng
hJv7P4ogD2TA0CH0yRQVPLp+qcusiTJZiQjgoUniF1ZAu4h0K1hYlkOf0AAAW2cm
MFtbIOIEXeNZdFd/xeKqZ3gSRWONmFWIA25j01+oyrbmRTWRsUvp+6Grr8Zh90gV
ISlYIakbPV5B74weRH8+ZZOx5y/EYk63dPxOgzdzzKPH/CxMotaV0KyRdynhz5rz
nHtV3iptmY7MFgwFRxbO6lN8U8l3btxbUAY1kA/H9I/8oD5G0IDvrWoPqAo0oXBL
u43DjJ06CDV78KAnCHYGVsQe8AF4Y1zmGAFHBupA4S4ORUld3ene01lPIosOCfX+
NKnrWY3HUfils3U7S1BVykeaorgDObQmItZo85QnIukbZbTPlR6LLPVPmdhZmA1O
6xImN57XgKktIP0rmp0k6udFmyF0RWIneh9zffkVMSlYyuNmmRqnQI74dB+P6MAf
Py4Us6ylD28NOe4VzRSsZ/vTKKQwoMA00a7htjCIkrkqH1eadZzHRWu5lfMiRqCT
IbtUFlcY9FyAuokmQWGTzzaq2XR47PPAnOAbmIwHYwXWfYBQDvWmNVFuKC1HOJI2
trl6xiNxayO2/XOSEpucBehKMS7ftltzvUtV4bDW0uWRdYu2L7c+tr1yOozRYBVg
6zAnDTmqbimvVACYB9iuzoijhpPJmxxFatUUs77B9lfYQj8SoTWnuTWS9BwJf0eB
ABMJYleAhXIcnRYGXz4rczShaJwaNcyaJcjqoVq0V1roTS2/+TUrD6CBMBAQ0bsk
DM+38OU2M14WPUL17id04gUSjvhTbvbKsXPjGDm2EqrY6Ia+zhKbbhL528btYRko
j8UPUnds/mwyXukBrlZFsZpz2JWpCoZJ8HTXNXxvqF1+JH0vrJn+FGr8fS2OruqV
mKYiqf4fXJg24aP6EoSRQG+uALxJQx8O3I281m/PemXIvzdjB3648yv0vcfg+OwI
p8zdQZeXQaVBgJ+q0sfyGlvgFBIfJV3YYUHtlx81Oh2QWdL8u6S72Haqjtl+Q9eb
zsISsZ/RPXcv5u77obCorGboKCXDfHmq4q2mZw8TLB5A7CdxGNzHUbJWTNxqkY3G
RTTOM4M+pogtQs9txtbXqcivQ9vz2lUNEGt6po0BNtrxKTNdGMACvYmqTn6X0HYP
TgDXqGUPfAxlRMdPHRiQjz2NwbAk6PxpTKfU4mF2d9QSb3dLZPunfjRok/2L9q5s
NxdOO9SyL7oh3hq5cAL1/tSg6TZB79LmVnl6bmrMO+zdXbOTvdvdypdBt51dV1zn
DrJxeWMqP+r6eZxFYcfaBjywreB1YC3K9qHfHbYPAHcj2nBwx1Au5n2iKtCZFZwy
H/3/Sn0koINxgtbvQk+VOkfPOeBAKLMd5E80eaQiyMMueHUYtaXu3da4Q/ktFc5S
kYhO2itesHlZidm9dhELPy4xipgJWmmSPC5up4vCcwE8/V+6mPfH85yxLz2UHw/r
VpgYyNBBLNf+UAGrdNDHFdxx42BdOBnQSZrLGlIdLGfW3ciiNhtoninkzqaGkQJO
GuaN8mlgHr0W/SduYrOkqd34YrVvy9b7VVXj1k0PcZow/D/3AEZHLFXDtp2ZqiWW
NjKd7WA8XWGueJ4lCOlXrNHRtOPNqfGrN1yNAG9LZht/jP1HPEqUZ+pgodrPcbEa
5z8KKXqb9dTy9LL000DV2njzYspZJNOztbfqgg7x/4uXHL7KWZeN0T4seamtOP+e
PSTRsi2l3fgnPv4k3HfSuDzQhdpvEZwcKeyWj2NR4YkS7kgBLbcD8IRIzKv/qulk
Oy+mTrCEgDLCXTZnldvRGnuAX5yFx2/TK7vAcMpXgW7kLHG4hQjodM5JFrB8eJ7P
dDG90CdrNbGFfjnHatByysJ7guzVpX7EyYyLjK+HhnLOS/cfxS6yTfFr5hfWO5qJ
5fZdKMaCGaUlSkikhnzsY6F2FCMaJYoiFZGYtaiNj0bFuweHF023Etgp60rMkx4z
lPERrYbYjUwy48uLdftinMh0WxKs8GouonK8jNW/gGHopiE3woZonIPrXpehsQKe
OyWe8atzfRhacOENO3IRmyKz7oEsboMHtYJQjm8pZcG7h3e8MqESqcKY18GULusd
NDlV2ghJKjz/ARen+My66wArhn7ljUYJCSKFDatb4h5xK96TxJdCLEam2oQB3Ojn
fgu7QNQnoJQSoxfBxFIsEk3V+hNjR4oQbbsoEmCD4dKZkcZrHx/qKYb+01OlLuam
LZMiNkmmgGyhFmiBG3n09PG0ZbwwZnTLGTG24z7sPbKg8hRoKEq9g3e1TXLoq7eW
f9qGglWhzulWcfpZGfJhFOBnH9yccK8KTnki6IiTp+LkEaxLeU8+0CKjuJxyLKHX
FpwsGqul+Z5q0vaKyeu6jtkm2PnXm0V1VLumhGe+y0oY3Cy/gP4D1pGrWfqDa5gs
qVJ2XqdRrDU0XEyKqOanzVU3XSocsEiuOZQyIKRhb1sIxJBv4W7M1tkFmLMlGPi5
ciIIVKam/hP1lv6ouGRRtP/myKk9oVyUKzKDE0y2DD9TedHQhvgSe4D/+rCwIumZ
mr4K/j39J9LD6b4wQuTbiZVWB+o7PaFViljga1TnaNA5kK01ns1If3YwJoqsaBk0
ii5MXAkbnuQ/IHA65i7au8EZD07jU0lwSIB+l+qKOo3Dfk3q299dgJ8vvXnvQyWf
XvOsEhCAKI0YD/zgxzIxJzCJsB/Guc2fyVS1g1QferuPaESDmj/GBNOh7FBOXL7A
CSb3yD4LcDmY9xrKZLeNdp425YugjuatKPuR8sbcWonQDpcjRAl/ZVFHrHzGZcUv
dxuBBohwlRZroKASioQYQtIq1hIAFZWrt5G0fQQq5C0ovShEeWjD1XdPwgTCuV9r
UzrYGSe79Hf/WE14ZbHr89BeuzgawBpMef/JgV2Vg7MP0OLALzMBVieYjXC2qW9E
+IC5xwPx79ZuWgnCm8eiOHwXvtIaoLTEsGC7uSePq00eR+COcM6M4EPlXTIQVcwP
sSq1HbIJMcFNfE8lj2urVpjEaILKRoHPJJR+y6v4RlitaKT51GK/Lr8SdyQrZ6Pu
PCm04trfUhYvl7wr9mfE/kLWg4dkC14L2pAQAYLgDMQuCLHs6EddV6q/UkyhOiqX
O+Lc1N1LhXn7K8ZAc1LvwB1y0rNtUgj9EDdGJPID5svftcGEUQFWwlV043xqyqKJ
KpLpaMkz/lSHSt++kNKjywwH0j7Xj+PMSU86aoz7K31O0k8qe2l076YX7O9XihIY
un2ZiFbk0RReJyZ9VkkWoGaB1zH5MGaoG1g8ODRtfD1ycxaudBprqBB1Oa0cGuMb
aQMAtDdud1dJU2uPzkqsnRdb+QQTYHCsZId1LRKoc25VOitbfo0Kc7U3DVm7N285
PENcyRm9morHzOmz9A6h6AgO1lYg5Sfq1iN0DoOJbp3eACN1Qu/BeK5ka78oNlDq
XsvHZnhU8o2NlQfCWK/KiO5jOzavIvWfZzNab9XHh/YaT0BaN7pavLwFuVZIM7CM
eIsIxQTdeXYXikQxmahNAAo/H3DlbGKf61q9hJIcYee1prkf8V1CHT9qLtWTkV3B
KFDbqfxLMSM7faabBjfrHAE8dRBRnnKyAZRMLT8zLLUg45WZe5WYxc+FgNPHftub
aav73o7YcdLVXLf4Fz1eGu+iEzSKJaEZ2ZkkXewE6q9Xm1PW0BpnIU3VKXJJloxN
j/elH4HRBFB7FP5kZ7QIpI0p5kZwJyhPvvwQE1ZSCy+wb7cUXpsQeD/58+km7QOn
pDzYydx4Nt5R58RuHgZbEy3I5cqEvjGfsZvp8zd0TgEVMQ0F6cb7p5IKZkFdAYsd
lgucvImYgB/Peq95KR21+Ysgee6+W0K31jRrQp37Aez1a+PkUZZE41nc5irHdzY2
zzfnXKwBA+SQNeT2qWojecsnHe8RQg42U5FQn7qUThNB4DievbQdvfv+2nqZM2go
nT2iI3vpG6BpsVODJQlu9nwZRoeZjWEJRCEOqPVdmbwWGl4Iqdn5+Eo7hvwbh1ax
3l0mYUz5Ue/wIU8s7bGIdG4JC8/fO5kj7WVnOPlAQRAoMgqzBs6RHW28FHxjXoZT
+41PBTo3j4O/3tOaFDLSvTeAqxvgHcsBISYXoNxmY1pA6twr/LO7AMYOAnXH+WzG
FxC4QonnoxRSqSqF4d5WORugzUIkUXlIOI82I3ZjYuV7VeFx0KMbPy5t9N1IAuC0
bJCcmx+BJIXSu96Huj8qcS4CSR0fpwT4uDd1oDOAUV0N90Wj78RQihbBkRqrpD7t
a+gHBEZEfHBhgL9QZC8zyAvkNiRNHG0PTOPeAA/BIaBceAfFSNoQ2h+kgCluuyev
MF85mQ3FJnQK7Ez6SVojDnTixMroVYn/Sqp+tsR1/U9WTg5mSaEsySw3YDME4nkT
fsvhzMPCAf9rRFVK7daoH6/BtSo2z1OWjBTjll1I7fd2hqTdvGeJ9SlYCYkTJ2Ks
qSBac425fJhdHmdHZlKq2iaPbc9TLnnWQ/n2fq7zw0kJzSvDky6iroPjURF/dzxu
jVobRgglxegop2vxiYrBLlGOI+QjB/yvbUyJ4BLlroTdIwskAJkvv1dj1y81XTVN
VdrRkYJN45p9AMDhPh46+O8ediS9V4gY3wc57xxRrV9/YpRJaVpLE+rICwW+WW3e
Uzw6GAs2XitXSOeuKETWKpVuSKXz20dIlXPVpUy9YtE7SzQiAIGPoyYKekYU6Rnf
XDJbr0PcaPQxk1I2VQmWOKabErkregji/n9ZeuZXS7QRbFb0TL1KU1GikyomgOT3
RSEkubjfo939YTDKGbyFVFlgnqflN3LoPJBjUV3pRwme5IVsElS05TpgmLjucRKw
OK2H0XVlHmDUvvvV1n+7YPuj7cixCpcNbnGfFwE129fK5ELQvRh5+eumHZSV2nMX
poY3WbzbnKomB/c9m33mGL6M92tw/i6XNFLcFYERs4r68EsIqSU/kuEvaSC2XyGx
D2nfZPVSH34r6JfBFeh6dJVT/VXuPljyssJJmn7aU3SYY0G+0ldnP/RTq+0ZiQno
1khIv5jgEfvfuOKCQO22D4h+Ka2ydVlW/Nw9htx5YMV09/H/R5aVxwS+hIJmYtEF
DDguwuHZn/Bk3cQP2N8uVe+yIaNs4Xi1GSqYAExNbLWqCNWMkS8/u7oGar6WA1a6
VRpellEuNMxjzQtACQ+akP8ThRlOwBeZGxjwGuDz7kPBlEL0whYgsrM19i5BQmCa
5gnOzqMnbkHeB2/BBxR/sjH88oKAyyIxxURTQpOL161Pa1pC4O45ox67+aYiSLVi
JzJUErueBcjKoLqvcdPf060tQkklLAq8CYpzT9HYc0CE0x6PRN2CWpS0MUniOZRs
4Hzvl3OO/3Q3X2UBMJy92nmsWMa/xBODx+47JL9qCIjR8e3+Mmn47XjTR94/XzMv
n2Iw+VGlZyVHrTtoMYXPwc1D8Y7IpPELKF4atUDFkelnIFzk5wIQjMza8/VKKyH1
Kvt9GhNez5NeUm6PmDnWS2G20xIx26h+iJ36qnTjQvnvkIQJloozoi2qUYk8nRlX
55jsXbFM3Z/bGFuMfRsGN0J3JO92uKu0Ei/6x2N2X2TuTjqaCwgRrw7auoqe/C1b
MxFVOXxi8Hy5cv9P8ago7WhNR3eUackqoKJnVtItEH4YC/tMpum8VqS7ynKLLME9
y7o+yZKvW+SwsMVIUVpuWAKDCyneWTPRPBdfivdLKqpFuLQRKaZ3rjK3cY4s3WPO
71LzEgb8t//uuD5DAw1CZhkqEk4Cc/8I/an4UKi0qKYJs1TDYFX4Dn8cMyrdzV9q
a8M3pl4uyMRq2toj26qlnqxIYrAiSj5ehF9XMZl3+vMwFM7TFEQCj3iTMKURTCbJ
t/apiqmHclr09yq10grg5KfKs+mtIBnfu1mAHzeaGNFss/olgkpTA+VrfAXglvTS
GtpokdaqbGEk4KLhwxjxmu944AYDQoSLKSeJJ3ImFrvrJv7e3K4qcJNdXh0aMMwN
YaHA3Q8J4cMnfdUFCx6J5Q9WAtXPHFrQco3sbuEwCycM9Bajc29Cg87kN1A/joQN
07TrGRNeZ5ktPfngJvjw8WXPOn7SbFs3QICqSUL24kYMg/CyyI30y4i7e6c0QA82
VsRDHAUpEuJiJU2+TicIhkokFviggIN77hv82gOv2cTWEB9YSn9MMR2Sfnc6c8Hc
CkEWpOuKwrdzozL8tJb5Xa4Lf2gu8b952HUmV60E+mPf/Y+8HzMhj9mG/0XOfoeg
S37rKYewcXIHUs0uY8a5azss++d+uTn0ihCaw7rhsVGBeRKVlvGyWLwiwjf6/E8q
ArZb11rM+D/RyP7r5DJ3wCignlKxXL5KwyBK0Eli4sne4rZsqPnuKnxoFKYAUmDo
aqRfX0ru8LbPiET/7gVMBmM6UTOd8EAPj3MNbXKrl+wFllyPmWNcJ6eaCf6MAOTQ
Pb4Ym3tH64YDNYhTJ916orPxyJaUKGj65cXJe9rWiuBqPwojbedqIsLegTNCFp0M
dKZl2jn8xfBUWTJIpk0haqZ2Z9SgcnSRqHJKeO0+bMslT5lNq9DRZk0rcXCsvIk7
JBBmrsQS1qQUF+1VL2XWvZ4wlnFI2ns6jUiBKcM6Q9cErmbsfQRkusJYdnGSO4OJ
cYXcONE3mxOCVFs2mLrAKBqA+JLZ8giojh3zyOtXjvBG/mfc4TtWJ8lJHzRKfJ7Q
MEHGuCAE7RaJBqU4aUpmpctdH2Nmr5hGQPMErzBdP1+Wq13+jE5p1fwEri+5xgzb
bz955W9qk58NoicoODhgXWXeNrQ9e/2AKJFHQr4o4SsCiQvKCH4pXnCMbfGy4Xph
yfpX4hSqg8yiyl2+gj8PKZpGVeSjYxJ5VTk2qdyIjRsIBD6n6QtxHQa9vwNtyWEV
MYilDzcqxNZ+JvQvxGF0nLWZ3KK+5dU+VmZhYUPyMsxFQnxfTq71EyZYXG4Cs1Or
gNw6al3uQPwzSqPfmDGI6NLr+iTGfbQAgfN02IDRbMDQF5KPNjTDPVERoWTZAHj6
JuCO1fa1i4bfkv8iw1f5E2BZOaUrzCNlWZsCnAKFZTrVyvJYs71zMzKh7m+4d9tE
nWLkCzl8LeyZzEzdfOumcSxFHvhlpwSs8HH/fPqS6wEzs49lXHMQXaausnwdBxuv
kKr4GDy1zxU2/xaniit2QtSqd+5pKAiMQKI2/nVLe+2Nq+xV7U7jV/9v8ivvE4vA
lUMpLlBb3K5AZ7oMC+BF7scGmlkzTDlkwN++ul01Q46nLHhWk9GL4rp33A1h4J4S
LciDMHkK/Qrjd5tupmuD0CNHp8Znn1kZO4rPcH232qaXSSiTad6OOfAWFaPW4F+e
e6lHKVv+nGX8Nige65FHsuzN9gl7jfo6NrAiT+hopov9d1noKH8YTG4QGowV/q5t
jX08x5QpPWDGZIyZ1eH7vrb22wyc5Ccco3Smr/7H4SDxAqv2mATevOGmelt+E7te
2KrzGBYH+RM3PeIrznhftnu7uQOdV8dMlEVNF6Ijf9im6qQWrY/8Gv6dLfj4+nnk
RtTND+wPsL4NTCgv3JpSwQlf1LNEqMZtWBIptC20u9jWG1x8WqA4fvT48B8VkHwl
73lBBCO+8o4RtS70DIRw3XJPxHWTBFlHui8/zgFYtkLtHSKHMpbcsAKpgGszrAdJ
YrIyf4ckJfsYXGe1qmhgiULim3P+kitbN1sT/r2sQVlpfyfxa9oD97Y7zEMlD/ix
sxKZ87d1d7qM9deaGDPAfFdprpMaPXlZxCMdNsj6fvEb0ozuGSLAVt8KNJ9a9bLF
cg+k9da34Uw1BfctY59tTzpeuRsueuOaAWYL64J27QNf1xk5gKUcrPn7IIASM2He
dZS0iDlY9maQk1hCXIE2w0T/4ZCoNwQdzZRArDZUWWZAiBPSCyrYUXYbmHmoprdd
Ejgs5IQe5MABkwBRbqGYGVm33sKitHq95HVU4CHWNQUAOs74pAV6YUkofAGOEAs+
YqKKZ2NUrLYZtWfEFmQJTaFS8X+ouJF1M3Bp+phswkf6QaNWgLUi1KDGcyLn8k0s
z2bZkDO0Zr2TWcOzVMnS70Aj409ZYWIUj120j4Ucwy28erzJeEO76pihr78OdGZp
kx0Ebf7s2q3x4eTsMUfwpgBk04P3nVZOLOugT305m8kbS2I4M+SQxz37UGFElCN7
Fsq2VuMLUMV7M+LFDWD4JJJ/06FoRCl+7UaGPtDWLA7oc/EXAiG1nkC60ApiA+Zt
Q2atnPb4H0IKOF45ZZD2uRyV+WGT8IAvale75+ioaUWNNSS6o+OGKHSjOYzcP38m
aJ6k6yvd8GPs+5fG/fbEFjVtIJPsgyIogmbjTw6bHESRiGka1c2+pLqt5uq+xykm
MIZuIR0rekF+bxXg4Q/uNg1X+G47zBZuONzG91cqs2ISVh5LSQvq2UZSEOIUht0C
5KTbdGNcmLZo5ULSSDzDdOAlbeVTaiX+XONdUAPFw/HLwqy3BHkvLYYeTQeaHxIS
0B5MHbXt92m8uZaaK1fiAHCbeCunRgpoO/9AT+cpz2HBrtP2q67WT6GDSF2GIySW
cJ04dyNpCdAu0veVer/NJj+SR10PuP8ZTTzUPaPDSd+CPhhKkyf5WVPcPYaTAABg
XlJnkA8bZ6H8V5lX9q12o+aCAvK2VLZ+3c3tzzGmMnTiIytVMZgClhYfcaweqDYj
uhxEcY3KX6V5WjsCC5yDfh/5eCDq+bB0QEbPK+mRt17W7b08seL25/7gRkUBuSzt
9I9LaVKdSnwdxipA35C/4xPri8DpecLegwXIG1qbx6FrfWdSI80hZ5WqHOReSjmS
Jn9zEi66OiQD6Rr6m8rCOwY1Na3MI1Op/+iPPW1vwGt4FB9kiXaRSaRRjV9PrfV+
ZYCaegqvE2JUorK4tU1lgrJdgbofa1uG73/+Fzlw3bTEVb8LYI8jIEgDNLxiymrW
ou8tV92GA51stjv/m35plA6TityOEUvsW/6LMNbGJLZvNGNKNClp8tI+d9tZKjfC
iLLb+Dsyass5yOhNnqO4v+cDWCdlilsjH6Ilft0wr0A4aVfR0kqEbmW4GL1riV3a
gEoBiLDuZd160QxRnt9241c9KvHklOjpuPjY/VUkCmROK7n70KtJ93TT/itb9uiJ
/fuzCvxJM4nJSHA4YdfeIzYPcdcj831RIiZpJ191OciFnLvUc8Vw4hTnKLFOdyiw
B1+Oz87h3s2TQcM56snFTq9oGHr140IrD/xRp0PnWnshK8iMkqPTTvminKqkKJ8C
sBEYvMFbRMgUYCWiLSIQaKSv3B2OsJGnm+jSJnfoVFhSwnY7IH1+nvbb59ywyd2E
Q/EyZ/2SDA1+BkOkbLBQRtzMXPBxLk3x2Zwj+uu9w+qEcfFpBcipN1pa5lOrHjG9
mZJar2uK1hTb/3us5a3oJS07SZCfZiCQU3yTMllSx37OSAA9X5+/UpaocWu8mrm9
hCBZ9iEwqeWxfK1FdsD4FqRvgRP8cPIKKQ4V86oqli7SjaZH3l3OjIwFadhUIEJk
7OHGsVktkuf0HJQWdxLtL1OwXJxkbE7WJBVky32ridAPItCFOsb8xXWRKpTHuvxy
9/YGn50SC9PYBDrmTaxPBCmqd0SqiuL11x/1mNTQWH2FmYusADersbAmJPeRhGB6
wS9TT8cLvVzaqDxaf4aKaVRX1OB+bmn+9kJ6DDgj8RnOB9qokKtUVFw24M/ElbgP
lfoRaF6fxoXpVaRAKLeAA/h+UxYYw/Q4s6PNU0d7guhajgnfEp5WksX6rpX8OmRS
Y6yRBFyBmWH3W2H/q19vIwbstCGruE+9F+GbKF/gcJq0b3dXPB2K95iMb2iMOdcx
BOo4zwCppo48TxGDzaVCGA7oOWSBmY5fS9QAcNxLoMppHT1fqZadnlsdM7CIHCGg
Dh/7pZLz7qWEpW/fatUvuYhMKzkduDJ8yk906AUsv4zLz2oHFQXU/JZc8T5Xeomr
sefQZ+aCfq1Bw/F6jbQ49uju7wU8giADMVFR4979vNLeJoiRMYCwqZ9NkPCRcLt/
ZPwWzMFOpkG1y7Gx5ZqpLmzUSu2/JCYjFUF5ce0CW+nTlIQOubmhV0/JeDnUcMFe
klQkxAVMj8rCr2S1sSo9H8rBSmt8vblnc/HZzI81zTkQ0ZHOgU57sPRM4RsGmVvF
BvV6x2luADYy66xzzuvuFb9LuarAeOu5cZzTzJt7LAps/FYEP2f/V5IFM4NyK9nu
9jBmmjoykNCZmHMBgX3N4FYKFLMdHjgHAcLurUKGpvLupWa29i4PXZKZEEWspw9v
4mR7lMgHVPl0cnhL4M1aOqvtbnhgrOhl57ZRtAwZ8+cBifCVfrYHbMD1vHpkwc/8
dudRG1QZWgnHv9VRpMUySOhcXBrD3HPnvaPxuh57bz0Z5pKRPpUM+sWL72d6uY17
tBtWSAI01jU5sZenUasjg+X+pOkOIe+5QZfA75fbnGUIllsNTlppXFkGYgYAU46T
eZm13Y4zXUWxEWAwfETWu3aYhE5MRgaPbjCd3FF4ZsYdq9lTs/9kxNTIYrwp8PDN
gW4U9FJ75mIx3JRDzpCjWHbcnOOpF+AiqIOPup5/VyxUml9dG82Dle+b0YoAqEy2
Rq8Og5bWcoW5oIj7d8d5pHIdYeK8GGIaquJjroN21LgNmUA2xv5fa1JU+FUjSIUZ
cWAM9IlxB4XATYdyEfUbUxXd9dXO11wQtwdDD29fK51fE4CNYAGi/JDf59emph+f
FAnMtmpvTPSGN1mntLvkWzPpo6ZIyJJrxvwN5uclNyMTItF2v7mO+9SZdiE3haBp
hg4IjV8RVzrhWg8Kt47J5O3Vce2DaV0X+vuatzFAhkmasLUQpWyU2DS+DwAs4SCr
m/PRvYcJSXoyJRsyv1BznziUNIobC3Uwkehk+r7XImnKIDhomueqScsb9N9AnspF
2KLUMb4xCJXVy/OpZlOGtR7zz2GQlOofuKayC4osWPvUJZr6VWMwI9aEiUqGUib1
F5CJ2brMlC6uo2kueazn/KmHkbdAvf7NHGt96tho0b9CS9IHurda1LwcvNTJnqHh
0W0s6HlYukbgR06TPWmAitLF1FBP6w4k3+jkS3oQ7pan4ArnPA2rZ8lCFiGtmm8i
oMTALrLmAhaOsiaIJjRqmMGAu0i17f6vIaTzar8skaJgdaQsoLeXovI2qKSJ7x3x
7j2QRhatIEfSALwUS0jiXzh8BBFARjoNOMlKwfGFXdBb9H/hA3Te+oGqL1fuOyvk
S1Y7trPoswEMjL15gvP0rOk3Kp4Vfz82E34lDY3JbN45YYOPwoGkyzfo7mZSjC02
xSOewM0szU1DeraxBa+cIN4fvU+rlxyaX6a7vrP6VJQvW+S6l/8T/0ksWzvCzKJZ
8TDQ5XzvPUbxKMDL9M/bJMaYwi2UaLdxOfCscu8RDZ91bbEtnKx0Ko3iZ+mRxQgq
1xm7iMd/ZjJIzRc75fH3YjUxzgzKCsBHT8gK1vsztmYnIz5MVmJCScB6o1oxeVFl
sqOYveg2wT+jIz3DBYhnxn81AaggiBhA44wG3WA0eQm1jyWH+0yS31LDTYTC1Ids
cXJd63MSpnaPsBoxGAOoJs95OjT9rMdmYuRaize3kb3jujd2e5MkIWZK1LDUxwlE
PZgdJJvx28w6nNNwJLAB+2PW5cFuQoATpvOpeijzAGnRKSy1Z7FbFcjBMSYvW/+i
sSYWkHHmGGu5FgBKYFePDODnTat2fNaT/KZdJF/1BMBB7F6TF7nLrI/Tz4xb/oi+
1ttgMaBD4cuClTr3Or6B4JJp4ItN0FQttuGZrogKTgavBCeULvf/E4r2HMGp352L
HFVQw6HMbpjEU0q8aKWbLc9tn9LASJkA6qacqdDiUb2GxLm/Rdf+hCeCUHA/pKLr
M8NJFNyLWNkur6YkuC4sRAd/MwYM7XIe1OKVULtUOiEt3Hgs43fNLMdYepNa4XwD
/E2lWREkWV1dWVuCy682uTYvdMcf/K+fg5Cq8HJC1zFTTvPfJI+b2qWXTsyjFdhe
wCbaMpuOtXLX3TUXnTyZCtdH9DnZlyq9R28K6bv5zU1jNyN2fJTY9Hm+OnaWNNOe
woAD/SWQWeg1gN3fltugklaEBNSmgIVSY8EQEdtFf5Y7XXXXE5PpFkXv9zW5xxPy
eLbOBQbgtCPXtmlhvnBeFVZ1HeG7sumux9tFQjPWGgeTVIdHhKxEe5b04hV+OJHI
GYwscIClraw99MbLveNssVkh8XR/btd7jgvBpNcx+xh3sIXMYkFRpzdSkKQMg9r/
eCXAW+nKIoY2uDn/I2YEHJhRPQ6NaEM3lB2JSRMRuVOWySrnFaNopBo6fIP6KsA5
9wAoU0opFz9zDzoQneuX69rUaBbU5Rc/C9gQf4vk0T4AdvbudtrqdTavSpyUwVSf
mU3RxqXRdC2s6JNVglQ884VN1N55QAUxsoM22YffiG7bo0R+oaIUabDzoe/EigJO
6BRWmRf1yfY/WQfaofAgobwo6r3ov0BnNExW02GUfz5kba/GIj+HJQqSJR3qHCq7
6iW0TKhDxbGdKybI/p71W9peYmB8PM3HJrtly8AUa3BleX8pebLEQSdhpoWTiUIr
F7iBSmf0PI6h3KuLjICfBBVI9JTei+udnyBmeCNj6CyTcxESAGpV/eL9oIon4NiA
pYy5d9DhPMp1Gp3a5oxqLkioe8xyaVXr8oCY7zOVPFFvViPPowUvopoAzSmUhOih
RQhauci4K7u9bvcrwTuxnODJrWHHdNvDh4dgcToBksSmUsk/hypfwn3WqHlnCXZd
0myEkDNUvQ7f1JIeORIeUIV6jC+tUSHuLvrwrTzOWUONnKSSNyBEcXVSgBAJPNt/
bgQfpP9oO9gAMqxXd/UPgF7/fhVIxgnYVK100FjZOpazFHQbQ+PyS2M9KQyFp9nT
U1N+zcmrmAJ2etwqH5KxbBCDtc1y0yiBMlO+pHwKryqpCrmRvocHuqJD22hI9KB/
8b3iQ6spzEK+KZ9Z8wD+Rm/iP8Z4r9QC1D7rM9Lmjnc/MgFPIxm1R3iOTb5tQXZc
qh/4QeCeTFwDuO7Qi8eD+1EMgo/34w1V526qDStepHAp93Ygz2AJbT2zQv09/2zb
1cGjni8kvBp0Hj1CgNs5RFBZFkkgRT47G9qcKZ2OtIdgp1uby1xMq8JzSOFSRzYp
SkP+9GJ3R65QcCbIRrGOTtZixxfj0EOQzUgJQNBe4Zj67ohUIlaCVB9GaT49jwcJ
ZjVAe1C7P8otUFpwbjogSqR0TKavTQn6Ax+2W2QAz/j3cHHCRofNorioFuxz0++b
YOqtjvwa31vaF/v973qiNILZFXjLzo0YxpaXd5tm3OzWEiOReZQkKUAL9EZOVCqB
DvF4CvzknLuRFxAGW/6n3rUhkBRZLbMX3gBbV/+12LqLrar4SZsK5Z63609pOG5L
6PQcMA9Ihtt1d/H+9MDh1Adq1aTy+0UdmLfh5QR6plUbo+RIfbnxtkF0IinKvgBi
OgxAgxZ1w/jlckZJg3xat1ysBqVeCAFMXhFbfr530YhEWf4g06CYTcrz2bCzmC34
PIOYsSIkX9UrcwkXL7i/N2PSHuMxVFpiJbcuTH4vIimY6sdR4grVAIoeovBwnpMD
ePM98h1UrereLTF8AbNMoD6TcbTmM78pmAvuqRxRkDQfGi/spxJFkQslABH9HM2/
VBVrjTBJpVPnJdpyPRG5RAfBIlLehgdvYv2T/V5DK7RKJTYMi+N2FmDZyq7G5Gcv
uV/Pm/7Bc9bmC8xGCyDPmiQZptHdEDdcnF+6KvxcxxcE4C171Gqrj7tCx0OJD2Lw
Cz+z8Tvuw5ZhYM/rGr6Mn0AV1ATYl2rHiyQABrZWFl+/mWoHiy2lLSSotHZpbnu9
rUtPw1xXVmNuSssX0bE3IRaXHwsO0bHvyua30r2zatPxZ/Za7yQI+CyTxmKOuzZB
fh1IYBHR7m6RFN7EJRWYAS7qDxSupncFxr40ovlMzsM6z3oiznEKSeUlAN0V4/Qn
BQH2kl7VArbRV71Y6Nw+ZTsmI1Q6tOWRvcOcSsIxFaued1+R/bB7z0AGIMbkwPFF
9YSizPp677jITUjP+tJdSQoneYs4zoLDirqJ+lK12rtd8rTV3dTJYNNqq2DpUeja
Vavnfcy49bGDSA/VoWrpw2UwE3R/t18rlBnaS/9OKGh8++v8LsBCvZ0PLNxJ3tLW
qoAQuOcT0+jNj0z41ZtsWGCHKIcBDzfDec9vGYX6FU8+uT/8nWVOGweVYoizyg6D
Z/Wg8TQMIv9YZIhlfGIL19+to48wfmDrBhq2L9kmZ93onFzmd9BEzXdwD+wdQafD
0V3XVo3gzQax5IqIqSaheznef2bgHfS5qCFBQWMcx5Dwf1eE22pqbYbr6FhmpTY8
O27LC3LhmsqivLUsc8xtUSR2VUnXgtZGKIOSceqEfIm5ot6Kqm0NOTrt4YLymMn8
sdSS2oMoOXFMFaVZcChZxVdxP6+iHkhAmR20c0a/hpkwcVKkBBphuWuGkllvkJC+
gkVHyrPYxBbuW0sRn1KhEdjl6lU92/uUa8/a2Zy+FBnNNluOsRyyQ/l2+NeqM5eg
zI2Y7UfcyKNll2622gX6uzbKUvkmaR3wUDFtLdnhWCTOC5hOJccWaYtdJOOtxSR8
k7twYH2NEV8jYq3x/oGEdEA5vrdqNDSPeYXf5EFFplrF4RcUqsANTo7aFqg9grDB
Tm0rL6lY9/ugv9BRBIe4UVTx8XlLU8ahmMwfFc5tDnQSrTiJFzFq/EQM1kCg638V
w3sVntAG1Qm+dr7w372n6GDs5s91hn7GESXgfrgJhHSc38d9Q4r9knRZDplga5m1
UHgiD15nkCGTT9D1tQmCd4s3pJin9O/S4WQllL/PIHqPP5CBfa8eRTI4DOKzhehX
sbb3KiTb6sKsemoqGG4qNYgUBXVFzei6dW/a613whxGQc2pr6QLSbPWf8NNUAc31
6ko5QzM3Nn5/ju0JDnI0s0ErT0oR1VB34zJw3a6d4zmdFP1kyI1N6s/VYO2Eh5cY
hfca2c2Oz62o9HYYy1o8vF3yQ515lWlm8gsfhWBuL/iqyFwdKAoTcg3NuEtNccPZ
F9p1mYK60tMIcLs439pnqxJgtFXhwz8vS6869ypw41e/7hozvhTp3rZv5umdbWK7
fOA03ERHK9VYDDNdbPYBSwDZUQZ8Ki1q4U+O+w9V+VXo2lMAZZ+zzxznf6dJZX0m
A13aiZmaeCxMYRqvR85DLQEqJ9t0HQA7uoKQIkARS29aMsZG6iHxQ8dI8jCXK4Ld
nf8jCluaupEkAkzyEqNZ+LaRXhZ6P3PVH7qvM7G7CSXXqRqNOeR9Ui51PCFWVs2W
cbxSKsfjQthlqWWHGprBxPr/VGItcycVx+F+8uLq1oThpJq+m89JgkRSmD+0hTrJ
5o46fyD7bbuK4MS5S+rWoIfWIxttEUnMIEDrDFNLNTx1DukdoL+0zkFrhm0QpQEJ
FSnvsJmqfOrwkgyIAUrO540Sg3XTwIPZeXDvG+++m+6ERkYfh0c6NNLJxhPP+g3I
RZT2yamz7DNzXOFsrpZ+Dw6pk2QAvG5OCH3djSb8+fcCI+x6H2R3ZRALNKTfpEr4
+1jwwWuBK6lA2LB8GXd5/oOqWbs3eBjSEurvck6HvBLbbXT8y0uL0avBnMdYxv/y
EQsIExvCJENiAKZwokHetLHoh6XNadtj44w1AOiHEuMglqVKdd8oGJYbxfu6ZTnu
xZ8vfy0s0nxDkFabljFOz6wd5MZKS4Wh0nekgN3AbCi3C/KeuNgKt0o2m08JjmQd
eFawdjILBn5u9znRY14JhFaG/ApZsVpz6dOq1LM/HmZQsa4WoTrKDeZK0qagDmZo
iVYtdN6Sfl1DGeVtAdeDlobmTiFOiH7G4Y98GCZo7ETgpBS9AGRyekJwdKhLawcj
RvHAzEw0w8fLDMf4BeaNItXSlFsuot8QfrgAB6OWLmo+ktXpwAveBHk63fVQIx8s
cNRj99MoGZWmm2wRAl06ok3kk0WQ7q1gv+qbbpGjp0zCWQsZKYfbHMshWW4oURcJ
5z2d4QDNBP2yy3tbgLfq2v0kS+cHrOKXJ22woQlC2WNDwuGw9M4CVMWR6pOZA58J
PdXoCYc3yMhu0EDao0CO1mflxTeX5YCmCZoOn3JzMYz+AN9Y7WkVVWzNYcgm9udp
WFmLUaswbBhuaRHxqpK9w/654Mhqx2dUG6jCHcz1Iqhuodzrth6BqJVr6Hru0dWD
2MbdUkBGe42AR8h46AtwZPLk8FPaaPmawjA6zNBXAkY0f+rlGcugRVCcB7wfLMae
wVWfXHi8MrIVvLVTt5ZvNYumpadbP1U22ifiOnKdi7rPDE9bvIn2lYFeduFg4Pa+
5xo7iEan2m/BFD2wMJB7pKi/ASi7JsRMEDg9TSniYii5nw803/utTFqiouTCtdWm
O8eZQrBKhjPGDLoLdQUWcnfLpuJz5IOI61YIUfa9FMXh6Y8lt1yLbBYZkZqS+i0Q
29p1hFQ57bHn/iMvFNmqS4PW3Qxuu3F458rgy5SpNSaKcSDdItHQ86Ic0+MAcE0V
5Abix4Ln92NohENePLLQJUWTcSuS+RkC3cZbBpw2aaAMAzh+Y89eD1KHu9LRS1Cl
ZYf4g86RpNyZF7z35LajyCsUXbwhRdMqEi1i4DzgUy+G2QeOjfllqxzsnwfbBe/f
ar4wXivbNsAFhzcv/w8/D8yJYmVBakD7SWR0U2u6izvhUnIgzAKzFaQtfKSLvRe2
brf+GLgrKP4vAgAnThmi0KVepvAm1hzc29nI2i/vRX9/e0V0YNZ/vl1WrasTONz6
wdD/mdTvq9PbUajLVu/1+2VivJzMBLgDaqsxT5X/3r8k+hmzNkqPb2tz105byhQT
QSuhHssdVRBHvZIPsJBd7yPKmxbm6ik4mrP51rPQ1hfQ5SxaKlKwMmQojaqu3DGX
WjEePbhooFZmgMYAbgaa0CPnTVxmy6et1bcD3j4/mNK02FnDjQfyRcII9CxLRQ+J
wmm2jZ2NlEbnKWTec8xlc/yc7HB2+MOXXNheI5Ab5024+qtZvDjcQjyh1QkUwsa2
mYSG/9WzlsAQGb5Q8aUb7lfdyyw7fLWHjHJpQ4+NMHmxb2g3L49FE+ob+HvJD00i
4DHu4J7lWiSTN1E2aPo8N3ZAVP2R5kHWtDcQgeup2KlU5XR5A4AdTQmvEpAzJ/gB
eZuMNe3Q41cPkobcfCnOVzB7NoGBrzTzcQ214PRwGzCkoeb9nIlwgyfZsUuP5tyU
NND4i5XZw5C+bpy7su7u7fz5IgGFmiaRmZDdhoRbX8r8wRiByumb/ysTGNdpsXdD
aWcBHsBYCxyfeAN/2JPNY8LD/eWsFzVFfrmuB3HPou0nYhB4ahlwODWVtOvAuIEu
JdsnR4ebEy0Tn3/jyG3s6OXsNfHsmuavh4ghzJ4FnY/svXztGkaLaptyequ7jzKX
Cz0b/CwG5UQplGKfgtqZTRn2UPS1zEQh2xVUbeGdE4KT5IuU4oWpbDBFYpvrYSwd
wexZwwN6xVZ8a4sDpmdD0SsPJjevzi0wURx/JZ2NA2DlfVlU+SP8qmn2a7lLMbum
FvDREwO2Rfa/RwBkYsjmMxyCBLn4kDL4IiCHmSA0vJnQVVDGirTmexVWFFD8MrRc
wwoKG1J57K4QMSgv6agwZ4i5RPJYSZfIjEUbBDKpVmun8d3NI72RmO1m3QQuF0U6
LOCXWmlBOdQCSdL03qIcCf7fxvRlyBY7ecbejDzE9YZDqHo6KrZRlke4Goig2Vuw
Z6yETe7OxzhY15TBMz3BUJDjot8bE7SWDudFlsohBzKR4G5X5xDfuLeHCZx2tsUF
hAxWpCJb+t+4ikXS1+Z1hVWB4JSd5KUUFwbMur04fd4YSk1IO7/0ocy5wf3oF23R
BLgO6IhFoX0QLleFp8T9UL1mCng+69FOz1SkJmyo0QIPjmfIOnjiKdbATBUs46bN
OccjqT/2N21C3bApDRFEqjCFCeEuTnxDO4fQ/6y8PqJl7dssBrzMEDZmEygfrN68
tGSHv5NCIz4iZYWUrG5fOpMHVvE0sXHv6KqPFbI532e2EP7YKpxWNc7XDF0c14q0
4jNSi9kJxdibycd2hngkgzP95GaTgJhtvYVWkgxRxlJSMrPXVDApmBLpZ6q+Jg3I
QjQhVJ+zbA0CLY6Y0Mdexb9bjjDIWRtB8h1+JZxK+TOlio2hPuV1wPWqEMbZrVhY
Mx089fdDXgBMev65eoPYMqaUdV4XEqAQs2ndjXuPVavInWYe/196tWpnoFWv+KS5
DHq4+Fu5YffG4Rud6Pbd5W+N96BOIdWmIhqXl81cA0teD0WX7K7BKEwBw1wFzGlD
pZsZf0Xp9a5lNb6wdwIgtoOQg50d8CRz5rccANEQFEI9ssj0K1tFeazrFI5gD1jr
w9rcwTC9b2yVvR/z64NZWfMLP1sL+jiwlPk1lalUwc4fAgdLXjUlyXSynuHWLgYX
q4VpMctWp0+OJ/AUXHpQcFKZQWbz1GKtIlkd8EAxpiOVqCo92jxjFz4JLcDTjW5o
VA3dIfgpZrGdwk0YCWtvgEEH2ONHAIvpJXigJ/V106MUP3cUV4BVg9w8TKbH9hRa
0s1V6XCM0Hw/vnxZ0lvje9bsXx62a+PplhwZgslTlN4xR8etu9e8K6Tofuafvm24
z4L1oUEZ/bgmbDHl8oKvfrgwH91VUDy3KI8lqGSPiO6Wqp3HR8mz7mDJFHXzMKB1
sTWsvbnrYgHgeuLjnI6csabl7C2XVdPV8PVWmnXRFstVnywgmD2iVtloljjZesP0
jo/sWKxkJz0LKcXnjsWRtO1KTpdsCOWIBpQX2mEI4Zu60MWNgqycfb29bJS7t2lT
V91lij0O2xEgn+GBQqgy6kA7Ga9KfuALEFEJus72BwK259rKlAQJwkmjRGzvueQP
k0Hb/FinsI/6Cnr6uXY/fwUb3WKJN5fHHNswRNpUBlFpeh9wW2JopfO9/lzEGmGL
R3JbA71irsM8Me68AWHuLaJVzTH+Wnd+RwHcAVQQo8bW7HJbMa07IPdQVqsvNA53
ACBJQxVWHS8+8dlwUsHD+DmzQ9Jtb/N8LsRHDjwJ7LxsKTcM4wX7IttH2pW7rrYo
BWhoJw6Kh/eoGko7OMfI0SRyu4wx8Klc0h0MtHb0462X+AKYSHXqWi2kuHSoigII
3+VO8VfYhubbFb+1fNm+3TC+GXcUWncz6m/8HOsFO0Y+mNYaAeuwxSKnBjHMaQ+7
mdfwbHWu8VGb56164pdQ6dEHUnrkNwF2UV2I1tjZNbHO0t1d1RZwlq+n24UAJt7Z
BTRKaI8emYOw2gCibvmAcVfymRnO5RK7gudkk7XlsYvNzJfsQDyAJ2vIUTEnNFqK
GJx5+mONyff0CEIRtpsshl5k8PG365XmaDeuLhOi5XvbqIrvGfA52m6XmcVhlhtt
7V16WYOTx1/rE1dpJNs+dTf7wHcO6fHlb1ACnWJ52LXmHvS74fKReClnBxZ374ZC
D0NeRNRWZsA/eF4nPlTkrmb38QnxbSJ12x4iNuIkKPnnRX6ueo3g/FTlsPIyHBNr
u6we5BVyp1o+SN+S1liImJEQ/uGNTRqsJ+tkJjUHHKfVlNMdMg8zBEhgKVGkv3Ip
F4xpUCi1+oMqTYFlYSCD3SMlut46hwiqLAY8b/dba4bggIU94RcjOUTDdJezuV6T
VvEz0Kbhr54Z0hWWKYBbuXIvTzLnWODiSZUmgUyHvIYz9a4CG0ixgtgL6u1s5jPD
3h+XLaJpM/w8xDaQTnWzMYrb2kK79S6WppfQAwZ6S68IRAKy2mtqmZId2o4xLSMN
NPZLRvUENKXpOEC8tHUlUu5612RiYs6CphGrEX9/mIqVCkcW5R8nBArAGk2zjzJz
nSjZjdSe/P/c2L793KsTeBg3Ad/ku7cRu4TyUHoJ5aT9w0bn5KDRpAtjh6bWgA4u
G5hqYoGzxo1QpjUhssXcYfGDv/fXz5UENM4Ty0fwEo+e0smj3wp5ldgnoRngF0L9
FoudWj9GOxBOMJT9DZaxK6O9l4IOWOsHKAm9m8RxTENNL1/1fr0t3rco+rUyT04l
vrNOvuCNC3wW1ANieWskHd8YemwjGTsek93Rm5Oj26M8obhKatHaeaJIfwG4FO4O
RwkHkBZ4AiemCws/h3d3ptTe6ZK7DENLc62UnO50/DpBN7Q20JEP22shP508Oui+
DXmAU+/CrBXUXILPDeUCF9UVwQaMWhVw4tuTGVC3lbwDw/Nr4onVFe3gkgXzjYp/
Uy28/AFcRO4KZAnonS6hEowqOvqtnMee5GppPQVyNbqF/CjYzKTtuVNGbED+aYg3
b/9uBK9HHeBfRuAAeKoL/pdkCk1jQsMY54Y5Hf9IQHhE3rWwsR2Bb36n6Tsm+3vb
aBBEzTDIVkX735IkGtuPnAnFmj+RhH30YWVZPWPeGwlQzGrOSEju/dN8RIQMrdj9
tkiSo6OvCg7xK3+/gPfHpycQVUH8zL+497m6VYYmV+dUX0jl44RV82S7A3tCJWhh
zPiNAVqA0vUWH/FsXngVmGlDSP0GEebmiC7+D/2XuqPIS/hQb0Fwp99cMDIzVJEr
NQ7RDgmoP3rp8w8SCfAI3/JMoY6zNkGXUbuyS/cbUo2dMH0gKc8ylRy1/v1LK8L9
pp4OWS0Z+aRHcfOKf84GrgYm62M25tskKy0D/BusSvcBsoontOE82IGGDaRIxm2n
tMs+69sxUyReCSkO320C1L3eVLsB92M4RsM3toeY475Z7w+/4ejvpilcug/zbJvv
rph/WWLT97u+LgIwQIJoHm/82Nehw/b6bgWR5/PCMThkiy5Is5x+Jms5pw01m6tR
jkWTlY54Oi3UqgytAUo6jJs+m8ANlf6sxldZDNd71cZpxOrJDJogPfuouP4rQ0Yj
RGok/By/MUZCzZDVfWv6F2D8PfemOr2GY21UbRVvunuDeLFTdETmSTwtdRmsB1G1
T7WT7wdq++uA48tPswwoKamCIZxEh4SmcU0r2NGdMB3MnYZpqCmd0DohDiW65tPC
dVi2iiF4pQKUTxnGp40R35JUE1rP4pYJgu2QcR/tXFqIshB6a+RCRy4xLiLGLqJk
o4vlx8NW6C15JZ2+6ETRRnWQ4vre3K14IIklJRaDPSe4qXfFOBLeLCcPStc6/wY6
PTir8rVbykSRusjJWMvCUYcw/2ssof66jAmqGiNYROGDdpzwaNWt97G2dgc+5yBs
TU1oYOXg562XuPHA238j+AIXLNkYogI1IE5vp6qgWZWalbbOHR6U1sRs1d5+Yg4B
mjmuvQvxw0j1FZjnNov13RcUX5HUKtxMNY3MQMkkA6Ive4LE+MC9QMrofneP/Iim
LrB4W5qjSkrU2EC9EwFqBcRzbfR14hy1xfyT+fH01pEbJtTdaidPDmtanc1muf4Y
2x+nMe9PWGQZJ475b8vtTVego0YyuQBl/2XERqmhvAXrn8iiOYgzRapFQJgNC5NU
P9vYHYLpcIsuDAZybX7d3WR/3tCJJSwXtupZpqk6yUnVxMb7TEWjW6qRogzSJ5/5
6CMKHVWbm97fxOwQCCAIglYZ3xg2IQd0VUYr+J0CEwyANbuwG1XCsxvSB6R1dRzA
ofP18y4A1y3ojsjeKwhSvVZBPJceHLUohMPFwiLQbpWQ4MR8AIssZ9k24TgZOnpO
NYffCogr/7DEM+j2Wqd1EHwd3D2+UXp+tkMyronAie3rwZn1I3i4M3DrbrzRkLzI
VC8oZ6NwnVu/CWwLWwtVRrk1RjlRil8bCoSHl7QUXwEBtD5SUJFC4yDiCtJPpalz
ze6pQNpddOEMxB0rz8W6ZOoVMeUn5/AHmZckEJH2YzyWhp3HVP+9+EtNX3qh0kjK
1Oc5UqpKMQH4ObECK8871BQb1VAtXzrFxppM44U7dIM86eQA9hfDZqt0CT5p2kv3
aX9px1WKXWOrVPqtWj3uo4iGP5o6AM6y9q8dXDCYaP8alvz07PCyQfKpMG8mQLyA
2QypdxVOrg6Ofp1RNUeklm3d6jhFDMRkK/rkj/b3TpA04GQFxh0AYd0gN3FCPuzc
bhJapmbIjyT6rSidtAgIkTBv5w3uMGE2qDKRxxL2baOTC2QRqnmmARnPW5argM6n
gztCPjUSZ2kNiQvNjUMxKV73grhVz3yoo/HYfcbceXeQOuDRHuB9aqp9A6gXTxzI
w7TTftezG/Fp6GfuTjd06dxC7lghJtpHeDGBAlL6SYIaswztP7xvq1jpvvnRsqBW
BT0vHOkl2fB6zmXI0k7D8uS0UJ4nLLLA2XpaaP18ris3h6V1Ws7uR92iJwg9CgeK
lt7MTuQ427mMhBQeC9UtX0elo8to0sIFHhokZ7hbd2BxEPbQDV3zXK+Annxvj2zS
KAxyVnQ2F/bYvQEG1ECgIRE1aTuBjdihNrlYALrePzzY9rXqXs8arVSnKi/roC+F
mW9E7zvbghy+dRYOgeCGP5TPcVjvKV3KKOT3gDcty6ocRWHjuORU3SAYNUucszn7
GR7LBUJDXupS+0eAKLlwFGHAzhpKWQAUo6YxYHdKX9IiPyh3n8zi38jk8fKv6RKt
iA6mPvB0l26I3hDUPSSWwqj1VYUmYMwJJmopxydSKAJ3MkbPEKOXT7Ugqgx4I1aV
QEKqy6Knna6DAe5S32wEg63OzaE6eN0Pbn+qt4gllmQD0pLPPHvHs0KxpVDNUQk3
/sfT6X2VfyZYasw4kMm1xXOEEWbpwCIL6P1emSmJKpW4P5DzwqAudFa8lHTYwfqa
muea0MIcZQDfU5UpYhINybXXN5HU4DPTPAa2R2pUlnSxjII8xtap3x58H/8xIU/8
C/iPhlPExMNJ0eC2sp3t+f6k8pKYfhjc8AMYr28qKnlyj0QvCO52qrCV2YhnGdUa
RZAVua8hiEtIyXP0G5QAp05cg0vGNu8Wtl48Gm+uQtdGrLJ/XnDgfIe/Sv4Di4ky
eHFd8EgvPB93M+YuJ47CrLddTOivugKnvIiYKPLln2vGHw85EyeMuHBGVLSYFZlP
vNGf9I+QjKXxx04DqfnEViSu0r3xwc+Z7pvAN0PnkrXfUqOeZ9ZIMSMtHePQcAzE
vEMD0LrafG4Mz7gMK1Ino9F5xDmhY4iv9PJKZK7J9itsGPXXlNqIhlPUSpwlJPGI
Wgrc1nEQfYBV+2I+v6rAmII3pG/2eQrjhISRzTtLTS2E4nXSY4CrLVuosWnZTTAi
WSd0h6F7+TYQbsl6Gy4rAB9NDQz7bv85MXsrMx8zCIN5CYugRE3cyFm5AtaXhi3t
2msjmg246ISTOsGk+M+Z4kWgMr5UnHrcP8nW/d4Wm2suUSS6YqxO6Bq6uLs9PaXX
50VM5mVXG70myBy8J1J2hzCu8gaeUHQLGy/WCrUooHiSOvxK/l+/pg5z6leaO26w
J1pypprm61LpaJmmqmdYq/tNyHuMcF1fT4+0mLPVGJwSLeQav7YYSHGk5mXAC+al
4Uy2kC6SP0xG4gGJR8I63Yg4aJKs799D9BW16f9RpwxXg4cJY1QNp1uNfxYD/QdN
2ncGM8mTiYmB1DWx6FpPeKhUID+u6jCxFUViYQEfHUuRzpV8VRD774ZQrB3GPTFJ
Ca7GgU1+i2MjZAFvYnu1jhims7lpfOFFTWUNOquYo1GvParXvOPDL9XUfFUSiaZP
aPk5ZgGUTaO+BgzDwG/BuA1wgGCvh2kgrfeSVTi6+Yn1m8fwuVSErChp4RCdZo7Q
+R3VoY7hbG1Hyda9xaTV7Dh56P/Fcg61FjNQBK+YA4ObgV9D1YyptDZda+kvd7tJ
kjV0jdUPDvhwqQrx/0ClMQBhLLcMQpR1aLTMv1/47Y0+s5r9n0Jh8THz6KBFx+em
2ER7AjxZmTheRpSg/bc9sh7Xib+1469ZuEpJYF3pcYUTzabFPDqeDU+bB+mZAgIG
pkOmbf5teLtnVqg0TsSFHB0nXDuWNjevuws4LRR3Jk0WQjzMKkV/xaslh7qzNeVv
y0bO1cdG1+H04Mk8CYgklWlrKyaTRlv185C/Pu1fpJ3HmPFaUB8lZYQsVdSMuAwo
bYM4AVclHztbNA4ooMvLU/H4uqp9VmeSO0oHNrps/WHJFV9tdYtsVF+WkHxKlu4E
Rqb/la2fBUOtXxSXPPuYI7pf56xy31bDWwVaklgIe3P3ygRS7Eq90JUvianxLiR1
qeWcKo7GKSJE9Cl3lPpLmIGRBecWniNtos5Kil7rvxq40JpYudXnY7lM/PriO31W
bFBWfFlnlygngoaheT4PPemlmJUyJ8qS6ITk6vrUQpaS3H7SfkSHKM8XHDZ30Gxs
W9cdCS+J5d3St1Pn7ltEYJN8Nip7g1BQtdj+fL/aTaYoyB503tRZwxGkvF8dQEuc
joX/BLMVSs3e/Rq7fWlyaJdu5r6H9pNljALEC0a1buF3U0WwFX8ECxr2YM1VU/2C
nggisXgI9A5B4pGnUZhf9hqO3po6R+B/4pIyVYoX8uOrQ0JS8GmXT7rjp/rcMl5a
6jbOGVeR0PkUkXjvaKIvhE5+sRgXG063BBRb8QVbhlFMxPvKLm6joEnK9u3ylvBU
xykyTfdsu3f4zCCIhAQxYpXndB4gXb6qw9G2oMrO9zlTV1BwpJ1NqLKCKAnhcpPP
Aw73SUVqmUv6tvn55/NrSzTue/WcrVipw4KWk99H4977B5/E65/RRL6z0gkJQO/9
znv4eAWE3+3P/z81i1Kdbb3KaBvuvXR5g1jtsRMSNU0DnLcv8mD6cCxiDLOMSx8X
8yRAlubak1IE6hWB5E3UUVI43dpcQ94EVmwyUmvAxdveIq0aVF5u1mK9hX/Xz5PT
taGQ5c3kK7lxTwmMZwuSOHUAklHZ4plUk7B5DEklEKgAbhubpL1sv67QxsVxCs1E
ohNQoTKyTIaYacWi6Nf0IFinZPtUgQbHbAhO/bKi1zFcNC1nU34yM+UbwrPXliXH
xxV8+XITnl5c2nGU6ghBXsTnbqzccrJd9Xiltatlcq2lCDnW/fssXhuiEAvZR1iX
Kifq/xJ0VWMV4SoohWpk3CwQ+XeaJUCNKcWGG22H7RvYWkel3j6ldPRiRPbis9KF
SV8cz2qrbtMWPNQdtz+shiKf/vGrC80pbO8iRbmqF3E6zX06VgyLW2gBGfm1V6op
h/gPIXZwm6hJ3wzqkWK9VpVYbXTe2ktBFCogU/dhJcx4P+oIGzUZuB/YAvj/rH1W
u3oeDyeZtjXzVy6eg0ygAINNv6SF+7Ya//ZnsnjQjiG4kXPEtF1gfU4S9vQrj14J
Yn8usanozDV7+wemjPav2lzt4BisZjyM5uhfoQuUFM7CCFhShhUTZ7QHfL3ZJHIi
RfRzADEwUWCTipAoQ6FijUwmMDqxGtjv0frVprAJnVOSw8i7P+OGxl8aHpJcsx3N
1zq+BKGfh6LnGo6RNUmoQNHPyFQZNM9lVBHg9zFynB3pMtwNECY4WeNZoP5Lh9Su
V9t6KJYOGMCn/mvCUq9H62pQ9BxXOrAfBB+vN7kid0TY2x5vg42VX+5DnWra1heh
xbmgjlDko+1ywOvsRjhQPC+fQUgPxvKGcNGOUZAuo7Y3VQ2Y8aS0sJJgbE6CS0sl
VqfFk7Y6734ze2u5JOnnb+8nBQUzdAnhKEbgpkquNigrvGSh+KYDFaOZdzcro6UC
R2xcHalKpw+Xw7CXas01QlzUu+p8yFF5JhA7rScUaPhtVAKRdruQpuMBCG+nS5U4
DqDwXH0iRvgFVSe0c4vu8q8ZiQswZlhMPmYWosZWCLSUK2UVanbU/fCR5MW/MF10
b5Rcg48op9dFPVCHr6JEZjv2AKJvlUY/DRiypStlfXakoq5g6LBjwUadhNNDNalu
uOu5aLPjdCj33kiWaKwbz+M57LapSWJlIRqlosIjKD4uPFje2lSo2HyVKCBvVFam
dMGpQ/V0hTy0E0kMsZH/q4ldBuUpLWMqJl3n195dVHbHPYSzksgGZyB04g7ZlLAE
JLpdPlv8S1LnBi1wfocsqyONvZ54lOOm7mRocCNidaSEJZ/CBA4nGOkBJDQBFVsI
8akmR/oDMsnGofiJv6dFm8tTXBljnZ7vZyRzdYOZ5YjO6aZfN2aooyESm9ZibpWP
tlDNEZFZMSacBn4L6nkPIPLKpokACa1ICWzHiTJWRZDeE5D4lzdHeXN+n4ZDgkCL
6EhUDykNpOJyoX3nq+uF5ZQOhcek+YUlPqRW1E8h3OrSfDi6UI5T0Xh7C2l+ei+d
hH+s1gbSgzrQ9TeXN0suuAipv76v0MK7HaXJu8XJXQscrWdYos9ENWt0jFzvXt2h
rI1AMIST9RGf/zd7FObNd2PkFIat8pa/Z6IbsGxDdvxKt7vv6jSETzmn/Fv7ifVc
JD60y7D194wzADizd1qKu9JSK07CQJmrJO0lsenM1M7lLjHK8y8N9/Qy6+hfo5Ju
375KtaU2t+vLVjvKJ6cPG9wc+daTEfqh+G5tpTv95Fw04zxtDi0nG9apQIV7lqw/
P3qRhpzdyVhMdz/EkjfwdhrNOW9Q/AbmF11yuENsEuuyW90LypFfGiU2GDfzFvOr
sU+yNcYVCi23LQeloVwxsj+n+MEpwtewMHmYXY0BMUADuL/xYPttV6V12gqnDkWr
ClnNWA0cVQCDm5x+PWrEGugrdag9Aw4EzKiGQUpQPgCKODv+tos6Ja/8nVWMZ4lY
jaoB9ZNnAQQJ0idDslydzdniwGnniVFMCl99pEGxjdhKpZs9vggHNVZWvWBQcADf
OcANmrkL+CbLMy6XQugcIZyHI8Heu+DoO4562vAnB5iyHzEWoYmaZKZiutUPB8At
9NyjDQibfFKGQ/U1plETcf4mdgBR92LKU/lta4FGGNcPweB/5ystrhSUiN762bWW
8OzduCldV1RMu8B6L9JSHz47qBvRgYFiZIzUnat04I62XxFPxXZvSG/C+RLnQzEX
77SEkte1lB+UDh4n3sQP3oq+qN4rY0fEo1rC2+xVjL43/a5aOYcg8b7wTq4zeamf
B1wQpa5hGlQqDh9Fwj9QQG/35ZddRpvVM2KTv+brov1e5Rvsh4s7i6A+H5qUEZ5P
Zy2VSMvlVv6r1MBwlqprEKyEVUqfJekxj/5N0iwOgQgpjW/GB+vjeWnix+BdgcxG
F24tId4U7S5VaOyZFR8Ddobg4CKF8kAVHJR6UuO7Gv6kJRXAAhW46j/LB2ePgsOW
Z6O7zSJP9SFdIphvqvCjA1MeC90LHiCV1a2Kn2sSZAYqM6oPYMdU3bUF8eUZWVFo
infwHBy24KZh9SJia8sZjFdCrSC1ZqtnfPp7S9oN1DwjV0wH0mqcyVhcsRPCmyqm
LC9TBw7kU82F1uCXnp1Gg0EaKMyMTCQCDeqOlETtJDAB4V+ckVPAZZy/kUBTjfMt
t+NrK3fESSIriR4jXSm29n5F+93NhokCM274OL+cxfxyaC936VlEdL/5S2XVNbiV
Mvws44dwNcNeKAL16oouB5VOjQFRUmIA02ME4x6E2AFNKtabE/vLPeCbh+Ti0zCU
ksShgtL+GgmB4B2S2fmW74U4+0wJ96J52c6ecjWhsQ2dvRi11mRtZbw8ZPdooVgn
kpZQmg4XBVbpLJHr8bFeg6NP568MVlqwrBZ8TnkZS1HrWD1pjYhF8B+yylBqMrag
bW2GYi7nNYbVjIGTf62GTlodRtlw2BJBamvtCwmhnWREnPU8oHA4qZrP0/TzYsDM
6mdlOfDIn40b7jldmytWrXPCWUoJuxP0KiBe8oDmRuYEgI3YPRy/fHq8nmHVlF2m
+S+vXRplSzgu95Vrf6zgvhPCRbC5O7/EjVN9Sxspda9wY73zC+vXdruQ2CIsSdsp
DSLKGhtun8GbdCntB2UATK7IAmO9Ea4/GmkEiTLD3BSNRmhrCBbdpZKC3uky6Pk7
DLvXbZqQ9+Yup/ZtSZxfbhV5f8qEXE6F1PaVbn2ZmnH9T0d0+0A6QcmGRlATj5L9
YqMSI/bqoSExJU681P+1gFXNu2f2HZW5IKMFQKjXWCPWQQ+E5bhaLof0CO+w6Bg1
SDiiVTrEN3oLQfAOwRQOfGa68hBx7MOpG3hJGmuvgo7ZB92z8uAf2grSfO0+X9Hl
QwtuIs9ga1JiLLgWmEp6AtV6mN5ECGaxNXtIYasOMNOgCFEhx1Ev3i91Mm041rIo
FsxG9B73P9e5s1YNY85gvBOKZjbWL2Ql1+TGwmc2UO4zj56BiBNK4EbTbYVQAPsy
eVMVJ3YMMWFHw1dDYddSbfhJb7fsRMkPYLxOSso2hjSCwtzVE/t5RUy1pu6J/dYP
iOIksLN9JD5Bu/9XlvLXiXQFuHDh52ki/8X26+vTCgjrLRGxDSQ5Yznvrm2BinC1
30Z4scPCaJTJ4LWM9EnMoqSJbfpiCn9VPcEmluKDyhlI/FQ0Agz3MvifJ1mpTdWr
SeZRgQcI/ACsNO57Mlb3Ficd1ukKLQeBAfxPNf3x1qgV76k7SRwrWOp1l43ZW7cb
76hbtmNZ/biGlIUZ73dVFbIQgZFuImT0BoGJlVjTDoKKmGeDiE9awoUwrEleI14R
nLygReTsRS48lOMNsrJl6+R/oPw4DB132Ar4S6LV3UmtqlxWX+f6JToAGwRP5Dnr
gRa9I6IyDXZXVWlVgscnde9t/dy/7xKL3Yt8jN9iuuIV/nwU17FpEvgoqn+2fBXg
IGjBG6R/1ts2AVZg1feu7hbFBCujc0bhawCizdEZSHsg9RTfbrtjvDvw0SdiikaU
7Tlm5h5m/KCLh/dQzr2TzgKeJhh0lRjR+KKnFqBkxpD3XhW6fyxcSK2Qvu0ITuqt
Yixo6X81jgjx0wtdX8ht7dXaRTEbwL5GLY85BkwpexVED9yYezsq7Mzw/ih493pe
JRaItKyKnkXembKQ0B4+SzE/0sJs5KPDAkS5oKohkDejplxUUVit3TgKhnm/uR+I
n+0DFsrDt6Mixl6ZJ0Ab8EiTx93EkR7JLzkmn7NgFYKbWBy/0kjtDU0NjVuax+Nw
wzatAks4DscU0vqjSlgTZzP/35b0iTh+aaoTn7cqZ6yDtyBESz6mQQl+7JdnFi+X
/ySGvKVMhygxuIWsL/0uyjUAi44WLItZXpN4bqfAIPeAVxER67X/7H/DdNUE/7wi
PGyOI/URxrW1o02T2LF+z0RKGysOt4YDlJqeGABDXwMDQpircJNaLH/8QSyUrokU
jagoAFRG+NU+Um52lVefa1QF0caxwhDTc9PUrmDRiB0lNECTs/k+XpQkaXgegSU0
Hjk1Uf5zetLY+7MlFCkQbjnnJlgBFxAy5TVkR1kSUrek5pirHO6JlnUSZmqcbeqf
gU4uf2jJ3aNNOt1hqZS4nlWzTs6f78rR5Tijb6u/nHzNh++/UcXSfRlFU/0jEGFB
cnaCHdtijmesA63r1grvHfbRm5U2H23HF1Bf0uQeaBzUKZxtMzQgcLk1A3R27bBg
f0XYxdSvnG9n5VWii9OrBeFR7zkkJJssklMaQ2NNJYkuhtkWz0xMXM7Uh9zO3sTg
rVuR0Zkov4KtkAigVZ6hA5kXl4GobI3J9Q6uOJ7ckgeIjfD2iGaHSVacU9VakXzu
CuTLU61DX3ZS3n9/085pOv9J0PTTra9hGeODtI3Vu4btnMRMuHCnhqj3b4bpZs3N
8ROy7UTwmpip9rB1jMJ+3yA6kqanoLdSTsz4lKmW3A3i1E4Wv5eR6GOzrUnV+L7r
nEuwCv/aXdO646fAXntGvevbaZ5nVprWP0Ch6gf+QQIAxsUzicmwjGHPSEm6J6iG
LzCVyPCUThgHxXH8HTfXD6yWC428KSj8zCy3HClKnfe0JUexbjMgq6fvEo5BnREk
h98eXbH9h+QailiMbdt1BGur/61oLx9F2NaZD2XBOitvkt+KyKeZ878XSO2IZeoq
nhzfwrMazyMhR0qPmQr1iHAD9aZcmnhGB4lZGQyqRwBk3kLOsSsVCei8/GLQzpeU
WZCvH4OOc1IsBdMX2H0D3jZ3rCIAjblQUr/6dNtUhvlD29PNtzB7uLAef6Q+zNCs
/Pa85B+RBTqGTyhFAnDSOturKoRC3FgcHiTQJzHAnDgwJAgaBDnZyPk7Avo2RAQK
DJ4jrEA2i16L4gVEWwPoPoJJ20MdxbRFOyNNVyQvmi+7iFUhoEu0+aw4OQktbsRx
0ak+5etL680DqCd5Y4QyjKVHtB6RyCBJ+wQP7HB5y8Tg7mOeRi/HlcPIez7oMb5L
KEA92HpgX2SzjvJornPGy1uzswATInkUM7GYGfU9XzTEqcO7lzBnR6OoB7uAwitX
taF94GQfLv7TQg8GSeuwq+bnxHX+8b/lOb/EDTzDaL2++BNVvdnAjmfvVYNyVSq/
wxJO/vR1UgMhJbvQfZj0kMId1MsdfyCo93AzJR1M8vAyYUsUK9KqvO6vmtlSmsxr
DN+ou5aHVNoG7rc3ReHO8/Bbn7QPjkhyrhlcC6Xa2oKcYmQ/dG/brSxyaw4QhL5K
l1u1ccXplzgkj8WQ2s8zO/way8ZLX/QHMx3O6nVKMPiKBaZaz65dZFieuDI/HcIT
RaT5fl6PpNIHn0LCUEag41IRrDeR2F8/JmPNafS5thAjTMCY37eKy9pOglBuyI/Q
xjBycCVzaNVrl1ky5W6yqfLwbme8XeHO7g9Ja3DOA+AtP7NRMf1TA6EmPQVn3xkd
SQraSSy5oOgB+LFS11PpI9eoftNHjp88s4OBncDKieJPC+0v0dXIXMj44rJAIw1H
3HmQWBm39DOslwTZl2YLhD2hWHhqSEx7IQmlNqtvYxq2/q9DdpXgG90Zh5H8ZDG8
rEsd5CouaPopHnFSC0gGNHp6QTvW6rTgMyd7hh4RvcuxkXFdeb6VeJtirrPPRpag
pLXTaugnvlKnfJNYe2j4C5PYc/f+/rm9vFEq5Fkanrr7aJglZF4+qmwRglgkqh9+
mKKNanM/t7+WnxNOkqoQP1ZX8T/kDxYK+dAPFL+uFgfMHwYIg+IeeeNS/CUyRobi
r8RbgJtHgGyBpmE05Ke0ddMdR077p8aMvI3vOtzXxoVUn52a33guSgyk2P1sD2XB
cHxJLfOwFlZdMLrHDe+5zgekwpzzbwom7KLPjmoJk0nt/jA+VDo/vxmeBsYpAI8A
HSKrytEvir2E7Bfmz+WT5Ye1GSVb4gLqB40QE8gyKRAn5WkIhKDWpGXazypeSeTU
bEjpK/vRRMwHLxLkpIVczWMm+TxYz/m5Rze7+gHBuLcOo7gx+NgXRODq2GHSmW9L
/dSadSMQc+Eq1L222dfv8/EY5ztrb4Ly1Igf8qtA9m/vHQinFfSlBYFbeaSnA023
zmFJD3fwdjaaTZwEm1ONncD/cvBaSpAkh4Awzg8s1RiWvt0VMMVaGwR1qiyjQSOr
ARLwtUXUtBwf6b6LkPjblrBNNEMFzhRahWpXvn3hpclq4CPMfx/3CWycbbwW6pzV
ch8FSxR12W+o1kjnaCnJ80zq0IWUA7jJZOw3ttCatstQpxG7mzumviimMewXoqhr
QFJvKaglFmnxiYm+uiMnDhFh/eX+AlktxvRkfEji+xsf7gyRWgsABQcVk1IUcPKa
tAHZ9Fn9hYJifwmYJBaklMPuJQgzPgjwjROSwvdxeYKonHwXN59rKgw/UwJIHMuW
SMr9LczhrsVWpFKxzF9fTxlCgDZ+R4ZClOkNjMcPzH5LFIccNawkML5slg1skntC
UWwoXxMTLswZE7hxvDG4r0zUhrxRqgApq5fW3h1yXiAtA9PZlgONdXdM2dHCfW+H
P1xG0Aj2/2n+5gL+aYhR0oTspPIrHk/wvuUqs4tkes4AB4IjIfT/AR8z4EO1O4P7
JHXDr5w8DZ7/6wLrWAskKUURKh6cWcKsT+8T3rmTuXTKpSY6H6/pIExbdD3zd31F
poIZJUDJRqfTxsViuSYZAemXyLnUsEVJoNoiWeIkj2sEvjAP4HxHB2/Pbx0WTgfy
7rDxjk0QrG4N7Cp/P8PATZ4jE/u8Ov3T/WKVA+GhD4MG4bOEskpmXLT45EORoVVe
A+wYvy0t1OVWpdG8yBim1OOcPMXxpVRzxsOOTkdTZ970H12dA5UAfrDtIXwg7Pj6
LoqrlXFGJf79TVhDwmJKS2ofJjPAYr7wLXM5Gn66zVsDjPDtHDYRsxI3iq2hWPrT
8PYpxIxpV/aO011yxOJNazjy+nfp0bxcYTPlrNeC8XTcIkyzNJOilZvnZX7RvfET
HkV8yGCSAro72GMDOGRQs4v9jlkSe2BH2VrbLIbBcBEGWWoRp4Q9gO80xesI+NUo
Ny2+jSpXceK6DslrL0Tj51TEsCLUJ87JgVA/VFolntlbU8rLTnyRvVa9+lFnvVjq
WQG9NsSYdLJYjuvzB0CXuwXfk+GNaJZrnk+LL2B97mEirPLBTuu4rA2yYwP9i/4V
Kat+w8NIXqepKjOZRCCwa8Lj5C8WOPvFdrVYC/e9Bgbr238jRChwCHmsJxmMrcto
rgwBkUVuDckqF8azZGG1z8odjxPnqlJIIEpXlQusDPeT1q3QzqGePnSSHdAIA5qV
q7N9+Va8bC/Y+Cgn/rbinbxkVsrOnHCKfBe/n8tJQ9AoNaqBa7oMKDdrg0HD6vyW
qYr2J+Z5nLR20j//Ouuad1x+UQ722yFwG6dLFZBuQWcefUUbLaVwENVg/1gzrXGM
7RX4l8fiL5sr37xqMAuxleQMIyxBUq2KkLtqfn8U12pO4pvnb8hxD7PCl5I867ae
ITElwhwkVhXbDFXeXp+VDA==
`protect end_protected