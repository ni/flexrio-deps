`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzkZGdUrjzQR9gfRaWjj8jjJDwjPvvZz1NhpT2yIh5+3o
Y6FdwE5Hy/gN1dYGh4DDT9pguAGrVm3eVnrD3NBPsLD8tE8s66W87DNCaIYi5LAm
ijyUiJjbmW0os65bwmoXE9Irih6fQimhx2PXNSS0t3MuB5Bxsj0YpqQRWur7X3cf
gHGKuS1g2TCDtlsNwuOyTF3dH3Lrt74KjpY1jeh66U2boof0r2g5Vu0evDtiBLzd
SsebuopSooDI9nC2//bW9MGKiYU8/A4LR5sM6SuXo7+2WXdaoG275Yav+M9RZHcS
cj2YyypL5BYVTHmgCkRO9TjXzhug3b4z3C3dDoGVur5LOZ1HCy+QVMAvOIYv+avd
cnnobUOQ8O77NWV7ir1TieNIGW/R1Qgo3SPPosgnuPC9T0IDtl60VkGjQGHDmxOQ
9mrHTrZB3chZ6a8wO2zR9kXHL4NhB9gbVEuCmLxMTnMtWclDeglls+93GSkkgrZ3
v+ZUz29J89sTWGW16YfwJPgN2tSzqk4JqTg1Rsjo+ap71GQsSD1nLgem4jeoYFIn
mqJVmRYKpBya3PZYH362DZ2igqclD/A7hDatFPf3TkixDngxDhnuqgs5Zhk7rph7
58YkMnhNq8Sho++IlSi0L28Rcjy5ma1QFBUG7OsjdL6us/A4m8jNda5RJPDnFpzg
LrfvY4anJIslVCioqyUE7wUMybXcngAU7bwTcfRfW96cAoze6MSKoVM02jKkpW0n
+Ll8Iml48hmrUXXT4//fSeeeR/LL1PQ14F++SFDhiQbgXAXg0J2JuPFAu+0LvexQ
/9PU+ut6pCTRdxSmiAJ2NW8ZeJa7/AX9PfpVDgRckspFL4NM7rnoOFoDVzxYU0WA
kSpzRlR9xFES4l4e9GqwuNj+TTNtBFborjFq4ta1yo4wOYoXAAmi19oveM30DsNp
jMkttuRtyHijQOh7zXfKpesMdm9rhYZI9de/a5+caXoK8e1cpTfKYmB1ipKYF8Rr
geg12KJZPzZjkO2UCQZgpnZ4s3buMnj9DiX0vNAQO41BLF7Fl0RqFbLXUO04pgMO
BpYCLnXvGyMtlOp1iW5akQBQ8G5vWQ62eBMG9byIt6LlwFjo9457FRpRIiJ4f6lg
gLKhxaMmqbCiP2/SSky1kVaIpnYeuX0BZy7Q8uhl+e8VEwSw9PccmdfsobA4/98m
5cRuWs5QViovYiMIkbyEyjtXJTKjzFAd9fFTBqUmP8PRl7pMxmi62KTpyzf2kvka
pF/ZZCPkgMAGXzq4P2+9GhbMdIXASm/l0ClZsJiSLRkl/doxOlHw9Vvn8Ku37eVl
4SsPNknugwLRbchtv9Du601uocJSzDh3aj0Rubu8dP+om1ykN2zIJRhud0kaslJE
LBBkGzdm+xsGX+TeqJrXM4G9z+/g7Lq+jPE5eKl2k6NqLQi6p1q0V5MoH187FQxo
Xr31tkALqOm5+2gek+NapFhfhgiibnumCGHr25abjy1ggfQe7IN6RgNJALTLUZYg
+KS16628H5xNRhcMXL69LWpD4T8LZgyNPZoEKqzA+qfU/hDt8vUMoJ9G8T+oiXgN
c7kfLOH3duj9WqnhsQ47nAVm4WgVgFUUP6Py5X7zeg9gRrkZ7Y6+7qYxERCMJNv8
Sr4ABJCHYZf3QwgHFm+CVyHNq7qenjmcg8hvubL9nXjrTmNAiXGfLHkN47TDaIuX
wi4krxxqaZGwpCbhu0pypFPGF1aWcNcX1G/wGnlsQAaUhdfzTTHMStZrE3MRW7P6
+A2TV+qIvTui7H0Fmtd3XRqVR00iRvwO6wNeIfx8VQAgGIWkAm73B8Kjbb7EvrdW
84L/VgGYBJeg4oacZ8+xoQXy812TE1l3sZoywmwMe1Tr2RmFIrRtai38TRRbo3S/
lITOHxISxMzTmpCmvMWT3r216H3sORCsgqxkvVve4qO3CCQ0YpoJFgqkGmpAjp4w
TX26HVvRNONVaSwzVluoT//Dp8PqXAfBcaub7BP0q+xEMJm9n+7hFVb7xYh450PW
FlMglpPgiy23usufjfw11Dl6gavzQLRRPlh31yvYNtZ9S6yfuHHb3Za6zh+G3jWf
urzvVUqhr1xVr9TdAWFsUcyhUolMOliLT8MqEW3HVBrnPdQ0Q6AIL1oB9iGCXU6j
jQVs3C5UZ1CBEuatJrCW9neNPZIA6TEPhqeNayB2noDNetaW4AVTZodSOSlVcj7u
5ZfXGCNfiCqBhfm67TrEpCJjPKS8CMKkYbLATyU51G4IgHPC95oW0KrIuF1XeNxK
ngPTTOQX/SVPDplGwgpdH6Z6h11wiBHNeHDmItokcQ9oUlx6VCvF2OzFpPbQK35A
TUMkTzEK53JxftktfH9PvP9XDacf/6G+rX2FeFJ2kS5Pd1bw/+s6spwf0DdFmhuX
AdrvWbdQCqDXJqmZHEoLbgHtt2wiU7/H2zW7XAlMlemiHkO5vnmvxZXthc2EkMhA
5oekNW0BWV2QaGWBpabICxmJmOaLBDhrGTCeKKf9ArRPPpil0bYyIKjrE24DZdh9
dGa4X9JFNUHe3zN1zdN0VmJkqTD9eTFXwYY3d8rSfxWcR1SNdMCFGmtaxdOlxlFy
8akzdVDo6NcXVz4sw0Jn/QNxQepTiXXjrl9vUYHm9grhmbXcHDpaZ4uAnT7uGNQT
btxHYB0gdHyaG52GuQtkShn8+dUS5GEedbFHqfSn6BhKRzJWFjJzpRn8BTm0si5j
DhoFYgbh4ayIZ0aR5MNBEi685Qy/d3zAKViV9FD/dETSd3eCS0m7FMk3WLjDfLL6
GCgB77dL7EMAc7wPNTtULnbHW8CS4TA+229iZGB7lftzpbU8rZo81P9FFOHxOk6a
VRms/H8mfdNaD60ZmXQPNOQZgqL/h43xoCham1Nhhe6FDfj1NvuO/RbMtNYCPydJ
bYgejx00z9VlxT/r32uAI8UX4KK4i6PS9Z431gni3I6kpnXsYeqgcdp4hp1lMUSA
0yw9gHPJNgpT4N9eHf0H6JNVIss+mUsOgXvi5tr6MrZXZSH89yQAgKHi1efmuLoy
DecUhij5ZeMWNk7iWI8NXWXhvi7kQSP43CvBv7oA7oDShmpDYNmRfcDQHFjWPXMO
gOluw8xdsz4sewLI9cPx4F41XBr3iwgh9A7Sd9LLLTJ/I+7vkqqBoTsyLAb8o8Ia
sxAE1464Mem4f5+fmuagnKmNvWfUEUTWJLDO2dFfAgVZB+3OElkZBSW8DaajslSL
j74cvdA0dY1UXUj9keIujWg3d/T8Xtr4kpCKogrC6MOxpdg4fgnewM5l/MZytRhu
ovTGq9tUP4GPhrtSJXXw/mGW8mda5Jg385/4eXJtqmLaDNWXmN3khsjXNMb6xgU5
IksO/XYYrzY7RRJdcGZXlCUY631j1uZUU5WZy+VGSOfCr6l8zx4nusvEiWnfsTsa
EJy+IUrv7owzPlnbK6eoA3Oh7xAQtfO4lQiAqE1qA3hR2az+DUhjwtQuRlDvB6yb
zK7Jj+3DMCTniDmSP3O1A0kxZi0q+q9lvDAV2Rn0D7GJnS3zMIbLyRRpZ0Ak/0D5
tplg0IF5mS6aKZEVwApY16kq6kN/cE3rWn6rVtATDIUdDLvXL7ZyEfiOPZO1nWLb
GUXiF78UxaslxTzdY8kP37j0Z5A+2ExxUkeV6uZ2ZGh5gi6li2BYB8UKKTDkXyGw
p19kkqpnuBlfPS7aCNuWys/9WdukoG9xD007rWylpT60RHE+7ePAUG8dtGtrHB4X
xaxp9kx2j73rVYZ6qfwj/InwX+A4sDG1FTlH/MsmJgkMnekCNe2YkE2SBIURRySs
xtnjjcK9FcxfIGKOuloD8FoPAaQ2TYCDrv3g977LQoE58hDP5CxNrBXXP1CD0Vln
St3bWrfj8/gObZIIzJ358A+cQemRP/CdkdN8NlZ8Si8C8fpEMhSCbZiJuRtYO87L
OoPgwvs3tn5FU+TYR4/w28RJVzKhC4z/rHrrC6upA3OPmVQfCd1AQYP/A/hsM2yb
iv7LwvqfL2m2W9vmn7ceSSrgirJxEc/FFDZ7Zz+ylt6C9g6yeCqprQE4eD5oS31Z
+4dKa8D91h2Ga3aYTKm+D+JsuWX926RnSV9izWguwPp2prqI6tbirrt4JKPE5VmN
b+/Tn4DgVE2+dCvXycgOg976mZ9n/ASylT59CqACXNWgX7h5P43fiBr0YMTrL0sM
Df9rVH4ejIgV1rpK+bK4IPKMtSGl2taN0dp4qGmLZuk/cIj5zEDmadNGOPXnFOwF
UOg9WY/EgLp7DMlET7aH+Cj1VINO6z0hi9tR9I0UTbZQc4142sUaPqEeYhjhbhiS
t8/+gLL2jTWgtCJiSvjHj6oKIrdLnK7NnQYr25mmtbXPRkCX0jS/X8h0KaQj+KCO
69lLYvehrlguKWGBon905QcdD38GCD3rrAXd/Q0MI+fni3BTDT31c7EpAMk+mhBH
8v7Q/vw2IflHNTUdSx3PognVFdKJTzPJAsTdLOaADVVkcmpqV5Fe6k0KIr7xsPko
nY5Rl9RO7TgiGGN+4SgFM1eqybvxhrzgowF0xd+L7RY8ZwKyrixWixdZjuG8lnVm
q1ro+ObhAL3kbq7k4LwTvC8JiCr1B46QZeG+rNE9/Y4o/IL3iHJxTCbwZwAFeqwH
vMVPAjRtHcUXDviLZ11f7z1u6igInfBOJwHHS8S9dznILb4DwkaEU9GfeY0PJ4Qj
rO+Nv35H1o308NWnw9UYjoSLoC3GnNKzjtcUk2+H80a0ekKWGXvHv0+yXd+QNsuH
JqLNyya/YedGQ5ye7MPoXSphqqP1ZmywpBGHfed5efykUwYosfamF3XRJM+A3DlW
ohIXniQrxYhGGLLKJzM1szibtNTguIsz8mYtxhFstwT5R/lEcpEsmji4kDKJp/fi
YXDRcSSX4lpQ/80ddXhdu3MlFZjnKhM0+8gF09fDGOo6Nn5gIXct40ZUikSZHe6x
47iYxmR8XPAMCYn/bEq2GRaOAhog0lPRNxETC4e8KMZWyNb9H+rvS0g34AnZ2s7s
lzw4jZCx9wylFhvYy5DQ8wJk7GuVT7+EEu0qqv2Se1GrO4Y8ZkoidX5lmzC3d3bU
ybjtb4YOWTI5a1T4Z5Z5zJb0G+qGrk52Q9k5z37iLfSOCZUGNZ+6TDdVib9/I8RP
t5DPUDXSLoGq83bG5sFYxHVA+AJ9GuEUGGAKqdat+AnVAwNHQ0wQVC3ChEMlzVyu
MTKGFORS6Qi7rRKpgfzz3Orih6dDo6XNDj18JGTi6fUVVKJwKWXEurWYDaEKnTgk
qkQUSmPyvgajOd4N335UPHFwm9SOTk/7VXkTevdWEzwjy7AINSFgpuJWDRbkPlWr
l9dlUVERVYh1rZ0uDaWGvlhsOYgkTj+MOgLDGoGD1tGgtPJ0sK4sOKFvH/+oz3uS
mLD12voJdNsCIbkbhtn+f2i1MmmQujBi04CBYuidQ9I1cs4IdjV7cPdGlTDC2z1R
GyhZfF2/RED96RROs5I0gtrblO7yWbc0xpSi44W3d1YrM4Ww++Ya318U27ROK0JX
Zxh33wC/XXghA7lfq0H6PsrSbSjNg7zSHxn/iVgT65QJVYcUbpNgI9AmWjguevrb
KDDnebrNcMEkk2aqoFcmY4f/VAg37iAYpRXTUZXTfePprlKrZLRVg/msBgjPg10n
sffB1oBYiRLh4N7nXTzxUg/vSgazN5bwkvx4XgUoBOgmi5jX2254tTwDlqIKETvj
pOs3kegWvV68wOydPdY7bFbOI3pbtumREu04FBRgEtOnwc8VFMC6plmA/gWvy5UB
HvJ01aVEwOysc1XHg7nNhq5ORiQJlddZUC5rZC6/EhAb4fFOCRJeiU2yu0b/RCYL
pm10suNpeMZeMboTRq/nPcb0zcvpVSeAFtWCieOUSkLDcZ6pWQpsgtOrOjmyPzp4
ZOWAIJOLRYrpElPWP2Cm7U5Nb7AnipDXBvxbGjDLOEFenhcS2Dgjpl6Z0gb1XFEe
YNU64CpTVco+IZd7UD30ahAHXae/JCG3zNqf1Spu5m90PtkEL98K4/zXxo46VFNm
oQDk9O6mUGiFVGeODNEnkrq+0MmDgDGDCUmT1wmU9UaEb79bGSJbil+HS15Qz7eQ
Od7k26dUjO0lBxQu40rnWwe87Qz3xlf+OmyYzrRd/Y/gyZV1jQdC/oOZbZ25+SvD
UsyMkG1r+MXShEG+oyrNu9ZTlEllqP+PZSG4cfLDbOsyerBdLaJ+4tTMpX+KYuhh
v5MDpuskt8aDhiiBIAQuFYbhoQoiJ9xeR28tL3IVZMTnX8d5MLBXHvoX5qrC/xWp
bwCiUVIPkm5qGpWhZGFa6YQvL13S+a9Nt+QIItccVop7RapufqNtAddyl0m+P/aF
tEtZAsom7bbxrZN/T+VNJYG5U2rCRrUEMCFhqrHTNkQqd6aRQP1hxi9dghtRztCH
pIbpQz6QR0rnXnwLu91GKBuYn0ivMr3C2W6qJfCwxYRaFCUI/RAbR6EDRvBYXXlX
JegplbdZ6dvpPVX73YWDhfcYkKnBrDg/Sjwzz2rkEvhQSuD84cMWBmoDw13ui6Et
a9IPreV10kw8mQ8b/YtRJa65ESalpY88c7R53EoC4tp2PJCoEI6tG/w22dXqErsQ
6hgvrTmJQkqtrXTHtrk7/7oGBjyYDCyfW7xZp3aqRJcadSQXJrseoT26fF/1q82G
RkvwisrIWRxF7m7dsIvJYcQsufxwYJrvFrSZUy88T2gJ1GGJWHyUI3oujE1gE/1B
YDl766tcK/5rmhAzbuTc8jy95v36ntr81NOtLj3LboEMhoreZKL+LB44j4hves0Q
4St2nd+9QNL4wYr3a2EK2CaNazSF9bhLofczVL9a2r0ZgZTRpp04TXNIS7P9bKwt
OxCXwN7ib0IaEx9itqTktx0W+TafsH1p0rONBBdlk/rTvrYF6fGZecznfpEbd9SU
O3u/hkzJ5y9wwKaD8HTNkmqtQv6eGy6SANuuXP6jyK7qY4/2ZvJct2/Hdop4uX3z
sMO7GaRZ6A4++8w2B4GVrAmDlALaCSNW4pWpUHq3TfhxzO5Kkx385fcSMhFBdFX4
waYIIbWhwjpbDgJFpKL1v3sBmarRAvM9wo5EoiGizYdkezZpjpnFBLCpjdgz+074
zxY8Reb3keCZaWSHXTaUT6OyaSxVuoF7/eFsBfSLqPZ+4KC8/hyinHJgKvU/gt0x
8RJPUORun+lIBFCecdLkUh3oaeioHMPItGH+EvJoA0cGJxHOHeTlxU8E4zuU29al
5lbnnizF16D9HwLzH3pHL07PieilXgWNyGZRcMN4SbnwZXKANf9UELR8kmFUKIuS
4qYYLIxzR5nA+Pzkq2/Od4mtjsdrwf62mZzNXe1vYzWUv6QoYxVvA23AoO0BXK29
T6g7YwC5Ik7VcUHwY6QI+KjBJXJONGtlDcgeXM6OEdtm7A09+pTKs3EuCIzEMAbk
Ppi3dCGFyBnsOsl1gSG/9S72bFrnbeoeEdyeHx4jzegUCuZkJTN/ecIgB9rLYeRO
TM6r2bAQrkbFU3o232qabYe7VyunSinnT8OZ1f38Adi1guawxWn0ClIFwOXZ+BBn
WdZGFk9JunWKqPlqei+WMiPbHa9HLGBHzpRC0JxyBuRS6+ZcCDNZEXsLbcTCF1bd
CRZ3PqRc7Iw1VDf+MFIwvHfNbRoc6seYSBh7DXZuituDoI9CDDRZrZTrC5v/hDMg
fwZZsWRV+NrabZG13TyuEHjIqeArPsMUWCnNU+cPQyu8PsOtku6ktz+UgBuiC+kX
HvpcbmqtVK/azq021fIMhEvT98VJZHTuiDrMEOCrwmMCt+h4dZt7PrR98C/38Leq
R4CZjUKIvacnQSZZRMeVeKpeyFiksf6qEd76YmoVZMxRf/c7cbqs7Mstm7fqMRcD
fbLTJy1881RrGMKlhUbLE57Gg5kamotE4eepn1J0v+ArX71t6oP45rP4U/Z2g4zY
aMMJldp0HxPRO+dgl3iMeUqD8D0siBXaXQRcWC5Ny176UAiQGZJ40UG0B4hxfU/+
yUDHli6Bn14jKpAmQG3FAMqmlSzmkXbwYqAJoPvJEYcTyZ9DFey2g+P05+F56eE1
UYP+jAkoomaXafRvtAVyNqJ3UnBvov5ygn4MSE7CzGV2wsMyObpdqu2AatknF9Hu
yj4yyjhngWZJu4+u4XlASihynnQad0XCA8DFUkhZczW836mngYxPcFHde98vh56P
+jz6hVRDtI4qrHtFBxYEw/karOvd+Ieev8isXZURT0vy0MYILC15aiNuW6JMcOD5
ezcW3lJ/7jrZ4CpgKLKTh4c9i6cw7XYysfnBApqDiqzBmSI5/pJF52X2xH7Hy5uV
GF9KmH0WEfi/SV+ZPn0kslckGvNSzSB2kjbySJdphG7LhcPtdw9TQI20tcLDiP5S
IIBfVgpT5xR9+2XI/2AWQbHelZCxTdLCoPKDUfGHXnS6XOsxezcFozm+umbbbgGS
ritzKtjK2K+OtO5Z5rpFQCYUsDbZOojfzyqZxshkopn1Kh6o+1SbL5omTyIajUPG
HVC1E/a8q/UYpG713XG6qvlZUQJkE+qr32iSxiiRLpUSe1sBS0PAtPCJ6ZwRcxEd
yTp02gvWwqA91ShKmIOva+Fh/tMXn1BHpOouhwakkABRoMgrXKHASHcS52U42VV/
YON0us/sJO+Ys1MTkkw2rUVkRhy//g4pClO2OLTDCnxd6SjRsUB9OgktLS8UdFiT
Scyz/fLD6zOpV46PP/GEWgpb7AUpimuIeaogD1TV6xOuyDdSqLDEwbDlrKqTw+ax
BMCriPOwuKf6qTfWTKD8Fs6bxWfQTT8+I3/UZ7TCdM6LOlPgpKVEDQT045HWmMpH
1tAuw3Wsdfw6qzm8QwHRAqmXl/EMesqAr3RpokV22sbtjWfMTDw2KqO1UuOE6E08
lyJdb3zWciRHRbdbH2P+v5XkfyjB0l/aCcLHqY6gWQgSL+/Ws9alTPepyvNWiDue
d/A6HqViCWaf4ZKtbRzumawqf6OYWYFYmfPhwOUdP2KCCwrgFiZQDe4njrOamDS9
RUU1CgoKhoW2g3WpR50Ms6GMBqel7Yk8PtD0YlONKZdESTrck1Vd4K/jiw8omEDX
7MLnyZF8190PkXvVrKdNC4AThVIu0l8Boj7l+R9Z2vPG4fCPZlSvR8xitC/X7Qpo
d5ShUtqVtWtLieDZYJJydi6fgn620KV1ykHKdVO/C6kR7kVPgHieWZSHlEEYYd7h
ORtusAaE++DNCbhD6A7npoPDofHKyfOCG2PM3r5AET8Z+lwZzbcJDbTSwPFh77js
z9ZO+74Dlb4p4zotpSQWfibcLpjO6OJpUHYAdxMRYnz6Xe20DhzYJvU8DBVzuzSS
bzC3QEIq2nzhbtLWHH9MxtoNfZiVOJGgx/hgFFnQ1PXSDRQ9hYLOWrbvu7tHI/Gt
76wYr6l83DK8oB1YX64WocLHTK9IJY0ULCi2VitTaDOv4UF4e4LxG+5Nq37twngr
rfPIleJSoCntfxO82nnXhJkFJNQOeglp84dlBERz961UDCg+PY41B8W67flTrc8T
evFwmGtZp0QAXoR916eoDXGXJKJYuxdIzPuIWHFFMyOVARGRqPUQLqDrpXW3pHps
wx/tY9A9T4cP0k/uKAKVbu6rtyEDmQQdBy+SE9UbNIcfRwlnhNaj1oANQ0bz8lC3
3fYMrEZq9eJ3sFzYwE2R/p9xGv1rYBmAxj3OF2D8pElVjSIk68SNyOniFiWOqFNe
xA3qBIq9BjMt6XstZSBRHmUVY07vRJUxiNgaSEMPk3Nn7BUegh1PA5LpmhbLZ5ug
ECQMIUAJ8Vaups/VvsZzcgwdhJi2UUF9Soyt74xE+KAea9W5Azmw3DASWKwKvbfZ
fJ2jk8DckJtueGmIbasNScw89m/evwz6ovVUAMuz79AoRZ07IFkuzFDz7nlYn2i1
VWeFQfrXdIQo2ml/u5WP8xiCVeUz7MLfZeSIDKRd8zgi6ofrUfIhVwXl0LTiMI8z
qcSB8BsIvT9j2H+T9OO4xyF/Gh17u6646ObrkEvZ1PP39dxDPIuu2JLlQwF517Ei
VN9znrVkWzVERpPJbB9RyPtMOFyuZ70llS/6FG5bNHmYb2dKU6Z2kC2tX0hmlhZn
1vQtuedBimNP1tZuy+J5YIS4SyBsMYI25U8ZW+ZfA4Ke3IBd7AhgbuvAxJLENcWa
EoTiykTYWxFMPHjCg4kxp4c4iM06eeMqUf1lpw+5PmZxQbEoAp1fTDfkiTQirj6s
Ym0CZ95Tb4KIz3Kn2M5rln9LFq9jDUfhRCG/KBc8lTvrlY1+wFN88a++e+L5QFpg
9D66Ziip1DlBfv2b6W2kiix5l/2NqXmlSnA3aZmiRXdN4UxqSC0gt1t0CVxz6F2i
fR/p0iGgC90moY1ieAED1jufF76cQO4OTb3effzlRaODpsPZchHDM2Oh3kuDAqPw
PC9MYHeC0LzX3JNhCheejN20twX8bvGNy0Y35nPKEbbEdewtT38+F7Gs5OaVnoHY
ipf8YEkYSSn6V3PSNvVFRs6ucOitRuSZ6lwyNQ+uId6GEcGQq6USWA80tQqCG6No
aATDsaAhPkCtjdmxTO2wQcryAiGym/kw3tRz1I6ep/vI0jseb0QLHGQ4ognj7g7e
iUFP/cK9rOuVr9D6VVTJ2FccH74F5cVlx1rzcjtdpsnRk8NGJHYO+cdxdXpL8/5W
lLoW8bSeEafotZ7CR0xfRIWjtJCf4ehv1gAyfSLKvVPHmV3Zyycth8TNAuIFNSLW
F/soA9/es1vpPKjiYQvvUfx4KxGNpbUEMhEtInTDRadY6wbaWp44FRB0nEF/NUef
4GQhZvlEEuZfdOaiSMGv2jd+KwBwpCCO6dI8wEvLOit5aEH6lSWBTV8bEli1yyv2
WQTSdc/l354yJRNyndrp29ysMYkYTb60My6K56zVkCEq/cwACa4uFqjAgjEXTfFi
QF8++FIFCSCYHQq4JN9qHthj8Bbqwa/8+O3ugMHoQ5nj1H1nnkaXXzfDN5Ock+Lj
VgR4lyh9fcFKOL3/SHZIiMAsl/qqJqyjZoubDOYuIvRc8vwOC6Kpq7sZSZRYg17R
1JTJ5Zta6osjXfnYQEiRBiNzBaqKAa88KaL+aUFXMyBOUJcb7Q7dzCyZZq3kO3iE
xpVYgjGr0idm3HUS7HSJcUuQyl4zbvH6+seb1y9yZroCVHvvZcXf35pWry3yckAM
K9o0Slzp/u4emrkF35tkjD+KQjWsb3A+KqW+EziXGSgtsKzyeZcBHn5MPbl0Totw
WoeIfUUO7MYf5orNPK2jT0tf6fAXDfzjD+ibXpNRTMjHuLU3uSf1NiUuKihUudt+
cF1VBh1RbCqi+GPKwhliNky4M/5nxS23Skw5VPP6TQV7s6KEXT8aSFrAbq56h4G5
zkS1u2EXwzciQ80KXO+hULMoRZy9H2o/y64ThaX13AlhE/wl8GuK6+qv8wowc1qZ
dA3txRxyu/I1GePxgn86eoRbYOKEZYF8GiL94frBQ44a9WocVTIoZKT/hSYEpbu8
DRTfbGTTjNprpz4UUutR8kYd+YfT5Q87cgQ5CJcbyxKL6UDiYjq9KoPNtnhH+6FI
d1gGK39onhPBNGbyis1Fc2f7PTFMwCxKsKuVBIVL2XB3rvtUGYQDTR6f7lyvfABX
yBp74L/0il4Vpbo5mf4DQIxoK4IsIshaSDERYEtpaWQuGObkTBnx28z+magw4CIK
yddgPSNDpQM74FvuarEkb1/K3RmVZx5NAVFwD/w1M4OHfnrzG2Jt6+qVXsKO4sJM
Vd90BRYJrcE34JgAx/UVmXyVX9xsUqvwuVbYpOhzFFF9EqflyblME1HY26A5WFOp
dD7ZsXOuXb0iVEn5cjWIjGIKPnI8B2NE3TS/XOYq8qL9yVylYPhMj98R0TIMSS/O
Ykyae/6+14aF9Al9Mxs8DauF0Z0XTC3U7VKAmRDIjUcO7pt7paUwy0BCP94dLDn0
VdZW6HGQGG4nZBsa1Vb9t60KYRui0H+BFt2Oezysm+z3BDm/aDJgD80zh6yNh57+
tJiDvidPkV70o5DC2pdBEoYCqEJBS5SnEW0FOB6PhZSrJwb65nF0dtDqS+BskmH6
LvsQjMMMIOqsEPHUc1uqkmBUfLCo5p3dj8hsFhul8lBaNfBNfTHN7WvAKA3MWg8q
LyvS41g+vSBhKxQ1HKuoiFZY/XmHGbqfFLjyoFAwWKY2ynkTqM0MAGqJ7arBPkhL
1ybi7b5ygDBHpHTmvtmy5khZYTRINK/1/xh0jOSALMeLKotonR4K98lHcdWvWxcX
HCGaOGh5sw3nX+8IRM5pQ30S7bHeTSctb7Xbc5EB3oSxRCgcEmBFYnY1yxh3zSuW
nz44hyNF+hpVt3rwq6m6+h0okSX2Vjoy1mBPxoVCbe2rWT8ulCDsU2LO1TfUTK23
xesEngFdYOOcx/GKBr+JCZUSe0+/7ZoWOI6WOAScvJ332i5PF5hnk2RWfcNuJTF7
36t80vW98fjFygwpcLR1kB3fkAocz6eO7DqYse574ji/BvtjdCLuGdYRKnlbQTew
lPQ4LCWjTSeAyl4XCds0wEzBPYcGIOTeaw0ZbfNZD8Wu/mCXFbRjh820DIyx6VRi
TTeaiJadKfzOw7nutdFi+uvws3de577N64lMj2Nmz4aqHx8EqD/qUtlyZIl0RADU
OIb4XDD3QefMyqHWQvZ8i3uiYH7cUn4ZA9qTQYJgAOsV/lEgFZ0WxVF8L9vNMRuA
v0S1XPqBDQ5QYwLwJItzbIPcMhiFbBR1EpTFQt4MusedJCaRZ/ukhiqYTosaTASZ
EONuR2t/8uYZqcqjLEP94jFbpGy2CgOTDt1y7VlOkXv3pCJ7t7lPwT37xuv+mxYr
u9nctfFrxdYToLvjjrAUsL6+kEdjrkU+HuuBgF9ipt+dGCSqhREV8FWdW17f7AL4
jv3rHtDBg07me0O07pSh9KwQXfdsWlo6fargNNddbXgN0hlXOCWdAm6BXpRdZm8T
1LFC2D3TmTY7/NXVSB7xyrvQ2vyLa5IldJiLTYk2lOFwstnud+Tl3xQIvQQsxDjB
Lg3D4CnD5wVsCHjfJXdDDs8+5Al9WE1T5Q4yUIItNxCDfaBp0uNJZoMJywTT38zx
YH0vVXv/hHhHlMBIcLi3pV4BBk546g3CMmNkAFn0KwlYkrwrUUEPP1wOZlPoeXrb
0b3qX1uNgEwEA70oLG1jYiovl87MGHgEAKfFX7arlRWjullGzUo3ZBCdGAN2LbVb
TIEIJpMJK3uKGKXnEz/AeoC82Z7IAbDwKuD0z5NSHxaFfmfTZa+EoG1OZdEPhfL4
Jg5QDAK5n/X9iFe54z8ZPqd5XnX3hQnZc2bKPs0FzEiNlE31kyoXuezw3049QHxQ
oBoxR0nKuJjb/fn2gcBasZg2gg5VMWvFpHzZpFDxzp0Yj6rsZE61jfIUszmgYNrd
usWF41IVULgWWezNPETir5LT79QioRUDF9KHEL8dHUx3rP+KfMRapcqgVVBht5Av
PfFznyfDRfXvByvbv48Yr72gPIZTSdIw4xqtIagXLs8jKyWDuPnoiLcRwn/C+dJT
Fp5ZH2yK2IA65/63v2HfLl2tC3GZPzQC0QrE9e1SUPfCNz1TV5/hFO9/AEKa5I1P
CbBN1jXxN8xfDuxEOcCLa9XP7Zn3VuGDnt4uV3qsvaZ4Oz1Eon4ggJbNo3MUuz1T
VA/lhUZySY0IRTrs/sBrIV3Hps2E0JA48AmfgOGv3PGk9WadsIWnnPp7FV8PqBtE
QJFzIfAbkI0xvWJCLIzvluWqoKEQyZQCzprYDQwhhgUwC9fWE2UTeTPXQ6xoHg+l
BIdmEnwgylYjpIraB7ldPqGVNhcCvRmEZQzQqdMOttwsgLf0N/O6mQB5vmY9Spf1
UZ+FWndsBzys6z+ybzUTj6DWpzl+Z88nSjQxAql1r2VMiT3l/tflXOlaOMAbdqZ3
hybd7vUM+zf6LmaIZmzwIMzt7Un59RZhF0fl6B68zNWMt1sC7JfgAnG4Go+E/y4D
hpRitV9aJkm7gGqXkpRbBw2T0PNOa+CXfBF1a0L2GltUuOJvn8nkpjl8oyoHcFM8
UXUNn9+UEUie/NrHXACS5BIa4OJyeyi+0/BFVbW22jzmKJkRdf9UMsFXWcj4HCEV
ILCcLpBaV4Pm7L33LDwcVGpewWAIHtIj4RnwSkj4xTMVHmiyF7lKufr0qTB8YT5T
Boqgyh46xQNdTevVIhPe4UWYrggtb3oyxvaN6iAYdU8Fwxy3ncBikIiZeAPkchGk
bCThsuPtgB9P+wIeoZBy5zbIZjJ7/GLxlt3D3CrgZd4vXyfCT7G1TFcAm6XK9+GB
q90IMQfdXEQoAxhwBeUxDaMIs8mRdCZjKiTm38p9TfXUyUSvKOF3j4p9+RqhC1F5
+oPelrhFj2ySbpti/sQT31D4eFJge4oT0AM3r32x0TAH5Uoou42/wNjS8cMr1pT9
tAlg7eVxfMuA7NGKGXxSoSfYJBSlFdo7HP/QZbL8TP160Qp3nRrhbOS8cUe9Qibi
HRz74mfp82VPlFRZdNOKvHByrjYl/weQz00JqNHZJ6WcRW29YkWXyFw4uLrzg2H4
FruKWQwy28rOqNcpDDFDNoTTXdMwjFwi2beIMSzuTcEJWHPWM1Biuem3wqf+a0vh
etwVNFt8eEQdoSspWNTu2AK4hSm3ur9XCWHFH3MgaG5A1b2Jc6zS9uURAJLn9qs/
Qpjn3hRNBhovxevOXkxnNPLXUG3eE9OPGJ4Dy7VJXOl964PIKNw3ncAAsyubeIXU
BkCmo1/XxY+VHRogXTo1J9m/lb1WnXLgnbfekxEKyVhyOS8ALnFLVFb2/MyggO14
Lexvt0rwLVGj2F3JRFT34A0KFwxE3ieCPcEw0IA2aRqvhwvp3VCPSZQ2Vpb10XT5
NHnmpiinHQI3LLElyeF8UpGz+3yD4Gtw1otQsEQdPVehS7kc5rw97e8r2W2uyW6F
8H9Mp4cT+ZPFhyC4gz3y0z9NuZ4uyKk031z5nS5GcGR+XLMrWuODBgl3rSkvsFEU
sKTjUFeyWqLQTorRXU/SSi1T8oim5Tpx3yCjleEt9H4Uo4sSFoMGntPSNyp+YraY
5aP462jOwCkfacWYhrtR6oI9j4BOafQHT799GvqJ5BWT1q5WxSvjwjT3lifPgSyP
GprIM0jDNZZ2U3r4wUxvT7fIpY1mHj9+yof5B+nBi+L7/kYbNn5uKHl5lAiysjQx
0vXbPaJTVcckpcmw64AviRgsLuIKZgMi4ZFaA+HUF8bjOS5nXaVcf2Hzl4YAoyhE
s2qzvdVTcZ7CLW96wQuHUSLADKod/QXbDQMAkBlWbcZr7cTQ0TWoE33HvpaihDFA
yXC9UvtySzwtxPX9JfdE1ZXRTZm0kcOih+WU2yfi4JRp85UECAp2jpcRr6V8DoLi
Vbhg+90FNUwasBxQ4N8ZBIEq/ssdRDqLJ11QFOPAiTFt49cmIpeij9pvCAxmJgcm
GY1yqL2nJGuJXIkV5okGFYuYSnGEx1D+Dc39sBUBGvVxW7A6/u3xYctNmPzRV49y
yNWje8nHsohq/QGvmYh/4zG983LLqfy+FeISzRI4MBfrcMyWGcmvENCso33IQflK
suB5e1VY4q0/PK8qGIrMPEStrfB16OC1GPI8BdwXNbd2bz7mUkCPg3rL0Wk8InVO
jFS1/n7oiy3Uf2TldAm3FRq6YrwksTBe52lyYRAOABy1xa7rkSc9Y+TeRvyMEpjr
KVzBE1rsYtXH6LT4de7h4qBEq5eQPYzupHG+pN6JS62ZcmHGk/8bt+t5f5lEKoUA
dDhOmE0iPbWiqvxjtrbVSZaMaEjyfh4nELRyaY1kpUF08lfZ4rTLm3Ec3mMXOr2+
TnlfLfEnd/xkiniMxp3RzzmqHJ5B1hAFfzpk/thrVUuIMRV3J77bVrmXnH4OVjQu
mJG1dZbQaeXluyFqVdhdTTI9FrKwGAvVaicxhMl3+ePfoJm69NbBO4tlyzGvrGgS
dvFoFNwvgBfZl/EqXfGxOA==
`protect end_protected