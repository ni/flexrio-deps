`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl/FaAgkiOwC2yHsDwDNDyf0r+Ya2F/3+Yw2/2nC6rDIx
XPlbBbGDs7kNhvs1Jpp7LrCidZ17O8/Gqq2v9YmumGcvgsEAHpZ8UlwA58HOgZa6
E5UA0A+WSxmFcIg+xov4b+pu4fA2IBSpQjffPmvbAf5SfvbSNWtJX2G697k6u3aF
Yf/KRg4GHtT7643PQuQTCpHTVPa8hClg7m0h0EhNvWIjhYTqKdkaLsW66WyXUvxg
KJJxtknWOczXrqCTbcbxSMZkkKefVBSn18EeX0k3MdUtIuE65Ihb6SmCCtnCwapU
V+j5UA7lB+61P1tK5J+sxi4OggpmUJxg/9q0JwrgpEuEtIEo0q4dmHO9hTM3fDIa
MtkPtOhiC7cOt+8HQ8J0K/zl5uN/yMcy0Q6noRzN0S0tolcNQjLghuPPon6F/k8u
mm4iS3tmEGqdoPkC2k1thlxYzX8/y/mPvTPFIWHMaViimD6By/itNJdX+mj1Wdh3
PP3u/GWmA0gFw2Lir0IlP0fU52tJbG/17nlOM5f4c5eq+otd8ZvTek8MwND4hZNK
ZaCZGPHTP3eHYWZ67fGpu7oSVW/8TFcrnp+5lG69tRsQraoDIKq8Ezn1385kFDjP
CxJACoEsEgIFmOlEpTTP0PHzMKr1SfUjo5aMGkD0267OBxFrJV5a6bKaR0BhamPP
+AUDbPHTcZqusSikvCxOH8n4Lurw/9wFpDTSQXCikdH0b92yqfAGp0FHZGfYIcWz
NqVPgyV5afsDgeLzm1M/siSPvqSpoE5jm0R7Ulq3Q24/bqZhWrjcM2koiM0HO57t
p2sc3FLVJEfY5tvEcZ3q/7Pi72IkeBGzqq5/EBq+9nuzKwzFnLHoJUU5Qg7a1asK
70wTzBi6RKHsu8FbsY65BoQ8tknM9t912H2N0yHbdUFtriAoA9kQ/N7LCcMI8QPS
SFLU1hcpVd6SbuxDxAYcKSHV50PaaLQv2ggkQXthPdfy0rlpJ0qu9asx6NQZ7YV2
hySr+jxUemirjkPnTUMXqb/BGra7iPYFc2hsWxmNeBfET8Rj4xWo1Zc8mTrGaDFK
p74hUc7H09FrovzT06wVDg0IenCTUsMV6bqLEYJFRbuRGqE2YyORZZKXowbvpBRk
fM7EAMEnRJeQhJE+LYesiArDR8n9cb3jkCJAUlkZobcHnfPqZrQrLYbosQH3p+1B
txpwiZu+6EtPqjhMbp2hBSoaQrliSQvSbdEVSDv3kUCyooCEs4Z/LNtbnHKI69T1
1lHEY0ggA2FBuVmngAC2mXuQUbhkeSWD1tRgA2drpKcSCQb7ivAnYmqHt0Z3MAdT
33hUffka6oVbqoHLuxMy+0ISFX1QA/tg5fGkTo2K4T0uOvb9s8Ux0+cP3xhLXI8T
/9rTAWOCjr1WVMCDwlphziHEVbjPy0aoGXE3pbk5JjZ8nlYaqVe8rhodBEfWdWW4
SLFAP85mzxoYdlYTjpSaM39r2vOD/P1WlZKtfcnOxcpHatrd63gvTi39DYxLpo63
eBGnR11IVuts0fBtPljO8r/pvUqwJnwgMBlVgm98m0mlVgKhsyv8JV78Qwfx7JxJ
FTN/FklDqjzWLIeX2D0ATAatk8SI8mkYWJsuUvULVV3kBz2P6Lv5W16rtjv5d3Sa
N5Fga4f8YE+Wq/zGkRGjQqgjh10UejrqKz8ulYcMXOX7jrHNodSzmPi/q/y8GXzk
HuwtCFFgtYq3taYdINIRDmAt3+oZGgaSO2A90kz3BjcyGP8nWqG0WnutrGP2UOmt
zflIihboKZaaKMkBw7oYZMoRbGgZWJJHGlIqDOHN6j+xy0v6F9fJns4i53hOQ+pq
aKY+mi74//VGjKEF5Bf0Yy9K2oUj9HoIQWdmS6j0IUH6ufOew/0LuEUaQHXZv93A
x824bRnZG+ZEaBEC0W/KDzM0A58Wjm+7RSbuc4Z3r7j1L/oqt09x1bIjB3AMAtOj
K7qIYRl/955ufpoe5T3IotWlN1UAE8AK6b7sr+d2A782x3FslhidTC/ZsIXYyJdU
e4Y2vDb3Len90RqIqoPtgzoTCgjE45KzViOVxFRwSQsgUURDRbaE6zQSzSZbbqEs
2M2jEjOA2PYb2q+NfZHQBDICRncTa6d438+pbYcwukyOMdClXZFnz7TsnplbXbjF
GkV9pM3WT0lLyNHIaGK6TKSvBqHQBAOl2FB2I70CxCq4V5+DTqW125JRSWroMRgi
Ar6tRFEH00ciBGmBcYkZ8l3ftXWDc18QDck4pE+nymlqldAbIJW/wIBKp/8lpbBp
u7+Y17QnnyBciuhadsokJZuMAo8L9gRyYhZXtkKLZlNHAMBqD4SihCfP/SoxH/O+
/fVgV2SP9n1Ka2VEhMW1ynODUJMhGKUTQkgbik4tUM7GaSFM+y6Hjrh6gHwEuOmX
j0EUQulnDorkdEFJhUv64hpFvL7j56n3k4vLw4hQf36KVu+E+XdXQOb0cbJx2Z32
mZ7e9lXt6u9vIRpT0goZ0ro8kOibHhwZrx8pEJbZwDtM6KmvqFV0lz8lsV1DWFEC
mQ/eOdNJVueWNKwqKB1CuxKrbb4bgFFGenzH+IKA/osuWbAyRUDFO1h0XgBA0M4U
zvQp52EySZXIhNRZUEPHhafnjNPLu7iIq7tUy4u7E9q4pFzYD0iCGfe6BwGXaADi
EbjQ4kRHRDE5sy37dO0SLhmnkAB8icblZ72aEDd4ADn1vThD/sUwTQaDqzi8ZyeA
zAKAFeYWwW6az8HUo2rgXI9/A5xzX6YlEpz/Cg7ocApY/kU9uCEOkm+K8y8Fl9zs
qTZ0b404gsFAkZQWjZfmEsfqp2M0x7r3I8SfWcS0MrzGA/4SzjYIvRjQxQZDvgHY
XdaNaeZzWUcLizHvB7KlzyrcL3v6laqqe9qrOakkfmjaO8UykYhWuZRCyowy6UpJ
urpemeJdmmpEm/yD0qb9gj5OYwmrWaagU4JBtsFAMTfWWrlZwMcrfccde2OYmQ1r
irVlLfk1QPFLYB9r7/rqcxvR7gAOBDa+gdDusFXY+14DpV81ieQ43SJuK34kM1Qw
sLrLPiE4GVrp3uEo0mDWpIyqgACfhZ9FCXVtsaWKSlZCI4ftQYZHlEXzb8kLeAnz
DQpStvzczrNMAWq8qwT/E+CLkGOgg9T6+dqkPOVr8Vw4JpUwo7O/5y8VLs1SzXlW
2OPi1PsYFaQWNJof3UKYpqEjdHsHBEdtVLiOdquHY6gFo/6/ZlMb5ZZCvrw8iRYK
3TrAu0EwJ9Wcj5vau+8rrhHz3ROr49c5Mvcrgb6LPf5SbFc1GcYpzMlqySIqKhot
NgA6JPlIXZGSqXwCVGwethd4od/iWD2BTK1nhQWEQ717BagEHJdGf2kFDPadofGS
Lm9KN+Bmuy7jel+v2Jnya5C0cLqPuew9WmKsHrJvsXlzsLoWE8Ufsn0o/cafdBHL
R3jMJLRQ1CozDIfJFj8gVJkSRMEkQgMYEIiV8xKAwpGwDAUWbjcHM4/WnX9rbfuS
l8SJQAXWmtrRK9LdY3aMnjpGjXpYgZ8n3Vip7VKX6L6p/sFCt0SpRZX9jkNO6HnH
5zrJp4G6Gw64dtb8mlu8WneEpsQiEzQPnSbzCUAasSqDtOojOB8yd8O9mnJlS7bf
bP6QnUgiYYnMKz29XoexXfhwCe1LBydF+2TsorSUcl2UgBIStpdJeo61CL7qCVCI
RAn4P85J8zwIaMdjzwRiE3tsjz+M/5jniGtpE9WqH8LGxLC5XxYGdFTfsWVel5m3
oldbdrFPiMWE2LBO0ADfKVZW8T6k0VGghpCfthXqwxxNt/DphfogBFmxzJaKOami
/hN1hJB/uLvvirRxwJfWQkA5iK9cW5H/WVB2VuDWnecXmy+gPyUuTGMs3P0wBMay
EmgFBhiIOVrEst4aPl5gFsnZj+575dAvRRHgP2KMZ7vkWzxpKhrXuQO49rymOkpf
4381A0Q1Rfs1/uH28tRgduwUBIlMMFwFKNDpNHrisaHzkEE9QzBZ7e/7Mar0csHI
9hJp8xBTSaLf7DsN1tMTArmLWZCF73kxiRK4GCQourPTWjQ/BSmOZVoKSzA0DI4X
/19ZY9CA/joEYupmmT2YqdhNg6dWZzpBSuLs0IEiUDdPrcGHGdQcaeKppVfuIgVF
cYOTedRdFBqs9BdTjt/HlPxA2YYHkqqx4rwGjxOwE7itcBUqWOXhqJoeTJdu5wdP
dCQ7jF3AHFqWyrOzX8l98gVmCPDDPujEXt8vJAH4l0rM8kIRLQlQGNiol3OxMTqi
TNOPQDbA78XA8oK66K27oQNc9v5wM2Q0O4LCFTMuaH/qkrDHqliv2Npul2T8GQhn
may7FfE6svutqofOxp8I7G6RevdSuSi34C9u40HDENeFlbfwzVpc+vgvVnIxmbYT
3oVktOD+6LuvGMXVY1MkoJ97pT7pq06d1bRb70IFtadEtgauT/dObzB3ozYUiVWm
BQbVQnSS1wRmVxAaXvH5Ai89CdvYDIEMSFVBy22L4fdn8vnQJQSJQl40OTIe3W7B
lG5BhfaPlWpGLJxt4DsVrCu0vVVjEc5CPu13gL1EO28bczdxUAUf3+dl/7hNCLSO
zWebCtQm3pc4i/5vFWeoqxRqlPmk9o+zr9AxbPT7mAo/XLNCzXjp+/opzPr5akiG
ZeKiFzoLv2ezC9uex1akDhDrUrOeM9yl13mf8nQPI7oopr3qnHAbg15ZVxK7IjI+
7Inphh+vvzVv8vBaPuiN1dGYWP7bNRlMgzbYx4Evt+Nw4wxX+thlxl9joKdZJvsC
R8B4R5noJGDVjZbt61kqvI86fnyGsDuUW5ecayJw7PVyW2DdurVAOB9aTG/KeO0g
0p+MnvYF967Fkdm8NtMYG6HPe+HxdEW18mnbNkWgVmSwI9jLxIJF5X3dksigL55q
O+XM8xPLo3/+cVvugxbsN0Gs4Lr/on/0JjigGqO/PEVMAe23mzo76bXToYK8SSrx
YAPDUqi/iKGNmcBFlcnAbdzt0R5s9Y2v9uUclw605bqMi9UgYnjeK2aXaXJ17LeI
wJUjiEpdRW1kLnuI4Zddl6+1z3L409eV/u1N0i87gU8C4QNhdyfNsCQ/f2zSTfnm
39xhI3jsJ+aV3gqgMVCC/A==
`protect end_protected