`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
EiorxhpMtoryJmXP/5pU99llRMYmPIBLU342qoA1u5feEEk/vFsjSDGg0tFL/zZH
vlGWz70sGB9EZ3sxRWjb/7ksGkfocVKxiE7S3WKNgomyWpdHBNUlv2DltLefMDC/
gN6hz4wMQur2Pzs+xQU1QYnUTp8xOGFFoIRANegqlfOO432jFJ62z5VGrJH+6K9J
iGMEZkniZzJ/zc4oAArXqCvFX76tGMSVvwAkhjdOzFf6ULNJZSOXFcnG1k7MJXv+
IOtnt7jDLMTJp7TeYPi4YUaIIR7kP/SmA43KpIdUuLaqWLZ8JaD0rQKGhyTqqMRI
V7sSoZv/mlfLdQ7WjK5z10glOMyFDxWsNiOUDNCzYmszQmI2ZXOTJZTGTIJswICL
yy9M7Ge8onnoeD/BwZNFGr6V8yfc40A+U5ROTRCbHOR30C2rK9rI4e8iRIYr5Bjo
QkfhZrkibjxJAPzilgMrc1gNU+e366qREm0amJBFkMo/EkoCa5lWz4tV3sws4eo+
kKrZLksq13eRiQYMRk60o+2K+5jsagRgLeyl9R2JAX3mkcS6vOcS31qqxA1dIjBa
HRftvEJHQ5NcVsIrT9feetym4Jf8WvPlOFEDO31U/kgQ8xm2IVwVOFGDDuYJbmwP
uO2qiAisPECg25KFzcPRYWekhcaqKXNVmo23heWEaVpsI/MaYzp+Ui2q4P3flktF
P/1jK52lIwXjTXU/LyCTtBeCphIVVBYL6U1lMdne1u4qya8s980r9ZBLZmxxRkWc
JQ+tY9SCAn3L0ztIn3b4e2mTh/bS42eCsBGnXpCW9+hpKvQPerTUoA5dfXaNak29
R+pWV15fXKpfqggqMKb3k74E/z1GvtdyIThFbJN+z0RJY/+ysmxJ64JxCgKhE5pj
cxeD/d7jyrX/26T+tGqKiE3hc04X9D7aWXuI8Gi41tVNufW9sF9Ouo1+vuQpx+eG
VLtySDO9mOfIh4hYUTJc298PiaPV4p4OpMJeJK2TqSC712RHTYrCZfMxNafS6j28
DuT/5HYzYxpZYpOtWDSPmWPhp+ZLAK3FlybESPsTSXjMv/Ex1ez9JGG7E5czWoWd
7/0stfP93mIo3G4j2Sr+TlqfKEqJBS5DEUZL7sGW0IyvZRWVE1PYeL5EG8aL2/yB
R0ROf2nKuD1fwHlsu7LwB0rctbbDxXcRQp5ZYoHGDK+asoKsBv9MT+nao1oWvovU
GXBKgfXoRPGY0WjOSG5NLNiFnDRkV3kxSdhImyZf5+9bOS5OCchi7yX+O3rJyR/t
pq1esdYoL0m87O3GqMzpe6JpqWEKsItsCNcsUXe77K8u/tV+K7Ts8Sn3VBo6kSph
x5q8AzP0wbh8U1KGj5FgOa2cia+s+cUXRRW4oXuTFwbFtnHYKtmo9vJima4g/DGp
7NgRHwvX8YGIvA9nBH20G4OvUt3QRScKMi15e1Jpmvr+QB9oFA2mqxkJcVgwzgD7
w8rXWhha60eh6Q4jYyZKPLDM3pKEQuQPS/c2oXShVoM/T5Ap85iZq3stk0dGMuLg
l321YF+cdJKE/Vsxdty6gTgX33j3g2myDG+dyu2W9Hv1Jf141ZzbEWeKW5pUt0pU
8zTPcSjoghuw8TsHBFTKQLvw5paGtJDrq2T753l3dCZhL1DCjKHpoZG4yLDne28s
1BbKoW2qkSz2ux1bONBzo+WZ+w9lO2ogS1PhMmb8npmadQYCE87225VNsZztZSLR
93lWKrN3yMyEZksxrBjMB1l37OqfohgN2wNpInp3tTURFrTQyy9wk7mBH6YUBgxR
kjS0L00HY2zm6Sd054UwZ1JfLVJHieD2X1pN4sWDQc+hjOZjmxqf9JFB/74IlxfF
dA5K06y2WV9Hj2tk32MP08wKsiSmy8kRtvJajC68XNAeG6pA0plOAiRaB55vBFwn
l7lOGmESRNJFNTzXp3tvX9F5i5qWwsRz/hfU8eDFowrGEekChZT4KhefHGeRnZ+v
9m1Z0tT6XO2WvYIDyEWUiuD+6gVnK1vWK6O8E/bxMxERypMOaoZbob5flOxbi0Um
Yo6s3ZbdUOazFVm6e9tTWFRLE6rePN9n3QmB/RuUhA5jOPhMlBU14sWCVyvcFji1
KXh1V1i51Gw8Pbc+UJl1kSMhfjBlldApy0Qo6eiLkmM=
`protect end_protected