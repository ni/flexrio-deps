`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EQKoDAcJ/8QYHXxJAKTmMHMEPyJxkMmLEubwtGhQfTplDw5fk814BAt1vyONzPiK
z3Ubytrdt1kWO7maZTq33Q23a6akYj8+fyOw3C/ebPMr6V/iTUZC9/cyITZUAT24
VLvNdbghqstu47G8Czqg7m+Qq2NiLQwbOT1ZaizNg+hUtKlecfRPMYsYi6u3SUwt
VtaRs/w1khVAHXHha9xxdn33EE5YeGPpJGuoPbcgLkr+im/NJBmMZ1P+aubppQG3
FnQkNikaMkbZkFshv9YzKhAogvtGEBdzJSxOZemGpbG8DfkUPccq0w4kHTstDaSD
5clgGgdYiBlfKbRAVVC99DDdH6Vgk18U0NcpOW6anWfr3C+z0seA91HEK5iBjQtK
+SA+4woy4H/W4Lewc0nCN3wVy8LO5eguLjsPuXwASROelIPZqMpGIb+Pxy1NpuXH
iDJp8h4fnEPR+4GrdGktO1Xm54e6ip6dqNlLC0yblSwPbCljpls5wGBN9CNnzRoR
NC821O8aV86KG9xgzNfqhNC7YXX+lfnH0nF6h1EDX+EHgpvBnRVzEY3933F0nDJ8
c8lMC5DLvemyJ/iYMd5ucNskeZIdcpL0XeUUu63UPY4WFAsoohTFWkYl7iHpkOmj
ExhJVxY5z6tykIpcJRqfjPgnaQmgOqln4otsbTpO94n22V0slbQjIxbUPFYblpa4
/l3bdg02nP7ZOa1XOvTusGSbEwzblsTzquTVMYaJCIGlHA9YtTlI9CxLItqdN5X7
wQZIqIZEyudhPfZGH6KOOxWzsF//YDIw7vH/nN/5zhmgSI/SNHnkc4CdOAiGU7ZN
buLzFtakFiUM3z9uYd5+EBmGgHsk3J9Uz+D35YgN8efky+NIF01BdGR1M8qqkR9L
4H2PJ3BPI/boAXNgUQW9/hBm+9zv2TRHOChgajqK/61bitjsmJ9LkjLI8Op9tDSv
BE3UQgP7I8Rb7Nh50lcLq2Xg4Rbg6wB9WFrlGahHSf92Dm3ERAhU0GatpXET0yBe
GHW6sw5sgTrMcEQGFtdCWoQj4l5tSfUgQxSSt4YmEtrz3z6/zM1jDr/X7FyDvHve
cZeEMBJf260TMI2lOmt48pWDSKiQsh7t++34OQZMLBTzsaEFa7t3VCJOMzIVqOaD
PQOa1Hu5+ByWLCgWq8J5Vx5hNltTdLFgWyB3ySerAFgldPWFHv6xtGjbEPGnumHd
eMBbI0SR4FQpFKJIVnmcStRFEjyyJZ1o81KeAesGxw6RnMi0qoFObhjpDfhJ5hxE
oqz48SgxjagDGTPVVP3RylGI1MHrvThS+OO8fMoDL3yJjIbxbBo30f2r8Reo4GgB
MBy16NHtt7fMoq60yGiSGhgJ/bnFGzgWEoSGOcQDGgaNZ1ZXu1jJlaUtVQdUZbi7
FEVUt7+Lp6sGcSyA6qtP/5iuOBjSCuZSmPu/S408I9bVGdNAXuOSs9xb5on0CtTq
9PrNy7gqlstqIYCc24GF7I3klYJP8SwXdhELHDangLZss6foSO5VvRQMzxtiOhD3
i2L3vZPsDF4V2CzcPK/0JVzzHXpBCt5M1Ka5WhSKtyo5klT7Ae4mfavdQBoYcYCb
G0QLuO6Qxppw2yvNezVVj1WlZSIrTzaYwQhH3LHy/bk1taKnr3ebBiqBk9SVRrYV
mw835TfM2gYUe2OCkY1sj/sLA2TS0SAktk6uiPUjbokKqov0eVhS0iceaQt6ymRO
gB5oPiT+hU7Ofrfk+FP5l1RTLxzyxRfPZOD29R5y5cne7mrtkUPCm4m47kpAr+qO
yviQUTbGrRgYg9k2Ez/Oyhm2D+x86rqB/4gugelxKK+XPGNOxP711ni11+OpEyq1
XcPhUeb0CrwI8xpyqbdE7G4udHw5C5le5J/xjxuWSa2OOfAPO9ynytwlZY0Q0IKd
tyitFrCaBR/pMk3bZ57kBzFBywpmjOYDl8CuW6ZWQjRqI+T4F/qpJIj2auheDQWb
lMbaDi9N/I+N6ZXA/2VdxVdP9PVGe6hFM7WY8ZL7W4OsoBLGRF2T/qE8wZy2g50d
DclTZ+Pmw4hSydybZWIfeYYMMGFNqg1VAAWIMv0TA7NGt/e+n8l7Y8MvxUkCKSwV
pKLxm/HMXv9T0VOizjhyPncHtl0jMlC7HN4xQ7KHPFTxwDeUJEp5isAYVmpbDY4U
kLF4gieRGsWKYKmEGUB7eEKYMwvc3CjBV8+lVl7MsSVp6E6RNyXWKS+hwGsQgUr4
0L/TYxwOqUWZSYKtw8RpZRBH+cQw3Od61FFYaoU+J9OKWzf1JQJBh0iNF5ANVVp0
ITo6QhjzLV/gdwEDw1cij/ED3QO5DMmtB+/0FVEc1UC6A79IUQSrpsWHWG/D5jqW
vgj0z2rvdhJUdih5cdgUCbFQxheTQrpbw4g55io8spLiGXqHvwV3+bg8VbasE1u/
W8aDJx/6C+lU17ni+kiluygahRXAPMNDUL0IKs36platt3SCNNB8YPlxUcOrMWMg
BAigpRW/LHsiSXhHd9AdNf7uicr9i3qS1MgLpnfdDEQ2LpPjEIksXy7fBErAb5KZ
BHyp09QTebDpJ/437ZjPWpDepZDTxh9D0n/sM/feyLkOXhKuqQv56FL7dVomS/8x
X7M4f7X/GGoqVI6QrmtJGfohH1hX0yowFFbcC7NvQd4x/zHkCNwqdh9fzsJyIbDy
6GUBgQVSuHSh4Yweo1e8UY/Ru//f9HX3kEc904MRGQsexaM0rXYMkIIF8O+Z51gL
WMPot788k7WjpPfEPJeLkSlEv+5HlVlI3uONcuvu2m7HOSgu9qVFQgW/RA6Jg0Sg
TFpcWkjD2CjJ2hmsynfHE/PNek+geHGuVrSk/8W3qyfw6XiQyvPjkcnY4hCEMIei
7ZCsSFU77th1sV578jTI8rqZtPqKsdqkZlf48O64ZrFj+MBUmBzaWfPnl7aEfrty
jOjI1ZKPjeag/K/2Ob8UDzX9mEUsb2aGuoZoDQQ/uSqdSKF95CUGA+5LwzcGKu8k
Ld0Q+GMP5zr230EzkJJxlA1kWWeLkE0DWCNc2Hd7anjCHx5v4cmDAr8H48F51vi/
zr+XZDw49OzGfTilznsPfU9ZshKfOfbveJLud2u5KtO0PubfMBVayG2Ae96Yu/Bg
5issNORgs5WWzgOraz4vE5JBCz0V099CayxOydvUBFUYWkpeI3AkwaMS02e0WE3Y
fDCTiMUxLPl9lUxx9rk9Iby+GzQDn12HjP17nUjY+eKXycUrBX3t11oxPXrREVVB
0p9wNHpCv/Gr5VzMU5lI8y9FmqCROaxdmuqW6NzPJGjkToDNq8zQvOoZ+KfIG69V
XKY9EHuIQyqtsHPTwx8wNdGgIex3B6jQ3iu1fcrHAhBvktGzjpc+hS0kN3CK3A67
ngObZudsIrhk6oAgvL33sPkV9eJ+j8L8Okd6jUUTvbYBjuZKLvFYC6C7osFkJMt9
4QVkMMhB8oaouWh2DGjQfq6dRHN1DmGAkxQZ3NElc7hUqT91y+Im/5JLRfsO8Hpw
q/HEeC1yWmr8UKbfEJ3LgJP2U8egVKQQCkfth356aG5Mer9T9I2VsIDdpQIjl9WX
8fh0azAXehv81EZU8pS9mrJgyyLtKrCmDKmcHRBxLltySzr4iniZQjZalyIUE1/7
EI/zqP26WUpzvmvN6C+z4UfZHf0XfeK0S4vVxmTS6x8QQdmUTDSj3/cqztyEhrZL
GqyWSaXyovDebXgQP3fP8rbNs/g1MxiZkmU5UHdJ01YI2qRU/2Ir9HqH+nT7buO+
bK5ivVew2Mh08efKqCvYvGXysdVaki1+FAL27mwwLK09hc9Vn6J2Jv2Le8eVG9Te
an0XqxDzuS/AacjZ5rEAGCdqZnmwS8sey9FtHID9dqSFLqTn5K+2fWh6Fw+HWGyF
3C/461h3h8VqP71rEYha8gn5WeueQvInPCDAO66REtYXH23t6PCOtgvXZ8S7ufyV
mVcF0rFGYpKEtTJkP01SJawOVUVGF96Q4SIVAhNytTBZJYsYuILIrjPXfm7I5VH5
DKx8Kf9AsR1ovfXakEH8i9IN7v6ZuTdPH+0VAlKB+1u4OCrhqstucmTS4uWNX2UC
Cok7FWw5+AKT1bm5ZxHmYVLHfcS1/0A5iArgOYjFm/sCg0y1UiuBDpC5stMIi/45
yP5lk52P423bqRvrmZw9nMgBKA2/TVHzrBTcvqKEAud9qXUk7ju7anGnUfKr3lc9
ovbZAuYofBGcRQLY00HYejvsKTiGNxtOhdPjUXNjb+eq6OuayQ/Q51VEMMqoXIkx
1rKLIa59S0gyvB2EG1xM29o48iXUwDHo7yQ6Iv5gLBlxvlV5YdVkXQXp8V/lKsy5
N1u6GBpfE/O4wtgtSBiy6Yv3mT8C13VyYvb0I4eBoOYOQnw9Blx239evXfLuUXt4
6BXbdzMKIU1eMXHR1oPyeHgUGezapuQZCrckpyXn9c0iZOO8DL0EMZsvRrgWie2I
tSHAQEyyHoiArk4GyZ3tzQBzzMphYrwylONvti+IW+2LTKmd+o2LJZkehYWhuNxF
oxgyOm63jutgm89+41akKeCKXxLOxjTw9lmNm/QSXQyv3cUbnEFNgrvNcfMk/nFO
H7/WLKJWAKwp5QyNUqbFf4qofE+/PifSrGle/v69YtCkzDkWer0XnemvV57ao5zM
NUaihycAr0JRWeRoQrgWXYP2e2wRZxBHHnxDJg/dzQl/o0zNFKSyd9uxt7qZfgxy
Cb6NvevnCb3FRtJKfpGTylzz6H6eHWczZ/hNZsMdAK1+EUNJPlnKBbwWSnnwtciA
7jHQXzyhl7Y2fItEgyLh03UDtPzLtpHMvi4x1U3ozDb18olqpOJh3fc4/W880hVr
qS2iK3pYHW/nIuAWn5eoT9/yKpJ8FR9QvrzZevofuQYNVWO08dbhNhN8cleJHYhn
LgWxLLeOhJFcSxT+53wRRGylozVRZTadgSPPKkSm2i1jNBQUwvVEHyZOXctaEPKV
Ft3J6/M1xwGql4zXuSyXVLJ4UekYoAWuK+D9F1PH0qjuxxlENEM77HFN4K23sWH6
Ixa7OPjzVo5peFMqd7laley+1zqGFMvi+PMFE5k6QoqaOhaH4P7Zt0jq+P9rgGDs
QS4xqzPJlVDUnSKnqOxW8NvxDPN1Yqo+ASj0477SsjNDkptxdlJFMAF+FvfMFMYG
+OW1kxMvIZnTZzWFDzk8Se+tcsmc9x1mM1rQeqqF5VI+YV2WKLe4G0eqBSG5Mg4g
9CQzjIbB+LymL8E/1YjiIHpGsgsAxeK72lRZOKKooXCO6ChNqKWEbvrqxu5HdTzX
PM0CYSAl82ZaFoHGuZwUmOJnStcjPbB0WWf8Wh3VJ2Gewy3MyGG8ER33qOFdd/0/
hubKzaRgcaHQUYa+yaR6T4/3IU4RMgE2sEJF7e1YxDrmVL7AkxcFdltEmWC7jS5B
4k0Up/Jfq1iOxrKo3SvzxGj4Dbnh3lrOBv7qQyM0zAlco6i35tmQ2lessD/dO0fb
nyEyWXkZ3e6HoVzsRh6JNFXEjDD/XJg5o0wOB2A7be5fcDfUzA2xW3yxcHXkHfVD
YU82fLFSBR5FiN9teaeUK3zwHe6qT37+m1xX6GruV1DOVnO594qJ+VZG9GxDdYpJ
jzlSAeeYekaTG/00+V1GbtPDqcOeMkLJMO9MRih5GzRau4AlgSMARGg80KPl5u2R
ecaw87v5hc3vbBh5aNodQGuyR3Qi7jg5j3COwHf87zpwzy88ygmwVFtSHc0++ga4
Hu7f+Y8JqXCYMZnspRoJ88pG1HKjEpIOTm6THUV8j2EPRP0u6lzfJlnX+3AwKGp+
ZSKCrLu32++OsMUAGWeDi7nfie5DeGsozVtjXFta4Jp/YJjlDux+99xprTaXmr0v
SbMmgWJVgOnJG5vvPAYdWib/E9i6BoeBTdac8ONVf9tZV8u1JYt6oDXGpj+5mm+u
rgmQq0Tum+cUwWbn1eFiq+zOKfux0Ka3z027hlQL2wr8+o6TFs7otJdCCFFeatIU
/X1DHIm2YQWJUK4HatNg0bqX/4482kgzqhGfnZlvujAr8vPDRalRBARmSPCyToeL
YlBgWD2E7ZWtoDKyj+58UDj/ry6my+l54zP5UHRAdtz0pbboKJrhJoOtUPhIjWQ6
XGTpimCrQ916yzk/9b40ZFoO0GmG0CbV0ZB70pdi+gZUM1ezJ4m37b72uY4YSiM3
lo5oVh4nRh+s8ttEVWQIJCl1r4rdl3orbbNp1WjJ4t5C2tVvT64Ga1ajh4jI4HcW
yl6WPLd57UNuwNbPeMq05RM5g9UxiSGuC4Obtg0Tcst7PUPMetStPb84dwvGwpnR
UDqrpfCl0W5tZiLmT9T0oKoEh8BMMR36di4V/vHUDlHXMYRW2U9ezkPWVs5dLLAx
ZVve/jLo0GweCYhKt50bOziSDtjzS1bu9F+8f9C3et0IAJWGoYcwKGb3MdDMQQBW
m3I1h1pK+Akz9jKT8o3a5q+a/YjR6HqOvyzvBJQw3EN2ZX94gIVwMnwSOlBqFB5f
AXGiWifDto7VWAPIsHiplq9NIXBCbIdbe0jqj10931jImbED7lwG2uFDEcV5RPNz
HGlD0kODUEQ3SMuSsLCw6KpGXHoG2Ts6q+okdtDfyFXv7nsVfiIk2WGK/7WuDvke
DeJ4Y9OUnZJndnVAAY8hoZUkPWpi7BkhHL2Xm25NthifHUlnzvbu61MHJhsnnSMe
sPRWvVa+WZeEgwwfJ3UmaskcLJUyP9G2u7+9ctW5DUGlEIFE2iZF7Vh7sNdHzPzu
ioK7zGvEn50Nh4xKqsUKARQpkvT7wgWQxh2N2H7//QILWZ9BH/SF4CzBK8E9d56J
3rgyJtRaPu+ww5KYKP7h6p6ue/r5sCr6LYWfisu87svlbtCjMSyjYncVYI5GQ+4G
5rbedJeHlRJG8zUI0q12FiyjS3nb1qpanFeLX1ZiuZ7LWarXZv5T2RfmfN46X8uk
ABfkSBAFVaK83TaOgXe8kvvAh7DjxDJzw+hZOfd94YznTBrLP5QlD112iCZgsK++
kpB9Xc0Nm6RGrdOdk4ajzQd4VmWXwkUhtwV5rIU+vwthb5wLNLK9TGR4fXF3upje
IpR+nwhhPHs3vPKSCQgWldYR0HBLuLAFyixkWT284ZLSe8nus80zzWRmrKUz4a1s
HQhB3IQLwOOu4Go/Jvgj4Zl4b57ZOddyUQccRHBuTug4SdnDdJujulKKnaTCv8Tu
PgPTxuaAPx9BERQUvgZ0dvnOJPZcEoHZi3xJ9+oT6yO3oonitGyG8/mDr8J25VG1
vQqqI0ZTQOIPYJigdUrkrRgCdlYlAOtmdj3iFAt/PIvnFODRr6FKZ0Z7htkHfyjj
UKvS0nBiWBg9hn7aV23l011eeNOijm75E+C79jljhcdm9wrpUBWGO8nWhEEp+R1I
GY9HNr/6P+DFotYO1aCMl+y0nJ/kAwAsP9aiVgDzKajuulFePCPMZL6uVqxQkiFg
G8JJ1TPVHRa22pQsDRlUfXINRsAcBQBNmie2ktDKqqWqEc7O7L71xuajRHOJx5wp
iH+6rHEBDCqycGZQK9FeHausNY8Z5Go4WWihci/WWVJphNJVP4AXYnDa8WzHNOcN
oNQBBETypcN32HaTcPKe+TvfXdNcfNwQfuPdza29wSWlNjqH9m3JqgXyRW9XQnbk
/onRqKynVhtTrsI75oOlXlxHBEMTiZj7mt+MZiHO2Kbahr2AKPslaWkg7MWqwVkL
abjcjndRYEGcbnQQfNojNp6QRL/ll+ISxy5xif9DhiT3EME3Sv4w5/1cJeVLNB2t
uq/287G6bAZZnDBkIgqI8dV3L19ltdNR3nAhVDD2cCwbuu2uweZFnciU/aXUONpU
3q7S1/5t/cA2E9fIgqDKtiPRZXNEPaccDeTmKbe43LGicMMigMPJ4Lt9VSC49CQD
V0N+cL63ijIAh0BgO/u+QNk96xWko6qIWMIb5+Dnxac6ZPU4yMXsJmCud1w9wz6b
0ewYIx5GOee+WB3nZ4crZMM7FqZx+6Dwm8NnriwLIj/O+F05wTGpL03piS1AWuN7
kprZ/kYfzomet/Z12JvD30cHYDlgK7H4yLujZmVmO50eBmfa52oh15CJs7e4Yd0l
99wIzExvRROZ5F6znTDUxTyR5YgOY+5//nUHgB2yX3qU8Ro0QKZKYlCztdvdU9Wk
gu8W6XuV4MAlWXYvj/TKgELTnvCIXY5IcQHRhbQ7ASz4fFngxEaE65dogWRZcKQI
1Yxf5ykAcWHkghR+tZWLU9SiP3GCQQ+bsGkBcQxI21olFQW2tvhO0sE/AJ7tNBQn
7D9+8W5yor2t7XXqQTd0dctVF3bovwLnSFhArfBUDNEZIx7BF1pAmDAse4ke7o6Y
UCbgGtpYprcR++RJ7gBo2TuKywT3nYgxFam1P76g6VVpXeLpq9EL33RKsHu+ddyR
pNW/b75NSmhjX0KTS/LGxbwonSYxgjvBzbs+Gv1bJd8T6upzinUaDtKGzwBMm1h0
cBXOuUXprXsApjoOocH18yymda2x/ZdE76gjc0D+DVXUCsxw/Q4NfTL+kgM6qglh
xn9PdFI0hgmucAQcW60K0m4DJnBo4wKNFuiKPRYNB6MITUTXZz0kP8K35mK77VD7
JoXhfeYq984sQlU4ti09DzFZ572ZJIlyZg+B8C8/EfHEybOc+IQcO14PvRb+n+S/
K8EbLx0ywI6lJyTS+/nd+J/Il7FGO3xFZGQ4kPwS0eoIXTdUDhpzldZHGbrOzZx1
BHgs7YHqi/Qd0VT08kOw1BROMz6Nd2Ce3XLikqR2Z/e9WbuWsyzFfHPt9puX4fgL
vGNOgItRb+vgSnefrvX9MVMtZMcwRADkgkHJkTjr79QSJBtWclWYmwD4/zhTx7wo
Yt3gicSWIFa45P+CWF8Fto4x7oF9gyNUao17qQVBUmRpQt61TMNz6Bgn5qdmNMXa
x0xNswcAyRn4tAV4/Rb6KgJ+ahTh39QCMoeKWYn6IGOA5NHeCUas5uui1ZWQyc5d
Fzfxjix+oX9DNZ/ryTyJtz53G9Xgz73+0D/wf7UHansP/a8ix2Fg2tiWjBrGQbcP
JeFM1LNVMU691WICrJ0RNl0f/QQ48U5n28HliBkpS2eoJYZDeXYONJd8MI8ZKIuR
n+q0eejnqVwZ4W0idY8SkwoTx+i3bMBAlD3r44qpQz5AJGsyGEE0w5zX/LpSW1rM
CrxLWvDnnhZIRCm7/eoXt6pH0lB3Du0AhK9/r8FQv7Q4Yrqaw1iiIvuT9xVFTMcj
8eZt0Opw9huOApHXD/aaWH9RNI30qx6XUhElsaOUDcAiOXcslEdtm6P4XRI9JjPa
p/5uWvTLPoc4AT5i2pJ/hKqxDOnA+yHhlppfj0hUlJrxeas70mj+TpC0Tb3LCWy+
ETbIJovi4VQsX9jGcA3CfpY/6aLFwqxJo81rqr8QO5uYpFVe4KAKzHUqOmNkq+L1
54210NPvN+G/RvXpOaYh4Q6V5Mq39rM7UynshSqfpTr7L9wuHHU/0a8XaReD+UdU
u+U3PJxfAZlkfLxs79STKufJc2h4RjE+dhqpZTMtdOmX8wLp+SaM84sq0fL5Gzt7
RuacNTVSMPv2i3qkHAs09yX+lFiZxvGzdQY8Mn+ABlCGEj8XnzbFNUdnipJqiEQG
s2IBMFsk1SulTCvJvemM2Red/5PjSaWwe8k0fW9JgPsfSBviMRrpSuxK9L6+dFt9
yIWn43usveINBbyYmgvabywjrAOO4oCzZCvUawlaDF9pFWYpieFmMcw1eusHdA3L
ZijqCfpR6p6YEme83z/zar1E5AvHhyRUxPVH9W+L/W/mxG9dAYlDsBKZDvTeREs7
DiqYSe8HX3Kh4DEc9h0frwYZYyM2kw/eArnRC5xwkPQHfvyGqD+0IVSfZ0GJ8GlG
aOOhPe9CJB1m28FBYWfwDrJRSe8w5Z9FxAuf4arjm5XKsJUQxKQ37f1mOjb/N0cK
XW3O4zeOl2OMAUI0qf+ygv7PnhXDJHSCDYfyNDX3ucKKC8W9t2eoLgsP0Ek1b1WF
6wIUZUQ8dV733oCVdjGvQf6+uekgMInNT+Fvtv8NgUr009uHZr0lwrY3a8Ut3cYr
yU603CMiP5WZQUp17mdOojToi1RWZmcTsfcySaWOEayAhd6CC91WZS5uI3ADNMZ4
vdwZdUhGBApkAc82MzNEJ5EIzYyzIOMZwDYzJZ+y/KmlTh+6NcjDFtOvqNYYMcvN
DZbX2Kfo9XiZFVjZBdgZxtB/LB7EE0TvgqWhdhN/nJ5AGcmnb5z6Asuog+lYUoea
4mXVR3JJju8uJlE5ZEvbMaRQJwP42Bs4ZIFVUNM1rOUZVn8PX/NugMSovqWBBWx1
mMLkgvL70B11SIvFrJbpRQIzRKddHSZY8/IK30rCczCL0k1ufriVb0eLYNHDMgBg
aHgP69lsk3qsodsHrrUMj3Qoj9sdNavzn6Z5ZOmp9fHsAMzJmcId0el92uilyKO8
YNkHzfcLlGYvhE0H8klY6ozF+180zcbeVUZSacIm+gHo811lZrCRktXNRLsCT90k
2Xb6Tzp2Af3mFg35UyYkKY/FgPStepOC2XCt/XxyxxxGbXMSy5y6awLIJvmM7N03
afUhbxhwccwC+krql/qrgh3GXUO9n8uNnXOL+j//XOfk3O7yivC1gyzKGjAs5tKO
iAZhXqR64MoJ+wzvCwHi+M8ZSPbwg9LFfCFPN+m0CaqPePTd4yyFBde3+gnajYPk
Hde/uDvO0dGJZXUENFCQf586MJV+J8gY68ZKCMDs65lBNElsIiCjubt8bAEsLIrw
3IqR0Ty6QO2mwZGUFfxxcjfjgOBN6gfzBBnCvqe8oDyrLgN0rzUKPlqohKHn65Zk
DcU1iTG5ONMC0eEaQAwn950gspCYSY6HiQM/o7VduPUTULPsjKtGsr6xaTdZ+7a1
aLcaCZLY1MaT4wLVdRB8VmMeCNBG3QER3h4Oux4NwO/OW3TDQKBNiqKzmn5dgWvb
XZXyrSlvT0mK8fBx/abt2kCv3auOHt94fV2nHiGrCzczB2zV/ml+hoX6I92s3hJf
ZDPAGgY8IFZjMbq2p2/ympt56tbNmz+oETp5rLxgdTxEal3yA7tHV2o5z9RiRYXh
Sy7o72bXNS+WyCg1MgSjSQGuxloL35ZgoK7bpgsp7jvnEtxqXH7aE79oPn0pnQ1i
ujWFnDIhPe4Aktrbjcx7UpJD9Wr3qB+PJWwJ6GPR5I+vUdCOZbL9OxmhyKNMYSrb
A3dnRG/sPyw5AViSZwFz/feVw7kN4jq42sH7H7O7PPAcyXsxQgrYQ+xOhJjeiWB8
5YFobKgKSTxAu+RP7dv5DOWG9QKeTHHrL4VCX/xLVAjHMX4w3xsFvwjHZJOz6Jo+
B4F6v0yFmbzqbkrPIf2bCo0nG3rHA/rgtFcfwsmf10iAJWbdhmdDFSxA2ZykCbQf
rBDOph1l9ex75fr6HlwbO8yQz7B+3UsGXDOdcFo02usIfgxInqhLVZ5Nil0Igxu7
HPZcA8wJW6pJ4S9gunfe6x2low06zLGEk3yovyejcaWV8ZXpoVo9dP3fetxe/b+m
ysHQHUMojpfzCvF7diMzep9Uo/uVuNz4wKj2GRYoOEecKNJebwYa+neEqdUy6aSg
fDM28UobL7cmFFjQNI17SNPqZHDqJhc0qKU1B6ELDfFD1eant2vZYSKdE0A64mYu
njnzSU8KtxOJzEWGlLSu4+7jm2OuIuSmiDQU8Bi5qw8zhLlpP5+vg7Ili1wOPBuK
T/6cNWRsCemrEdceJMgBfF6hO3c3xwhz/a4B+gvHU7PWcBtixyV56ODGmRnr3hd+
bbXCOpuS23AywuycrUKnes+KIzDBYwTPzAL4zQS0nyAOmpEZB5L1NwzpCXNMe+Zo
SfT7SvWU3uoN0fDl/wZnVQDSPRAN5AdMBq39JwLZNWI=
`protect end_protected