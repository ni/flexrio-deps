`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
wSlRvGACZeltNrdyZhP4eZKRp4i/2ept2VzAVdqVjfF64UvGUGrpjmih0ebTdC2R
VaQ3Lx5sPJqR4RTnruwoyzXp12tga9nxpp5+GzIakQZHx2Lp9RXKaylb38ZCvaUj
vnQ+LxFHC1hRiYexU/J91/1mDntvLI4+xxHM9Gon6jPad1xq6kBxq+5rfiKUBR+Z
hcUJLvTgnw5hxbyMyyJ/1JTS4tQR5fjsK/T5mzIIlPURyuTXCnvtY0t1xl4P3dRk
EK++vGuTc9ANVfAYyYT5klTtHBmN1uwyBQEWAwS32rzyrO9MijGfl0875NUmXZ22
azuk1Lj1muQv0UMZ9I4nkhtdcYcsvSHEAdB6tG+3dPI0Zioe43znUIv1HdcgS9fq
xzQaUZdnan23QGul8U79KE4NJzc1h7kniOQJxeUla2VhsKxsb4j/F8Wq89Ad6yLz
gEYdcTlClHV3gOI+4UdjF4v9oonFNKxtM9rcM1NJc/EOM56na6B55nCjBhSNYaBO
xerRoKAU9B7KBCUIElsumzURAPiMLhqlyKbWfySBUN/U3NXIXmqUY8Y1LpxYcRz1
oorkFXhnORCAty2MYR83q5nyJz7uWXdagIrR8ZTrzVG/LKJOeJ6RcrxXHZAZhDy8
IRzzUQa4WqD9AH3jfJIdEUv0Du7pqxID9xMDMflv1h9hh1QvbUIKDPn/Da+roJZp
l1z3bbMzg9vBEx7CBO1dff7VguYpKS0lDAP6P0vzLMJSYHVziZFE+xqkrkrRYdVM
Z2BnHJ2iH1tVSWrbik1TdGXNSWers8lT2JlaWD+h4ylJQ5LvkJUBE3MUMwV0WIWs
Apr5wo0Vo1mYUTvN77npYDRmLqFhfeQ/j6bGV952qJ+HBgYU0mCoV8h6jDHj3vCB
3YhNZXCRZC3yOWTFVXrTN/7oCTWrysBoCzH51Uq7e483004dLvaOTxW22RuRjWDl
sdE8UMUg1JwNCtsi4QaGN3rEyiqZaInHuSg/+5hJf5e0WrbyaeZJa5RtWL7/hLxl
B4FV4pQr/1IDEABAm1YaS3/jb6C67XDYnMc16/y7yv4hxoa+k66gJPs3+Fk/9NrI
rJunxcn1yOSl+G/isXgHSpaDXlfuvLHgJNL6tMTioZblAKrmxzsOfrX3Qt0gWWLE
ge9fcnKW7P97QG2fmaVhG8JSRThudfL8kiqJ6NV4nprzYxvRVubyp1xvVqqpm+L+
zKQrGEObUU8hAGqJBvk8hhX/TROWviJDBPiI6dOMAEeim/I+Jq3wEYEXL9JWUMmJ
GPxohQg6ZwhejmUg+olcmuTKkg64xXlViwj8MOFZOKtEhLhLK9roL0eLaBdX+lyA
8s4qstgPk7l9Q8d43rjui1iN43ldCGc2cubvM6Cd0LQnYgrpw9dgQExLiRcDI4eL
zRic9yZb23fU+tww8gNsD5BPlVhxaywyRXLPDSvrN1wDjEZn/2jESydDgSTUsow+
6fs5BdB2BNeRnRtoko63DbBZcHTPvzxHuTa7FRGWM0pEy52OrS3G3iTSqIYVZfbs
1w6zo/bfH8aZanC4IOldbi7JZjmjXEZO0CDXk+PF+UQQfHOhFhIqICHIuk1TqOjz
BHdjGgr1o7EphAjK5ZdUqeqAIy0Sdvdf+xntoOAnIddYen7mZGPaz8awxdnQpnY3
Let6I4o2bJTEPNOoqagvQIuBhmL5iS561y8+Li3eX9UiQ5jD/5IXBG+c6UqCCXvu
njPl5rp+6Y4a1UBREYBEhrVHDRyY8HDiWYYbv/7DSmG71hdv5INJsXm5TMCmhOCv
BzlxzhwzY5Ic0ruDHV4pfQ0AM+379HdTjjfLLbZwQCTwO/ScmJboU7ajf00ltyQO
Zg83lJEZeWoo7+zKAX6hSzzDJFSWkOkZzYMGYacS+U/070oU5dIcB+QM/+4c4hyb
hB3tQUZ1LgJP3HU48B5/MTDSfY6cY2YpJsAaPes4trFQoALWF/YnvZlC0ZGgPKcS
LH/zQHuGiMwDVkZIS8lxY9MmDwsRKIhcKQfpjfkAaAu8rpyZE6/UdhQRGsXcGid8
GDelihk9AF1sK4uwButDdOhWGgbHVaLe3pxrta2+Ekr/w2wEJcBKb0ii7k1khtZH
YR24HBkGhfdCfH2xXqty4R08MGh+4QwkP1Jeid4jaGFCwvq6BMWZGq7tYC1eTvD5
9L+BMKOTwqFrxWHrUYsuhVc0r/4zuGy1f95uSBUdbv58299kYEiTMdKzEgYOPkwl
5B6oWYklKsvdc7sYhGPGFxia67XcP8Cr0xY/DxoJfjPdpkos0CAJKXKVI7cyo+Vt
9BENt7ExD9hw5TRkLtW73az7WInG+67WrR0P+bhQoiQaqRcStH7VRIRzksPZLUjy
tLooURXP3rXqG3zMGy4TguqjlOaciLLmFb/t8WHRSfYKd7xcMfHxutqaF94VDEks
7jDKZeMUE61aCyY20UyriIpOsNRpQKgphGgVdocCTj+f17j4IefyOsMz6N/tkYjb
LbAw6rxAmqx6AaidmHxVrn10L2F16RYcYeHG3h9SOCRpEXevGvjqrTi+u4Wfvm3g
3XiwP9umfssNtWQN8DIgsGIibeynEPznl5/btr49IKWY9BzMCAHFylMcu/D9xdvm
P5odjt6qVwQhbYT2f/FtBTM5GQkPfX7Hp+yMD0CO5/77GJSYyWG9zk6W6I5KBC+y
hjmGMcNFceokvPViIw7HT1KEffPWgVjvQ49ROOkMabAB8QtI3InOdiNZdbUfnJ7g
00uGjVq2lDNYwTxvKaozOautVdKmznS1MHciDh01DE6agxnlGr3JqYuZ1aZ48yx3
aFq0mWBWQT+NwhYvNHkS20iq2pUI89/xMC8kQrugjhoN0G3now5+cmVHgr8JhSXy
gMCxW2t6aWvKG+NdOjfBvLdykXsIvCqxEcSgkvPvcy2gAqqPFVZOVAePqO4pi3rY
3tLvul0h7stIWwEalizm2xC9B5bg0x7T2Fx3Ua41UxFN1abWXS1q6SEI07GTdZeO
zPVknV8WNmGyHy/YOgMgDPn0Xpdz88eHzD+jYWDorOVacCu2vhNi8o77O/bJJUQU
CRrOdpcizb86YpHoXhvvG3gnn8ZJCKeS8sidilWEvLuZpdABAbuR5dXTlziW9Jl1
VOicPxFeKjWwGLecKAJYA9lPu/v6v5aOTl8WaXh8Dx3DrxVZHF7KwnVNi5wyWzku
+oOQqAakFGp0+7szlXh+akAiBISqI+s3mtD8ja8UN/YCyv55w5xYfwnDc+rTyrCQ
0HZn/wNPdWmIgu+He0jof/AmcUmm+Sg9eaBJS/rDTuxMdBWiDZootE2COSRq5h3P
QcNsgV1u18YBiOPRdBbeZ/rhxRbHgzlauqyXQVYpeDGjHiAt9zo/HdifsdCk+YxE
H+LUtyV0Cax6td5rc7a4zLlYjrnccjhh39sS6TXFGh1y+2A5lV0dlSRjVtIXaOa3
sGUcsPkpNcTdc3GYukxFOSKkqkVGMpw55JdSVh3VynOdqLBquQ1Kmdgd/4pvReCt
t5M6MebNH8mis2+BBbBlqyTxiWK0aUTGUS/0NlYKSbqg04ETOjsS2+PDcwomwvFE
KnMmp7gTv/m8nT6enN3xghYOqoexSZD2LFEY3TQqGL7geJgd7R9YKQNpEc2NrWKF
cmhOiUYcAHU1KdZ4BJ0Rde+qBqnT7LVPUGoQcJr/48/zemFtmE9mB3EOpnw+0Wry
vDWMkaILnju7T7SaGZkvInLwrtoN1GVgJWpf5Dzk2aH4M9BlVEt+1Fht1bwnXcGp
b+6RGYrkm7HZtN0Ai16yEa6fG7AB2mcTcfnWTSXiyVj0Y3dKSAvDyOAS/lo47xJr
HtTkvCf3aS71rwPkU3Dw3ieQjHiP73ohAvp+8RvIjHcnzz7gcZBj23cQZBfbTU9A
rv6Y/JtqBF3gjCQ8hoewEdsTQK+A3ET5uiPa1x4LIR21uywbLN57g3322POPAz6u
2P7GE+JfYzCkC5eVh1ABz2HjBogeYBvHMglSV96Wq/OPYcbth3KqasUrD+YxoRCi
eYROuHLcT4F3KUrA3UzdqRvTuPu1i+ogQ8LGziP3MxbsHQxJWWBl9RZymPPgioxt
xuJViA9pCINn9WAApUeug79WBTxWrjql3aABmH/hmCtArX26wVo5prBqHfDeBqkq
hdqppv33+zBlSwtPo1ig8HbQLzzodLJCHIJDOPOnk5sw6S2s3N8VsrUW5hKXK7Lp
ZEfInkFgPW7FQ2g9zVw9WWDhp+5LpVY/Be1sdwm40mWzCr8RfQNswgGkINp/+mXC
z/Bu2ANa9NGobS4/11eK/7YRYDV9mT2qa3JI8jYf6NhhpBYoTd8XboXFfcxyb3PW
wTbtdOsl2NBT0LCfaWkn3SHd4kmPdrTwJ03DK3bVqYuzqXba3/LhAWMVMD6eFIY8
Sw55gRRjH4UehW1wHLu0aWj06fQuAR82+X3/zyRsN/gf1cfLqmexLSgX3NPVOQTT
5uon9HNKC016oCskpDvrltGQnJXnTdWLzV1ivz/G9m//b+9tIj6le58jkeeeg+Yg
vo3BlmAUesbscE1olJG44NKO6T12gUjBySzL6I1j3uxM0c+XcDzkUFJVB8qu54wR
8FWbjuC6a0VBN+IbJ8o3rpTKxHgVGL7fw6U3fNVLJEMYTptEmoiNhmsu92ebkGcE
KlocduPTlS5Fj36Yhhv5e/H6SWe2RezNcfr/itKp5OVagerUvgWygZ5W6cOmfpUh
JwupClwidmKyz0Ul3yyoA3XcvWMgw5DcoSPQ1qhv20h9lxktUeRLyuzvjnjV9e3O
70f6fvinYmKtkznrjKzWXj+l+hj+a6NYcPVED2Rfsu15sig5v/pQsQF3xI895uyw
eRfUaetP42P/p7PKGYRunNOuGFayGlAXDrYFn1H9CqZu3zrMwK5umeQQt31Z2v5m
eonei6h4n7VCJol7OWia2oBN7CGZieMQ3UgTqdAQGKs8DIHfBqj15xWs3koprDJr
1T208jMVGPidCjMUDXNBQwjN1J68FT01HUSEgqpjiyh28TGsYkuYLC4Jx8t9BOKB
Sp8wi9BNZTQo8p0qm5iVG+H46/uFLcIWF5iiqee3E7oC6DGFt8nng+Cz9MLz9Mip
xIxxj2+lVdolawaPKWe8YfQwEnDG4Pt7KUVykDD55gasuorQv/03jfqv971zbl+I
ls4YzxH6ncCEtNhEZUn+ave6WY/dtKPLx1rL3QKLBzcSFSM0WCbZrR+sj174n8Bx
1DZ+oP/E2C8WhSTs89boPL9yd9Zl7a8jx0aO/JDAxmQfDvmQQ/1+nx+wDIRg5odZ
DIGWjXcQPCZ2Yk3crg6UGmtxYeir8n8eH39fRAYYyJW9IIDgu6h5APhz8RMgT7Gd
kmT6paCve4s7gsI4n/Iags6PcU2BNOR8vfh1H8mpEbz6q95FDWYgsKkul/Hgvo+6
x0y7KOmaM7Gn8YcdRxUwMRWlSdMmQcK9RGT5QSI+xBdi+0PlzMmsGSjbhKZYxIrq
30AVlY/pqDeR6PziEUy341Hhj1mevPg7U6dvfqGc+sna2S6h4uWRsQju8ZH8IrXw
WseUbVdrTQNAFPntNKqY9QHY8X73d6oOrljZvn6wkqSehsHMcSsDhyp17HEgHJy1
Cz5BmOchQr1DhFs9xJDYLfo4EIK1e0uzvy8y9Rfh/veVBXPZcZU5vnVMrnb8wEwD
gkyjZLSCourQXy1HoYRwyscWwAdtKyTBXzfp6oEgZ2ndYaWxF3euj0tDQ1rhA0RT
djfG7T3mSsfpP9Dpacof8iWoRNdqOOrZAoMhuSqNuYj/PUh7qKU1WIWvSU13miNB
QXcQrsn+ncfmJ+4kK1mSVsGLDad7t+uG2YoY57sAqMM/LEJszb2OZ8pe2pS9QlPZ
O0t1eUJKYf0z3MSoU8x4mvsJ0nPPDAjWBDfqFUC3mFjVK1lqIzfdGDL9VKkyQ7Sg
BDJJFLwxYVBM/oxCddnGnVKpmNQWIqPCXy9j/js0ezDtrIBqHiyOMSeyr2e4P+jv
JaWVxcVD1d6/LDLJz1DwCIfZRcQazqiyGpHZ2nnRpJZTDFRcaJmqUwh7r3g+DD1f
R8UExzi9JFxBnyfiO1SmzPBokkbb2KCB6zXVL9z4OZhrn8HCJjYo1ZiAhrns9B7S
GYnvAmCh4v5DlauQCsw5WFBByQgQ/GlmcYp49l0OApuZ0nuoVbbrT+ai5z3eE6Lp
xhFEwNd7qK2cVu4XHhTddG0HiIhCQPH7Py+q1jBL9W9OQe0eEov+G79sJH495WaC
Zv4r6pnnUz1Ub4CEyZfolC0BWtw8OrTRE50rfwxJlVsJ5NGGqoaKexvzfqXSsFN6
QErdOHHr7FPOUdK7c3Ybl5LQDAOKkzZl77xcnuXhgozyWUdA3LqvEokWavPJwU0K
1yVNzte1AoOIBVHlQT3iYWCP+5jo+s8ZwZhjeZaE1jCX1ZQH6AvzAUYqlYBgk9LD
6C9o+cpeZzcNUGhqLTHtyzXXmxU+gmG47DlQj0mv8C9BfhR38jWhCDVl7ssv3uGU
eBAXa2YdcYXWDZhNFQZN+FK6lWqzkEucYvZR+lp5HyhoyE4cIRKmh+TjCJGdmpLz
P5nKzobx9zIoRiGdio+OJl66+oYs7BxU6mfn5D/eTiseyryi3wui9Hr+R7vY8fkz
1reQpPRZeeKG154naUnkGWOdRFOHque5uDT+TByPX6hXw10vzL4WGEKZCYBthXi6
Xsuod2x7/v3CuTbhJO3IKvVqdduHvqhq2bU5/uEnSf9LyPLFioGks3YE3bEt+ll/
j87t0tgrZtcf042xBaX7j44V/5tjcNuutopqta6R+j7HHuoX0jYkgGeRn0eRCPnM
+QOzLITuRlZTJpyAGLHQndOnhoJlpZ85HmeLbo6hIwjqv857YrUTpt67VK44Lkjf
5CLe0IZZZSSo0CL7OpRfDCp4YsJG2svoA/IoGT/kHrSfTlueaaiihNaRoNmavH6U
cxVjyDxSPw15cLp99qMLN7RIjcd7D4g8iOd8UzI9lcDp0ytpyJRpAg2AcdAHWnXk
BJXQ3hsEWxdSS4wQR6qwgM9jI9qjYSpGXsuQG/TGZJs5Q4rpa0ItZFXNXkXezgv+
cZXJvdZwNdMFbiO/zStx7rsCa1lzoBrpzmgVTd+S5BS2O8mto7uN5VgW4GOq0qRG
lWV4qnWr15BL8duHKGKnQzMLSP5rvGoXZmPS+IMFAgKZ9BKBZugZ7ieLnf5e0pYM
t1wP8WTYJMgMSWwNDFOztSUGPyHhq3PBoMMT2O4h4pavbKdPh/7Q0Ttl5JGZqPL4
IASpC5q0cMqiJ4MM+63xrjJwc2PVAAg3R2QFL4ISLRn1fzmRHyckBwkXClQRgYTM
Xp34zW2S5mu2hE8DjRPy3+8m438AExMfLdJza+xtIubCjpeL6tGXx44ZFdK2aSla
OmNvjIRixfE4YAC/2GMGfKx03+ckfXBEdv7nb+D9SFhLdUC3V+ISIKN1wZnLz1Vc
9Ybt5dSoTa3V915bMex+RTFVxDtEt/EmXdPuKjY0/mEOydrfJx84nAUsR2Bl9hu+
mnpeeB35YIfvhjZhVcJceUvP+JwRbx+IXClaoE9r71tSSEoKAoTjm8DvyrbAcZQt
76LWHvgNBBSz5p7mgFo9feicR/HqGovUu4YUTxQjpWbSPOQvC+PMmubnpsYHhol2
pnNuZedJg3ZWPzeOE7YgLg2DIyX2DGHcJCBslCA80j+lQMSzCsVUwoZlU8PkLB1C
ycb9PkqprTqhWW7jCAeL8t05si1OIvs91aa7GcRbg2xMg3S4lJf0PAdcJejdnjLg
BUTRzSS1RGnh9t55hy0493WaenApMy9R//QNPCFh4PBFyhyfVk6ds4LgSKNr9yha
llniVOa58AxINVkxN3lFXUoeVQN8ZgAKWYrAaAiKfwSVWhd+NsQLBaBY44o8gXbj
1WNWt8mrN/iFtQkTseLyG1E35gpTsCGmJzIGLnd8DxK3kDQOtou0+77IgAa2ZLpS
wbMrMI9ja+ArSs6aMh0EbNLj0Xqa0993J2aYHRgxzUXX3iE2OrNFR+WdUVTXCF6u
GoWAYhipYLGyRWP+eOEdQeAL3LE1SFYgYnjFe8EIQf7TkppPS0jKBii/19UONbWg
GD/Y2jmfIalO66cIS+igKuGA751UZdibGZ9Mn3BfJNDtngmqQ6GzZv1k1WFhwUkW
Iuw934LmmRUphktXuccMWaVnElRvq+SutVCSvQhfllFotniOdENqFp+kmLgctZFk
ZUQ8gH61sCA+qjZKI5doIMvN+0gkgLawHObQOp4+SkChJjNK3m53sO8KRohg2AaU
eGxCUxRW2x8SvNpoNwTv8q/bcvknpCmR8T2qIp4YvCWmWekJjIRDlG2mXcqO4o+V
vKD7NxNrGSCPoPxkeZ6UQEggADQMZJsLniHoE6QzbLMHr7vEzT88FAdnAGC7cp2l
rksna+2QAyDSAlHKpJpw3OZ++8dT2/e4v+0J4YthQId2NG+cr7aS55MERb/4Y6Bk
TeLY+L4rc27i9g19Zm3PFdbeyh29HStG+ms1saIyZVbGcAJBHJp16VpCSmZSNeOb
wtaUYbBaLFwaaT6s7mUOscxlWSoqzbLGqwRCKWKBga78TxqkKe9/+6z6LzM0V7qJ
weYcEzYHQeTXNg/rH6D+cgLvtydmbq1WXTjqO6SZ0O5j/wm62SD0b2iFuGjevq6s
SnSgP049utjBGRC1vwcSEmhhGyVh9xdIz0xVAupQPTLCmuEi+UC74Qd8h/jArY7Y
fw56bZ55BvkZq1ztvf34/GslWcjnZwgH77BMPYbjC0P7Ai/H+BODnC44DzYA4RUx
dmPpjAE1qfW9mLgdZ6MW5YeC0wiob+NAycYCbZcmPcurqotHC5VrFhRClMitVcud
DQEuv8Cj+h/4tZuXhKWzctMH/tBlXBkSiN0H1GyX/MnGBq8nizsB6S8Fz2GF7Zgj
ekxNVwHbSHjX4wDWQ7t/MhyKxk+NbQzRRQfydsuDCNN0/zCdyTqR3/8z9DOIzUgQ
viLcVei52dgVrtxuXanUcFcEudKjL7UmsWTO0Wa2n8gs2Jx6anulMLJech1OLUKD
B0kPT5UJRZfh4hiYg/F5qwCLk/HyVSVOdm1FEz8WHLRqZ2of85R1Ot152FyBw2KF
wb39qw+YfR0elxkWJ7vTtfnmXhutGJoGPizlQXEgKWrdqYb0Z6eypsXfRpFNXKey
MFjP2bNv/EtuxA5/6D6MBo0H5cSCf7o31fgEZwqkAwsHalRnG+U9TwLCnChNG/7k
87TqV4axh2Btm78NhFyJwtDKmNtdHp8bVofGNO9QHlOovmTlkW5zIEQPRMhjz4+C
RPG/pHPsqunYiRU+AX1L4uv58OwA23evKSJfddMdRSpv+h+5FXd7Q7R1B4qBCqhs
nBwJ1v/y8s5ySnsbNTGX9+dOk4HmKh2TRTdoGR3a+CdK8dbtrfhgocBFmDTChhAV
9hrNUN4FwWIZyHWT+UWKB5f4r7/RlLLxuPNtogTEIavxX89d7hNSGX6Xn9INxTqa
OdGep6ynHLXIQ/80S9M9sU5J9bGdxn65+WcVGmMbvLlT3x5wLz6fUpGowrzLf7GK
5aLyNWwhstYuyg3nfdZwSH+xU+qmxrg7Bb24DbFAjO4yyvEqgtPxbcdTSdmBCixL
cpIF52mewlTpuU8HQunEhD3dv6aQlbpCDcIskiXrTdxL1G4W2C3OXaRC6kxFMf/+
RIeCDVk7PO6qSGgeoTQmyCfGopSQHlun8Lh5eCCAlwgkldnsxo50MoBUY0nB7JWD
QWj4SX2eU9fvq/JkgNuhyDW1fG9FW15jAL5+FOnvcKqS3KC3tRJ51Y/WLAlqNSrc
OY2s6Ytjv34PHLbB7J+ldpVRBHNa6pEdYgZVyFR3l+FbUxOI7NYBB/UEZyuGbbTi
pIS3Fbdz0ddm2F7musclUl/UiFkzEAkb2IXCDp2zquu7DslyDCbSM+1Uw7vy4J22
MXdEgvmwvb5hFmBaO3xNQ5h4A/nA8/UKDb0keQO48ByYuQOMYu7HOY8HTeMrD1xH
JeG7ljIxmxnfH3Zoj5TPXkdCiXNlPXr0AWWk6GeEceWC2XyPiEmMdjFfRgwGr4q7
L77xYDlqXYi2sGY2QX2mr+iRVQLW2MDDaSxkcHRcPPzhhhA1HcW/oWhgCeo+dg+G
AYe79RlyvVZLlWZ+TMdg9wGtHB3+G8/mSFt1Z2rbZhGGzp9QjBrXtNT2E/NSAit4
wpDk9zFmGft3nNGrQg3a5QHq1epeAXOiF5bMlAKd+qEUk0jPp0FAHZBEbK7XA0mQ
8siF5rrD2QTkGNaXcZWcmlyEQg+uqawBOTHoZZbkZZaPoQdOgonbJGRNFrpWg5/p
ZmPl8cZlvWKtpkgm+LUci4vPxRV9nvb1dq8WDtf23QrmvD64NyojXHROlrKbey9U
rNWdGjq3TWEU+D5NBLhdOhxA9QL5lsxYyMOc6J4z1+IdE3DvADmNorHUFy9Q9/3R
FqDCDYNUJbzC+2Y53v35TIG0AuvCaFacjXvuYFh7/HR/TwJWiXks5rdweDexVNYY
qhbHYtbCdv0fHg6OjH9SDS9cMevjBd49+HOkM1SjPPAMXkM963l4Nke5hJgmu1Ul
GZBgViNEKM2TbCi9D+0Bkia8pPkbsJHtlhul7ud4WZ8V4r5iaMateD/gApIwrgN9
zC8qPYU8c2iy3f/5wtTt33AKHHbxZMBUeG1YfOORTu5/970sC6dp7u3rqMAm++33
4ILgnOHW03Looesajw4VN4HnO3y6blpD1qwOHK3XYmlm0CVi4CeLit5pshM5GA+R
JIEynMUzrxoMxrEA/PywppL9oLlE15T9lHwVs8E921pZTXqM1XExh8bP5kJHytnj
2MISOFMKu1P8x9K+oh7c+skl4SJBT7DktjHlaTx1bRo/s8C8ImcjG0kgaT5NEkV3
TryH8xpUXg+8rr3kwGLjM6nfG/m32JNqZTZGoApJHAdTKs1sPNm4r3xR09eqUEID
fwYDcpxKkIYdU3ECZmUd1+qYhjvCkikPZm29vjolfwH2iDEm2bfWfA1Gm156YdId
ymkDDcceInfm5qivB2vpCwdugTrhoztiWt7s4WrUzluMAxNQ83SSXYI3yPWRBV5t
9CkOmYSBUTfevdtBxOqkRKSm95x7VhstF0kdPE2zeB+/wNw4s3lLigqkarLju3N7
3MuTCwQ9ZMypmWMrUVDjCsa8l84huOHUWWpwiH+WDbWlcxuYJYjh8/Msz2TupirM
lZY4NX5wdfZBwUI6df19oXbWQ8oeaC5UkW6X7Cl0mYzYz4TjwDe24IFxOgGHvVpd
gTiy/P3VbZB3AJyvC8yiD/QMoEwB3q4OYf9VUeMPRwaO5I3jW35YvgB9VwLNd43Y
RZFaHedM+3/7CB7iKLgJvn8uVj4E4/8o3c939TCOXvpo7Kq30z/iYMartJEBDzSn
F1httzNRnWEOQLsD9mjUyh2ddpBzRb7DNAwi58FtZN5n3Un91/AsKRTxbT1jq0Y4
6OZ+2pKEt/jpN3ySQ+3duu5GLD+KFwuVzSWSccP+eGm0XQhjq2HwpmGrBUXqVZQx
1tuYEiL1lOI3wLHFjvO428W3coOoKs1Z/UDSOnW6mSdBKbXD42ftmEHlVky5S418
vIhjuOsuCMV3Z1CnMQyhWiUE4HUupbTnRnisv/W9vkRmneZpLbVmY+yBU8/PXSTb
vOx8k2xTlHp2u+mdTzK5gl7iPu4+srHuVVP6ehyZr+EDms9GNAnDRgtPFw0u01qM
tQDilEuP/xFa33nC81ge6QXMHlJulSECoSRSZg3NdF56eKLmSAk2/wuQ9XKaRrKA
lhRF9GLCcPWtqSAqDIn0+y9Qq5YFWQvvzR0ntBiUemZRLY/OnjXJKk4eCpAnnjoT
ZMEyk0jazVXpcKAawNlNDyH2MxuC/8PuyWm8wtzzKXXR2AN8KWzTAyTEw1l5rUYq
6xSx/9KUovPSiGaMcB6ATZ6Er8lz5Gr1SJrsIEA0049JpuE/ih7Mck1SOvge1XKI
HARkHIRPF+4dIZWLhE8sRxiHT1EaaaMcufV3WCOxE58+6rGqnNLw76FuCByq03ii
6MUBIJK75cB4s1XPMRYNM/hMXP/AMRUmfdgFP05awp7RKTisgRu9dHYzP/itVngw
0rtxeeq74PTOk5LXWDUm/eqUWgn8c9FhhHwdKZk48HMlsY5p15O6cMSkfZKMsNQx
Jy1E6tC7Sp1DqddXtiYHtzaFz9is82HcmzSX4sl7hOnqXWatzcLGyQ2CwH2a5aoM
cnmWLuTw3mAPb9ilXf903+pIgMOScADqs3CetZPogyYmhtwjGwEncuFm0kxeIPCe
LCoaXUNDtA5olsOqyW0be3BWiAGRIfxGCVzPe9C+cy+vMenm4l5sdIMMKSWiDFcS
DiUTYoU3mskhW5wHqNV6f5T71vgTMyi9H2Mp9S3V/gGyByCF9K9Dy4EtsDkkDLi6
u+erNjBLL1QENu9T0iX7DiVk6dfMxrO+HtBQYnSiW02RukFHoinus1KA4TbjOLNl
+GSlk9E2beuJ7vDaJO2N2jGrxjcn6xsQLIi04gvmNE5AHioHVy1s2Xuw6EqO4/gr
QCe4oXvVsbv77as6bsqfgHAFi47JUdyPijGHXWW6zcu2jdqptO70K5Zpn9ukwpNh
qRPeQKtCUCjddWtehmL0VseN6A8O14RRPTdlgr7p4Px5IVZbX6HArrk8A7Vw8UBB
/DfR+XpVS7JpxfQvfZ/Srg7ckPWTKmz/GeoYxWHJtxNXgj1kjqXy5TaT+7bQHbTU
bEngb9JxvlwQMcJ+RWMsC8tfq3DtrcMyOIPE4dHegaB9NSV7ogmOPRaVPTUGnBC/
po3pnki1vWrzBOrDaazCoLZZpw2tAay41DmpkXK5WXov1b1habhLJ2h+zQL0NZE6
DG/gipeI4yWLKC8vJQy9ukFs8oCvueZQdfcv3ZQzmr6q1qzbnMyoUYibcqJAcMsW
fhigEYsuHlbx+o/dhONLu+IzX4GasBTL5OxLK10EgaHaNIhyVxjrk7EWmlWzruCo
rJ4GoY+LyBIo+P3/Laz6m2TLSaE8GLC/eANVf67VWxbTxeZvLmf6ivI94C399KKn
rVgpnGLtTlRD8p6ULS4/sOrBKH0Vvu4a8EgIhvkUwzn72yoxfDVMOJuoHIR3J0Ob
FhcPGiM+bDndQswJEjjZy6iGL8cRxH7YP4mfCVAar6AL43mKaUUshiemXsufFcl7
u4vGGWYFUhTyOZQHhk8baJpgKxRRpafavtIKWcu8LVsYTA1oI3MMRpwi4b134HhA
VKhGxx0GxVIygPVRafc6Aj+LJmkHD4KoZ4hTnKwwv4lZgEoaWKltNHCdj4pPPt14
slOIv5bf5Lifl9UF2PHDchZCVQt46lkE3OjOWrvFHelpjUWldk2ZTtJ4rfB30MHP
yD8kKD7CmyYhiOS/nztJG8MZgOEyN6QiYb6D8b85120A/BJMKCM5/KjD9v7ekYkh
kkK5hBN3wZb6ZumQ6ihsqyCxpq17g7MIakxunjnqezQ2u8M2RJcADHnY3rC60cfN
CAKMSvBdXxB4CWIpaCmzaqhmt/TfIaA5mc+/3hstxl2oofGf0SvGeq8ju4iMkdgr
cOgm6pWwvBXFZ0YFCOO6AoNTavMh68FBtWXGRpsWwnPp3DuaaNuLnmYY3uTXLLOV
3D+pgRLveqoBMUQoEC3pdQ+iU/A4RCeWQz5IMxLY5cV/QXgNlKTjBMcEiha/Vcur
85szcX88v/PL+aB9qBDjvmvB+fXY7lQn09lW60JvadIwanylx6PGkgFTgJWAxO/t
lwwSgTVS4Nf0Gqgeccndr9189ibh9n8VbLhoD+USTu3hytXvVkogC+eX9tEEEsst
KuVl/J/Qg3adHSJTOKkSZC6f3elQFmmhFkObaPxhu9IvycK4qhptWuSzcwKIKpBJ
LWpym+FiXqUgLOaRGcQVlqbVhw+rrQZ7bRw/AVI3GqdXgbPBGtXVHEc2QW0jt9hc
ELsXrpIA563riD0MYNtobmicTiN0Cdg3gqvyIBwoZPKxeXwFrmRfANEkteIVOYVR
vrB17QMrmPGPehyPWJBOmCBlE0tzr8DLC73KmJkPW3Ad8BFtMfTjJhNHnHcc2YdI
5IhzthJX4uZS9b6MV0GTz3ShacMzvF0DxXqLI2r92b1bl9oAX3+ah4mt6DDbx01m
XfTRX1mihq1H+Hbfn2gb6NI3pISZbZqQmtNO4vjPKPiEcLnkrWclHLBUXHVVfLMy
+VI11syppDxYT4syr3t2mpI5sBwSD1MymyKygjoo+nFmmKUsCUYr6ud6kMdgJ7jM
xL4xAJOr8qFHvMmyZ1R3tO8gtTTXGoIgocXmLU1dG42hUwfP5Pc1xeUocbTj3aYd
TMxr3QQogKQB+mMapeDh8hMQfvEgMfoFUOjsKozBoU12eTeA3iH1Bf8dUr2uJb8D
7FnUxl1dCF5eboNmmMfdTv82cDZfB0UFfQnKhV69cMribQGzStpFDwv6P6qYPklO
aOTyt7RuqwUtfWEAxVW70/uWqFTE/U2IXlq2lBUr4XSQ7aIk7XbwlsjEuf1JbPTv
5hfknm44MLXhjMj//IfIuVki0AsumwD4bf6JAWzxsOLB5POBxosnbzEnNUoxY0Pk
3GD8UU+K23QGHw8Z4FrF4j7jvdXwvE+rpX2KE4WkXD992c5G4vAqtHyVPbL+DVx5
fsk2OgIB6Bd2DBT4NQulrIFJnKSJsSkgw6xCsizWA58QvIumb544p6h5XvUTnWa6
LM/tTjhOlYK9i3no9tsEH/gL7QoDeoWbFiXT9JVz8380ylH9EeP8siZfSb6koECF
QkzcPZXUMFKZvzB5012hyJQbr4pasXLgb+N+TfvslYaFtsGqMYKbkNONkzq+7Sri
8Vw/Xaqajl0SuCautAweoprzMNgypl4DWbPHTVTFxo75pKpbvu/LOgZ807Yu4ut/
a8MBEGBlwKXkwW5AQVobpFkoVLtdXIZCJCvyOw965ulk5DcZEsnBtgMJVJQGhFbg
gSJIjWNRI7fp7brwJKAepQybPi7+HRplHv97v0HQ3Z0Ta+RgKGEH0k20TDurwPJy
yupsWd8N911IVwALYaCoACBJX4dLR10y++0SCpK8jQos8JGdSxDoLvYurkGFB4V/
2/VpykwL922DAlWG3c1oO4Mzxmqsp13ePlzqbXWekvuBOUGLrggP5ujz7fGlc+Is
f0PNx9hqpNBnNYNqExz+7uO9O+wbXoH3hhtByH4SBDIMVF/II+pBzPiJROUmfKbM
7ICLimpAshI/IH1QupPWXA/wOz9URJz6AKVvtyVu5Rces/GQrpaYndzrntYVKSHC
tsOpC1fEMQPeeFWbpS+i1k+SIwRnRT+xd9+wDPjkioxfYutHHtKvieJdLZHZUpVo
+cm+H26PDU6P74aEB67479LB5cjYPEoDnMvq+tmDuiF5vqgBuqKJcqi2F7sQ/g4T
TsNXg/en7woHsplJMTFABUs1oux2wR6trRjfpwg3cKvjK9Q2u5+QkZulEpkDzEGg
kK06/dkCotCOFxpgQMrlZ8yoU0P+T6fo7S5wB7aLhu8tXNWoSq4tJjbxEZCGdd4o
uyFrUcTLTPCBY7XinULfnyULEs8HTR1GW+qAhRqPKukxPMeSpsJQmE53eOuJS700
8fYcLhd7wPuEoXYGvNRxd/VhXB5dzs6hHoEECXpu75c3QAI7fNaAtNu9B6N4IJNk
FCSBRVomc4JtHb73eVp62PVMCuw4uymwhP2nI303S+W3nXbS+zcpMmD8Jspk5Qqy
5y81PlxZY4VwTtKGBp4X8KpsS8P/mERS/2WpmAvUCcb8OdQcCWDyuyPWeVESa13P
e3r7okxhGelt/bRLor85Nerho/eyDq5ePY9efUe9eO/xSPZA8kC0C3X4wwoIWUHD
XEXQmq2opIzwwAaPPCGKBTVr7vhpUMn6JAJbztKuvQGuVPOrNw432bHkSk1qygUU
MCmqTuNhs1gyP9tdJwjxwnOjDmxItVw2lQnyHLi4X/RKw2ApvnwH3ozTXyDUyPV4
9m53jcmc4JDX2k/TyU0J1qFpIL2Nauu4rJDaI1hy5W1v0LaQdcH1wOYqWEK1p/ZK
nAr7YrU3sStBF4O+8mlwujXTPGPps1KtPsrmN/NdvUfxt/AFrPbgNnF4fIV6bqDc
5c6ShNdGWqqr8S8LrP/Ko9EN5o9vGngBXO2pdDuAAsEf8HnufwtKQ12OhvnfvxwH
j8TecCapZkPKzKDbXbiUpVGj/PSt/TtWgsWkhH+Bctmlv82SH7Ud1pCMGuZIC5aI
DpFMb7TbX0mDaL5s/0p+XSdqewTlPV0ZrGL3iBnsmsr4DcQdjIXgntBy3qUgECJe
uCJkiyGFtn+V/uc1WclDLPWEejkcPKW56VEtMnTmsSoSiv4kZTGP0p7XqeRvsujd
9bGbZedb2dD4bDj9cWdYSHzg9tE0KMAcGIvoC9CNqs6jv6ghtcH/F9waBBEbziIE
0KGcZyKgg1fKR2MRzznKlBMrSs+NgHyz3h7l1HVVwTCLJafF8zQRCAx9jXHGF4kM
UJuGlYmuuku35KWct0Z/NAD1XBu33r1SB3w/9qoY99joQy0DHHkLqOCnTZYDebXE
d84ZzSd8rceeDGpeOP1l9qPBsaWGAMpfE2pUrIq70rzcY+wq7LQVSpMcR+xvQSqg
lckiaAcFkdyaFSkvHjrWI9gg7v8jVYbmPkawdWjtUBzI0xHAGuechZJeBMl9BfKO
2ndkHLfurTVp0ehlWIsNB9QBeaB1QIynv52RtgN2rN/xZFwkQ/cRr27fujp1UZsJ
uzh2rbAyKiI3gjICB/yr290zdatGaaYjoTWjjspjgyWPz2Gm/WSx/pD3Reo+3hZv
8+a8lSNgDdbw2ZDkNS/wGF8F0juSQZDR6tMCtpgKyLGYpQOGpdajM991qRyEvGGI
PRgDUhC0RgVSxnORT4qz7yBC/ggeFiLtAkUD5PA0JkMRw424P0Qom9VH1DC62dp/
fMqZIlaieDMgd+UfHSQpcWTxrGKTnTd5Z2d00xBV3vYTSrpziX9NP7Z1NxWlRMx5
fQMzzSErFtBOMg0Ri9axe44tIjHcen67RrkgXgBuyoOSnsuxI7kUhxfPQxZsD7Om
DZf4qGWulY47ZtcYLL+B+KKXnbT0/Xxb2fHudXII9odjVi8bmImr0iYxD6dQTowf
94ID9As+6Q67/J47+Wwe263UWwbBxREdT7Ed/wzyRGVvB4n9SEQFQi4Ptxu32o3X
2A7z10HmFnCSpLq67+gaA0Z4HifsHiiR0XB/wVTbLv75KYSUQR/nRj7385Ox/nQ/
lyo0ak2i3x5MCvxJ+1aEjBJWx2aZqAgeBcjJQmBYQMJbcmbD7etb+159TZyS++T4
EMSLoWyRdAhcQ7RlhDcbD7MCFS6JeNxIMmOV9hA4z0uKBB0G/06DzzytyiCQ6Q4p
8988wGyhNMkmamliNlLl2nnIT1CUYwU6x2dfspsIoEXQ7Xj3WqRoyL5e7Qf9GGvU
NZiCHEDPqbeAfsQcCyaAY52Hv+exuPS/njbp0fprkie3Rw189/cMVWN1seySo3AU
zKFFhN5wJZtpGlgMbrqszevwcaCGyPAA0U182DHuuYRfSarxOjGRfILP6Uyxq3ZK
OtnBU9nt5E8r8jFQkygzvm44HzlyMOG2/PJRUsut9SLXRC/1CHcYcUq6OGZ9WU7a
Yrz/3W2jqeGqk13DZCfE2Hxrp7FXVney+bJN6K3Uv9rvprcrtqVslFJHm2ar+RZh
glDO81Y28QbqZs3aaMde4BeGBfON5rI+Ul25wQaXU9BGNDKgXX7UQU11Q9kRPi97
w8c0DbJ1R8gO0GDDIMEerg1fulZUFYplHXP8RULS93H9Ts5uDQDiInIzubJUztud
hkdc6nsDeJIV+lUZrkZF+9m1ckQj/R+Ss7ed2phjH1L7Mq+LsBNl0uAwYDeBZIct
hY2/C1vuM8XlmUHx0xMIBU708bC9SrnYUTWLK1yES7maSB+XC6nR3c8x98jTivod
YDWcSNjTpVy6UrWwEqtluuyzQBj9F5qk+hL7P0SwhgNTUaX81vW5FsWA+VbLzVEl
K3sbhnD6toASnnJ+gugdDkCONKYpHFRJ0O/lYL3qsHKBi1Fq+H/0xaxVwt3zQG0D
Vfz0xnfsIUrUF+0yOpCJnrMopvzpU/29ZOSJWJVDcIf/gJ07v7PykvrKViFbIsNo
AVS3wOPGfkRvHSR4dqLH3rkgez22lTRg5fbWRAVb634laYlCpQszscl16miooxCa
VqOEpVcSA23NBZjGPNLAAsOdCxg6Ew7ZoZjkPQvi6upiPcMcZZxAV+9cNvU4lA/i
KuDJ96FPHYxhyurVY2nTo1KeRBWpYkFvjBFCW9fZmVgJu+3NYkEZoVcbnI72dwM9
TX89VUE5/U5sQSW2OZ6olpa7pRnLtdPwHlO6cc7IArSr4Iox/lcntlCU+9t6ktW6
u2LJouCC3Rq8NHTVQlQrkpHQp60JVnj1POtnwuzcGV34QOJPUnPk5kpJG4iZymkF
xQVPzDOA94TFFHNbU6VP1SD/xXL+WOsK+j5vR1V0ACAGOxWYEk05FP0YWrdKUBgH
R+VMcryED3WfpT08pN20892Jr/PWxKjaAAoZ42sijYWKQ56h94daezly5tNAIvXa
VzZN1FE7IMC8HBduJJCb95L/mk7wXVSLRzks9jJ+yjJ47LEf4Wvkxoa0Qljt6H45
sEFaN7/IGPqMYVc2BGEhtgNzg8pk5FyJVCSA6JkbsEFDyCVQE/1kYoWwfDTjNM+h
q2RYXJvj5/uwmE1I3Wfomq91/Lmc2i9GDBOX/8Rw9dMlRegSa2QnxVLiAEH7heh/
HzLlyLljPNKw6En+gbJV87LSHIkO2vC9kspqI0bZEgBFdr7YUSRLC3ozUifdx7ea
ZwQUygBaDZtW7o/6kGoozvQHAVjPauO5nSLmUJg/ggpX3N6GXYnvoqpEVAIyeT7M
Y1kdgC+FPR1AwKsE3m0BRNuzxC88iLghZwFXppZgEHHvYdkm2VUXwe0Pj8n++fZT
tQ2FYGtahaQmyRljE2lGUO+rHPZhAsViKjwXF3HIKKgCEQHJWoSsvGCcXdM8DbHA
WgxTunmCR1PIVEiAmuCJ7vZExlDQEEEAgvRtd/VhJHUPHvwk9M5/4bNWAxUcPuyI
lLaEgB1qKZWtUnGmqvWV6P9X8N7jSRu8NNcVaYX2wgU1o9nIoKxRc8Ou2ErrXjei
QTIGFnEYQZNiwP9JFvFf0QH3tODT3rCIkDW9taTBn2l2TrYaT1yN1eZ43pnWMIdQ
0HYrbZNATH1zzVTuJ1EfETbfwIUsPKvX64soBbep3oKW5MsK8qGY7KpZZ2CqiIt7
AHYxvhvSezK05TLNbao9CA4TX2LIvlr1LQJ2r6J+DTa69qYjsYvnE1HfgR7OMdM3
9LdFXgoUEGmzm/5eI/dtBacbAhyJkLe0F1EJv0te9xHjeDHvBwg5pjViFUgjQjJz
lqAOtk0EBkmmHeMWeQYnqoJQn09pHZ5ngQChSrO7L+J3DsWghr9nlHZHkCdZoeGi
C/oEVmnGlFoZwofkJVVRbQmH9IhwoQnRkAGIx9hXPhvL/iO1BtwBCXljFIPt2Ntd
uA62BvuBh6c7yUAAiE6PZjGSXarZ26AZVePjhRRcWu1ddVV3QkpIkFKj/6bQFYJp
dCXzzQ6TsfQdVE0M8+Q/Krc/Q/1AT42p+H1g4NYNNc0e87fkFrBk8hFu/u3HhztQ
JNJ1tIOfKrXtDWLIUyaazhzw9NBQ7esRmRhzRvDy08ERq9qBfNXWsV33+92AFEHt
6Dal8FG6C7yi+aE/7OzYr95fGb7z27ydb4UL3nDglGCTlzDwPa0BJQ3+zVZ5qeI4
r1TxNvwsm5HAUNgegjWz1D96wKO+1bVz2Vh74J+gyXmQJO5KrOv6Cc99PWjcYydx
4u8lNlc+8fOOyq1e5xhfAix34wVhHYH8POtLs1A8l7KdkfvNUbQ3MqkCCSmHRbS5
8qpv3de4b6EvBxKGDdifARDzGhqPT/NkNbdWhs5rYJ3csEzNy8SnoFGGCogkkqtt
vTv2GCEl1AFz65AyU4N1TtkDyBn51R88afmbT6rhYCCm8aPdRcVKsu0YZIYIE6gU
JqcJQvOgRLiIP8ydD9d5vgOE7jzf8INktcpOr9HbtkVTPo91T1C7pVMqnKSMaC3r
x5T+CaNmeCKnxj2S+/QXk6X++PU6EGbBxu8ZSEDZlBJuktJRdjsJ2HRXrwHNx2JF
xNP9cks3Sx4vlLn+16BBNobQkBo7+ANN2X/yHYgOCn3UQLG5yGIg3NvK69wZiiAz
OF7gVZFkx+MAgwQG8qIjYD2XfIOsvN8biGsFD3VEutniD2/ylGgbxOJdG97KyhmU
vZLpygvmsrqiVX7KAn/4FcpZ+tnhfgCkbhqtq/uznIKU4IY7gXNnz9sOuUG4ovLg
8mMf/gWy5Bp6sKdoU31pTCJOQRk9NU2JDkSKSA641iC6KBQcTtRN7cpjSz/Fz/J1
2IrlVNwfQ0K2/gS0jxgcQSgHPDDr5J8BoOPWlCPlBCU8wLs+j+d+Lh7VpXe5Cg9L
h0U/PMbGJgayR0y2StTyNJjVsn71JiTt8YyPSjM4mdbqJ4xnaQAFgQ99WLMh6mhd
Y2pO/xLG6wgg8t2JPyDUhNXgAqqG377HRi1AqaXA0nl8edhnnqlhqjQfaaAA3kCA
k6dhE5xJjnOSZCODTdxmZnUylFMuBiQqp7iivLL5lb2r6r7z+SfMwIklxKK2abQt
yTfImi/MEdjqmpQCnhE657gPDZDj589COlAx4oHq8BLdcY7I4DSt0XtA4bXB8RAY
kgQB3WYY/8qsOC8Uyce6ytPIv7ltJ9leR9Bes2cfGETRA0XpaRkESBRwDI8IIe/s
zdATXEtIcmhhkAfIrUwGDrRZTcrRfTqyj8vhuGUzqO5/CWeQmmYAprh/FaMJUhTU
ySwzvQln74pdfmUBeIvq5WgK8cVaa4D4vX11JTybxmjD2Qrw9Caw/9pRhRCp+cO6
h9Z0l3SRcYLEM0L9v1gCDFaU7TMZHcRXCDZrg3yM+7gsXbpc+JVbaiQWm6VFLXSw
kLZKWgl4qT0cZ9ww8nDry2TPeZZwa0zfaO8na3DN+Lc6tVWe5VnqmS+Ar4Vux8lE
9zyq5z9b2fHD89bfho51SMRzmh/PDbhTOX/ZgPwyUWXMu2hRVeYnN3uLMyvhRGZP
sHJ8G6biE6kJxTIbmlMfJPFAdHKvRledw7FZu2vLMkXUHrUF9ebS1emdac+/r/+E
VzOkDLvpWfWpunh6uTu7zEoY7QCEhzQEgHKVRFYiVbvAqMZID0ZcKB80O6rbpnvp
G1SSVqK2GkbGQWLF5AmFPppo14zjXU2rR4NabULwlp3HRTMJ9mKDA/MI3apciXCJ
bphZVNVtUbV+cFLPU//9q/xEf9YzC6N2lVBkQep5pIvrUHxUODxPWTIuddDWAKZU
U/tu29Cz8TzQ5JUsHxCo+aHO98AwMfNs8s7W1ZzRUVgWc4XMNMpJqMdIYEG7Oioy
zV+iusooL3LZZ2/6LEsJQjCT52Fxjx4rplXtfES5Jjwxc0UebnY9UR0CxjugGibp
EZWPavN1X3taryvyZFzoRKSBTSQJmatJQ6rGuSsJjhhCP2+PLbU9vToPN2H9pT76
SUulkINT623KiaivDScsHjK/MvmdAp5WxtyQYXqAlsydo7O/5WOB8L1KWgIvzBeD
53FkI6i/bhZicbLqC6thUPi1qwFczbbFWtNDB2XZ91Nv2zMeUI/8z8Y4ECxLWWLF
4dqZ/GNYo51ybj3DO1NEE3KW7Kd0iegLCku1ETYKYF+oDCajvKA9XCkaEbrqWamp
OiUNGRo0A7K17JACIqkIqZ600YKeruE6o/KLCpzaZkk0xQ3e2xWfNsbxdA79n/j3
iDBqat6gw3dIS0GQKGZi5HklJ14892yP2JsfQ5/Tr9mzWJV2XreRqx8JxeA2EwpT
9OwBbvkaEOPtOXSZlfQn3VgvHY3qx/zxD6acagrEBL+k1gaqbi9i/CeWHGp36n6N
2bzbNcA3zAwizvTKIZeCPZBAm2F8jJazzRJ2cvOgZRH/1pzTTNv5/UbTsl/h+wu4
FjqtOQuify7+Yhd9NY5kr6keDi/AduxA72f/mZfQFB9psZmJ+0aKLsMAAzqMn71W
pavDc7GTswUHxZXVOx/d/Etcvhr/RqmCL5ARr9iOxQopoKMOqxrLp/xkvqkVT0+3
rdRo5DaLsYpcXjb32TfqjIFo9Had8s90pQt8UwTVPUIFJLH8lE1noOy5zO1n+yAj
CIr1X+0FxQXnyjiWb8g1R9dCyrzE7ZWF/wvrwjByp2fFRI+ZjSym5bbHFr+glYij
4h/pqK6xT9SkURvoXxPbuhzV8Y8jQQWyyHOyi937TuiR/Vw9ErFiRrAMPgo8GAY6
kkh/GpAIdrmTPCeY2Ni7KJg/uyqWp9cuF+8S4RbVc2LpKYSZwbh/TwjaGllWs+AX
v8V8kPBnPCZ6gP8onK03tJdRa+CV/kafF5j4/yldtg/X71epnrVBX5Uv7vfa5OWL
ezNDLSYZO7OuoaiYSAeJvAGp/RcI+mgSq/XCXpeEUmrOOUJ184cgTt3PsvtsXozW
2OjtHcqAPdBcWlWcSozGS2vMogT3UYfCAi+wJbvuCbV71kLEfIMdaOPxQBEouMAh
hBSPrN6ObU7QcKuCRzICT54MQxlOo0I1DRZ/Ia8LDg0JD23zkr0iV4m6izcdde9Y
CokRZH6V+wAUSiEIsywduTpAnfZUPKukL8Z/i4B8DnxOjKHJyuFu1URmJB1YcJ9Z
9OJFrgA0vXMEAej/XkmMXY/lQD1ggwhMoLQv/PTei8w4nfLTN4paHu9EsnMKC1je
rUsTOtzmKvvJ/OC6dJkM/qO9N3DUpbRBBg3QegBSnqBwxzQT0aC5xK8uSoMlDobC
1G6ePE+dr/LmYUCX37qBDxw5vZPM4iy7ow0+mJLM2nyMYa5JHSmL6sXQHz0BpZaU
xs9zoqRcMRt0fkJXL8d4sEmBY+l6rFwJTFzJDeCfI66YwLBlb/Kvl6dhFJ2AF939
F9SqAWbu8Rd0Pt1qzq3nKoiwbY9Fz+ue0GYS1T1nO4lndFMWxs3lgn+H6hY2wg0e
+4IKqkzt/10ThFEkppDUUC3Fuc+t8e6VA7yLTztIptQL4YSv3ZNIud5f6EH1Sf/0
3MB+Ktkq8RUIzwR6zSWzYEk9+xQqv81MpPA8ucmfn1/tBwQLpMzzcpQYXs+0uGEk
0OqenPRAVRbpl17+FftbUu1blNfIOfoJhbaZpghjvmp20BYecuNiegjbQBuMSCQE
pl9fikGirkJU3rgUJB/O1GZZ6Ud7w9PNRSPTJI4z5aHd7Q1kUj/CO39vyIONxaS6
LvpGjizbIlYf3ZRVKn44x3f69woO4FFCWzhwLBJ4D9huxOGI3bO9X51UWNVtCXVo
Vm9s6aYxpR9stSuWc7A8CCfJUGywGTXo5KTXanpx+k4QFqWOpzwqfcKckDUQFEoj
Z4kwiCM8yicOaWcoI8C3kpsIeBJ/3tsamYFqxk9QQ4Gwg94OfStdcCCG5M82ANQb
daA/UbhyQFrRlgSgsCMa5wvFvS4dPX1dDXL9KDA8VktdOl5I8PpXvQbwJDOgyg93
jvv1vk8LJwdhp60SqOycvGUxJQOuPBVPlKt+nGysgTgfANiiDHsGFrZ1Uc6SNqX4
l2ox7B/ku8l2CTsergyCHFOvrYrBRLJZCdlttD9V+muPVYf9MP63e8lv4EYssHSA
WhsT0zgIeSrnQsge632bBCLzk+CepFyq74O/OrUcE9uKQYFD40DTfTq65VEsCW0N
mi0wBhpU7J8o2kYmQXunwmEEsYG0cUkuCymdtMbpT20m41KPTCwNaOzgRHO73oLu
UV3MSqZzyJZ58hV+wSWk0yY6k3YMxovCEu/RlCn4BajRLc42FcQ5tbqu4ThuG4hT
VBXq5Xe3EXjqBADA/HCep6U0MW2xCcOyXw9djkkbUXEeQm0/YXeYeC9ug+4JpmUp
9UGtTz4GzvgR1SNoik8gRGmPGaY7ZHTgItohYDX2EyUzjw4uFAB3oGu2OpiRWcLK
ZP5N70l38dDBTf5Coq6bvnKpF/X4mrcOapasu2hp6RNzOlOKBJKd+bJ0ujDLw48k
NoKzs6e5RTJu1P6a4mMH4g9aAfNiyfPKFPDKIpCb7QPdMiOwea2L0wvzXYb745Ur
1E7xXq7/58JGJNFUZ+K7mAs04EB6HMFlyr5YUhI8UWu6b8Ak6fCFR1fAg13e/F64
6Jqh1WAlRLafvDq61AyHNDAOvKCH78xstgonLw+WDd2Va7bm/znNXFzSYNYVJmzn
7nkZ5pz6/EwnljRhWNIVW2Q2R6Wz1LzykaTvJ2pzX1PV9Fb6/SGO11gNa5+O0aZb
AiV26o9RcUbXglxWCe5mzyXZF8jvbPH0GIw0kttYCYSODqinrNZ1rfK0LRlkA5eD
Pesd9AxThMjHfLnJJCVqJ/5CNyKZD0AHwRQpiqmCMXTNc7CktHFkRBIMoEDSUOr/
Jc/gMyd4sCXgViFEe9/SrUZ88JToEB9WJZEAZgqR++rvlUH1zj88DV2dXqGAzQUf
VaTRDyALAa2gsp7JBhQT3cp1mA/l8zlRDqfmn9v0Ay2R5wVCgVqCIuh1iub928em
/FkbWZlNeoVayPM4CjP9E7hpiG5HjeOXKs7PylOSCl3J3ZMQYtzLbFjimTrg8q4z
jyFfPXO1w3ZvRtlaZfKAVST8I9zOt99ihWVmGUhRAod19degY/BoDE6WRTr0LjQc
qKgXeQDYlldXaDyoLS+pooS/yRst6dFoIr9i7lIpC+tWT1Ydq/zl3fYk1qfw03YS
UZqXaWIjLzMlj0xvnAFb/nTKsYftD0Z9Wa9lphuoI9g9tSNVz5QfBy7FlkROTKXW
+Lteex88eW2hBivoYgruk9OaDn0+k0tt7aqWNTlmy6osmQ3/PCoSAg7aec6DEGyn
Ye+yMNxEezeUPZOXmjfPDYHnmyb7lAfL/xtXu0rmgmKHa26K/sroGHNJTGYjrsuH
hOcDVPHdT+BR7LvkDVkdvxtOjBQ5HDDdxtMlsL0kRxpnYaCX3+PIAINJD9dVl2ca
fxre0bu76Vd+MxAHSjC1wVfJSSXNjAQUpyThusAd5SQGxXIhDlzaI2XTcKCRVG/X
lEeGB0fLKpQ4PWLWc0t/EplFHspRnZz+WoAf8XNXJwe0EaPPz34xXdAtCfn+dfk3
h95S8NvCvGSfC6GmuxQMDexqRPh6jv+HL6TctMRruIPP9buAwhcUaGoZtzUta9Ty
LYxW29FySX2rV1gb7w9U9QNlsxj1y5tojtMh/HJkchmgfCIdzK/un9QcjCn4KSoE
UqxiSA3tv9OGtuJz83MNGD3QMbd/hStwSG46qfEzMQj+eIDbeicTLUicVRgST81B
QPbD8wpI4Yc/ytzbXcPHspC/ckRu9GGUnzcvAkKZM1t6KaiYxzHGf6EbeUBTbH7J
lPoexigQk/3zDP8k3fv9/UMkCs6ZLsZex5m4JKLcF+RYpZRSdCkOj6rM86KCgUwG
TTs+iWD8EVu/C2rORaqlmmDYii2djs+uzcGzVZv9XyTbF9t/2EdfRYHtdjafsDjX
GEvhOwd+/vVwy4UOxpafiE16+Eolj7hiucgnMRZdHUi4uVs2bMM4gh3rZqL7Dw9R
V9iewRJzgmnXf7VzLxOtKcCtrnzrtBm0JUCzktt9aC+FPMbmGKh9JszRf79NhaFX
XvIpOwv1P5btyagk3Rh9SLEL4lBEAEUFonHgWId9fzHDFAS9QXJ6cXWYiKUALRlO
93CBSw3d0wk+MKGtmnU8oLxEDBMShnvUBn4MrtPEmpsAbUBTcyrIAuEqF4Ou0h7z
sZkpLmUkBo9FApA6cXlqv74A3kFsdU+X/oV9F8fuAab7etr9eDGAvnePj3tBH1UK
NTsOlSaz4v0fRUY6tn0rl1c5DgPnc9cgIWn6WHVuf5lPudg6x6Z7f7mrwuxruWb/
24ArALWiCIze4+iWaTT52aGRmEovkc8bKg3g+hZxBAqWG4nSrmHPiKadgpl185bk
MSFyBQ8hf1SkRku2jb28gPGWEFcOMtlSnUmgiGNKKjiO9pT8wCoM8c4HhwxAghn4
kbLIl1FwEvRtiyJWOYiDDZ6twB7ohlJPyM7nscyKrj2l/Dt0D4b3aM5kLZKPSQZp
4yn94VRTekD6ohJ6sYmrcufzHbBdk01Q1C0pXyWUTTXhT1xIhd9pYg4NORDhwZDZ
k0qUiArVY+HEbzFQOuxrRTUzb0XZRpkLb3/UwDuetym2exyImTmzQOvapUmOxp9G
ZStckz6kJ75VG/tTHqjx7K1YQ0vwUi0CY0S9lsVhQywGtoelSSGW70JqU4w7zLYi
4vQcyzrapIBZgYr2tg1JERehQO/n8HhPaN4xnPlU6f31utfcghRzYDJ10HtYls32
0sdit9LaV8eQOaD7d94XSCxuYMCmXRlUvc4AJHT7oPufUdetAqGqZpgLm8mRDCVY
ufpIH7znrN+fPg8IXyc/oLpG+UZMPhJNBYuiGN+vsPkLUDFHRtkLBSM0C8v28nQV
N/SCscqPIGi9Wkxi4yySgEex9yiCMp8GTiRlceEQE0vxX/r6+Ce0wBzYcKQYIJXr
0XHto6d6yziCHfmezCfxph+emWo/YKKwvO0Jgzvzy6YDptlaegGjK0+5u+1b1mVP
Xj+wgnhZ1rwM28YsR0AB9Lc2iBEGH8/sIlU84eT/kMiZiGr2kg4G67Vxcqpgo2eh
6EQ3hygByu5Ct/DtFUqNupOE0/28hb1wzyzy+XBNxOTvj69BDMJk+phyHWdiJtNM
bXZXNBsquy3aUpQycynqMMfSEnMTAS4jhT7mka7KqM7jhXqeQY0TwmvEPXY/TOYR
NYnd1IW3fQ89L/6r6eKjLjYDGXzqUBf888qIHNkEMhT8SMSP6fJehRxVAv1Si5Cv
tPq8TzNiu3B/9XqMh8X8P0xD27OohaKukDBnGyvHoIZy/3HDQ9N3bBESn73sYocy
M7s1RFSLR1VKtYPt1gxGokvnyCkeA/sapmp8z4bABvcKFmLWiEBBECdzf/ewDr/S
Sv0oiuLTNL1muorJeRB08NaIPeO5BxfULF8i6uJpt6Bm6cJW03dWSVMXUfZTU5W4
+LZ3hIVtxt7qJ8OcjdXJMSFZwqPzFbbCheEdX8OPPh1LSrM8yRfp3vCXNg6U4OJt
tpsoEBVhPI8V8hxk5Rm9uoXNj1/DcKxgsklW8u2JWdi7c2WHJgb8KgdhVxbWmCly
3vOcjQAxnCHwOPbHyfADWITqvZDFqWiEkKlvrkCAMjOMAHs9OEEe4bO3YkUv9dc/
gQvIuvTLBE8i8yDAtrN2HVSiXG+WnIaXT8tBiHS2t1QMD3WThjfDe0hOYCzzIptG
hW5OArkvzf6OPAR3jTGlSZiWYj6XJSWvOPpoD+YUOEpxartJzdTspj+JEmjPj2uR
67njwHu/9dCh+29CzCHdT/pZoqsU6KpDtgKjJz3ixiHTBOOSJ911e1WUJHnDqpZ2
p7j6GPE7E6IhwmLcCqB0wFQ1LHkVZTfMoXyIauU8g4PZx/XEB3sPyUt1nQDXe1Zn
y4UuaKKki51NlZswd/iVxZOIGrJ78g3QB/RIKvYGJ3WshOLsXkmCwqP3Yn2jnj6q
j4wRHe0n/t/GCeTaIotYJaXDQZkCM52oC5xW2Sl53Y3pzBYSdN2OTjijYFjk9VQm
gAT9ysLFmbdg/xX3zrVqgmsZmVhBGEXONfVPiR7SxuVIsK4FmeTDkDlutu5C7Cp8
bkzcbB2aTGbPuOmzkXKgtQEh0rqq5QG22afAxPj9vL3udwV04wW+TiXpcsDotL19
vvMzUTCsNWiBVxQEtnGgmFu38fc2TZjW1ZMjWuKS6i1tUaNJZtugGZDbuwc00WL1
E1+znb73NtUHNVYC+JayW2cw63RexwA+xLWBCnwoA1mZkBFLVEzbZSJIUBD53XC9
GgcuzFgZfgRKLvPvMLHCufyx/3RwQScj24RYvohG1PFlx5Q5+wHcuYGzCgTwGSFR
a9Z4xDjWxC1GxFIhQyK5V10DKdfMQdljZDFTgk9y5rRLD3Ch2tJCIzLqW47vjdDP
F5mt+Xyg2vn+M73gMjObvoajgNzsrdzAjAPEgSayij5O5DeiOj9zzDBM+0wteKK5
8ljPFLAm5KLjFLhBP0QnkCr5mkdKGNwNJNkjBcxtJBvi4CPe1T9ooZScM5gTVU7b
prh6SdBwRug34Mgqqxcbs6+WI90en9jzFZH+aRFjzZMpGbr5DhkMr6xf4xlooCUp
kYU9KdNw5onGXKYZtNfW9+PrS196eHftD+OhYzTx7pT62ZG0UL+ZkZNARUYfQbnN
689PZa7ErUCWotTtDCccYOo/czwZtBmk64K6fc9ApfiFM3QPQPTYVWTNzhqxTvK0
qGpdV5H6rGLdRHLp9bGiIe420/lBLsy58A07CjlNvSFb/se6pOolsSvRxPOQ9x58
qmAykI0qqftBa/e2CmowDEpW4TkhHVslnNHI04NU0qc4jPdBhfMSHWBej0sJscC3
yfmU2Ql86fh11RTLlf34EDZuG8MrpTTTvgKCOrI7Wfwn/QYo2k1g2k07+F6Nd7ca
4cwoQQxI0v6eQehDLuHbFUMNg3ZNa3htSRpkmnIlghacuLu0GLgVWUaIbwg3SkzJ
rckTEkxvTie7S0wWNLSXG+T8cvVVunD29f3D3q++rgywClZDtRsZJh/TiZVr5Yvg
GIgpNYOjWsC494zgAXbk7mi4/x1vM35Um2MbrXkMvpE8DbcvUQUJOZLq+3beApZo
m/SXhQrV9Pf09f+4nTgTsIrlq5goJSIsKWIAVCZhbxtW8EwMtxMLLQzdZ8hspm0W
bPKHvCXpqSjYGfOwrh36cYm0VX1Lz0+2R71zqYufmTHJh1P+qdHdVCin3KMmgtgs
T02EJG6OHjlFqtqkWi8TWSWWMqwq3mdFeRQwMdFCDUU49Wg5N8t9tjjN2IXRPcri
VolzV7K9EjSiRoW/THbjP3ev4HWn5pWKlaUdzdUGyAqyIbJfT2ysZWPKbo51av25
FA95AEf+J0RnuS2u3sSeqCxEW2hHnTW9jFs9E31JdazWPSBPDQCl3nlXJpMqpIax
qB2fUK/SBIrlnIcJwV+q88XOOKIYv++oUueFyoSDu+FcYoDzEEIiU3GvuKSVqQHM
8qu5nBebpwGxH5MZtJ+U46/SpgGQrfGqO6ZPkFfyVuJtlTDOOzkrRT/nu7Xlt3q3
zwM0H2of9wEFrXVB7Te24D8hMCH5GwRRranpS6lo0ySPyDHk6HVaMuAn9Ij0AMOQ
oKHsbagooTjZ9NBFxBjK0vcIQPd8/FhUsispUVNKrFTPEhm1qUFOr0//OAeUm+xC
1mSSjG7V9ad+Y4UCaTUZN0/Bz/pzDiMV11RheZUfXyS1y0cb9hKQXEvpzAbu/RYP
k33hd9PWX++e0WDnsShDhoSDOSXpAxvVwBEUc9adFGXTc7+cBoeEZZT7DfZso/aO
JF6qvixcbkuNZ9PyIQdXJ/ir4yV0smEpHD5bQ69QBRc9/gKXNmBsYVFAamYuoUTX
VFMnDcekQgc+wVGF76Q+gs8K/kN5muSMZ1My1jPNiIDo1iCQ/Lj1Vxc8AQCnEd/f
uriYt9gQNRu3sjdaQUdfGXh+WbOpAk6tkOxdyKxAkMsP/pTV5j38DHqq0bsuC+6b
Cw31TnwBZ971vuZgdqOUskJHpx9B6OLfhp34TOwPKhprsjxNjTbxs/RYCHN95FO7
Ssv7dPJnA5x0pQ/F+t7QYJnquA2og3yt99ReZwvxaBGSmwhX87/f0l8hfCgFopkU
itgTUoqs5B1zndfXRO2xez8wAjQnvrnEsOboZROdvkFRpFr0btfCwAtHlEeW5iwL
kffcuwkiutAB2ttanOpC8wu6p0rBQzmg4K5r3mMDD5KVPoK4+1TtTv3hkBS+m3Bw
WitkZMTewHPlNhRSWGS1jqrjhUksqB6x4MktbHMzVFOEgiILjaHW868D4OTtu74c
IJAJGwHI/py35B25Ag5zDf1GimIraWbV5infhP6Cp4Ufiud2POmEVgdGkt7dgLhN
rBH4KHC1uG+p8Q72+hu0MsCciXuxcjWzIDbKBAulpznBOLDCqBeEPHTTFSMvih04
sieQ6J1M/j0HUoClgY2QNHoT71Ai5UJnOkdECM7jQkcO9HMVOZZZHFbAjEsObxc4
CzTtZWCkF0yRW5aqVyAp2ZBFJntyH4CxPNA3GWlK/2b0eTRzmjruu8WVLwytdvqu
43jddB4uP4MiHbf6tQMvTDhCyGLb98ArSBEtMf+Ilxbt+x6OE3HlQ77Z53OHmh9S
WglRg9piJSYsPKJJ0vYzk5MD/keuWIME9dO9DNJTj7/4olzZAPA3MBpkswFvWWUG
LRi0s2+HYkYlge4JHrfrBVhd3NcH7GA7GrPMgW0+qQMef989OvhtO1GwrVDCvvu2
ehyD94iKWOQkpqRaIT72Z1QE9sJypaNSmvhs2uvznA9++CLX1L/9Bzu8sRvkIEGt
IJSuS/bmkrbbsEKsbhegOZvRS0e6slYTD9PXDjySF/8rQSZKwIdiMdHMBK/6tKU3
Sgej1tm7WyINt62r8OUee0+exoYlsh+eq4y3dLpvyktIoVIVev9825+72xmqhzj6
iFlCZ1EX2Bn67nPhyPzBloKCfR2JBWkaVWNCGmAhfZMt5qwpU2os5kwpxQP5Uv/N
kUpf5iEewbEWlTSMR+umpJnE2PAbnJu5JvcePiiPrvP92crxHAttxDva8HYaz5O8
CPVqPog/tv0bvEcFtT9F/nZRiD0Pjf3ovS0TimUr9w7K9HRmKD7SIkOQTbVOvSIb
QXIqHSohpi2ZpuxAfMRXB/fhnI03soWE5yzcfvt72FqQueS8RFqxBKQ2sDZAr8Xl
Had97YgiHsYHlDg/DrbeW6GTzRY882ojqjw8pLW79Iuw9fW67heaYMO8Nyf7BIPB
rNTnrsSiFsDyjW9OQJyTSslfJw7VPqLjks7ra3f9PPM/crBgzW18TBZDUpvUu+7c
XRKKjsvSW5ugCzqrqUq2bP8aDUBh9/Ino/Hzt9e4VMTY6RkHOvvwKpBZyXqJpzt9
BX1kwmpXGT0qUKDcxcV6jYmbe2KIUCBt+VE6LtwJH2LNFxJFJSPtzukk/I3J/LGG
J9axQShUJlBb/fuTqDRDIq9xMXNJpY4AV0h1K7jBRCATySFrggwAugioWDgFhb3p
E0NfdEzyDoUJjQ693Hb1soSP0BEVwqKkhNCvhg68OWqD5ROu1/BblL8vKERVF5Mk
WGCxLD0JQb+Bfmc9VlAgj7QnnqbU5nQ2ayvLmgToimGvGiqMpQ3GB5fBs+X5YjX3
OYtazVa73rkyyB3s/ztLYVsZPhzzVa1IUSuMUdzVL5ngZOHZ9mcGK8IWPBhokg0Q
MdmVguUkVhVJr/8SXWGOoKd3KgEI8SVGHpTL5kzQy6NeHEsjMPEilIe0FDPRPI50
aWKNZOI1IZe+DwnwAj1hR9FpJ/jC40CcOF9QeQmPay5d795t08d+ZNST83p1HHP7
IGzhu62rPcok2z4JkBsYJMjDjztldE4ZxGvcCvhp7yWMAvvJ2GJHNK3/7AwK1YUv
yk9tyfZ1T7XudpS8XGdb6wmvlQt8feXVRk7PCuUmWJNVVUDUN3Tl/DKs1dgB+NXX
SMa2I40rNwf2goaZYb6lmpBmLCCEjAWoeblc9xXv75OYA8XJA862kfpd1mr2piJ7
spwMLdU6NYKvC+GUi5ZCl5MtRk/LDoEwIe1iW7cnrmgD6G3vCvRKO/sYRhYt+c/n
JVDArQ35G+CaVDQ9OPh2V3JCOH0aohIM0Zd0+T1LhMmWSz5/sbhOkW/uDYTdDPFN
7N8R7U64TW3ex03Llhvztm29Nc0R5yu4ZXrjKWhZoJYS9Wo+2scV0qpyNqjIrIOg
sznmUmQLakCbeTQuaYYI4o1lZ7KMCKwNlVhs3A8UJ7JbQmRMGAl0uv/dKCG6vic3
bWTcTCfVSJRJPldqRrWd+Vin3sfaKF0Z2KrAeHMlBuN5EPdNnGgFA12MD+PlJJBi
RhkId587NLNF/4k/OQfYNYQ0Odhg2EN7jAjBg+TpVDD+3eWWuHXXzHhu/9pEub1v
vJVj/bKMluaJkhp/P1pDUTFjhWR3GD3D+StpNmwa1Bd9lDcCRCRDrogAQrDDRjxY
DGKpOlLCaMhT1abg6sbDo/kNGKmbsJy4nqK/Ji08BQmPOu3zW2+8jUNCTv84ccbV
vKz5N6EZy8vZG0tygORBJuFomksX+fBY78tYiDW8SPqdQaOXoXwt5F5ezWtDZbw1
WbNGj86BRYPsGN81InrtO3WOOLq3VPO1kQ//LczMHnSquEz79N4aQUQuSp7NXpKX
axYnshl2xgmB1YwXGkMD9fa5mOwyYyrGD5YroRZGwHVwFNRR9jdBMQfJEuoaD8hV
Gucnb4yVGPA1L1I4aAMdHg4rqEP1Y+qxB+GZvAZNqnTo47yJ3YE3Plt8Tz+34Cr+
9tLniJXfikLgYRCBAgtqEBxtunpBbuwrTFLAatJot3gYw1Y8aHz+XAAK8y1wg48e
s7du+lxKQo6umsR9fTyj3Sw2aLSMfVWWi8FSzysf3bjSax1QXxN/QcSG/bfHT78Q
o0cOwHEzMJGq0AFtq1SfBxHqwmr4GSgzXiv1EZG6DQboy3T7ev2tYAKgl2lPPubN
U6eenRrl1IFreulR8p+zQEKlkYzQBCr5ZU6ubuyxNgcPo+O4CMfOn1918hXPccqM
4wtra+WOlgliqp6/Y4zNXgkkEfMrLnl8DfsqLz+1URMkZ9gh1EJA/DZKB+bHb5yN
vHAsi72ItSnmA+YLVYQ586lNdEkkBkh9VT8loxH+uuKiefZkevxqf4PH64KBc6Hp
s0Gr0lWlIEIZ3g1pF6Yo6f3WFmuQ0nx4yx9CqHsQDQ3a8GuP9oA8hQ6nIDZ7son9
G0Ap9l7w4U0TC7o1sdUz+Ioxnh3TZ9ZD5u3lu9WDBMhfVB19jsLe95B2oiZ8Aa5F
NWG1AurDWZuUQtSJvUyl5RtB9kQcjGkdpoUosmYhsdpPjpPnGzIcaUewdJCYRuL9
XFuPh/doZE+cTWhXKdmNeaCmMHMjojkp0Y2p/E1e9FD3h0wI9sReKdzyYk7osL3z
HUjXNz/6cu/zpeIUBs4te+1rwEXgQmtY1l4iy56WNGHQOrePJutgM0c+Pu7owJA/
sYPmWkBLWezGspjwHbwGKj7QGQFzRihDrNYJDPCcyQZYv7PUGLj51YjHj0lT59OS
qDYF5RN7TSKWsa9s3R8rNOtHI2yxXy8cd4E76+TozFcZgW5sUJBQ0DMrTLYoOSkJ
96UXoEWodWW1imjLSQL62esI9eyA4ifzRo3kqkgjZJKVnZlpF8z4ixE++IoD7Was
4fwh9hH12yc5B64hEu+f+v5sVJnPi4Gn2uiY3orexBoIo9qoYbXThRF35Q409yEp
Xm/1wrBRupzF8GzQckKsfY6wZCS0ljRJWZwLjQvQRbHdYLOFanvpZCKTdH97gX6s
czynAkyu+I0eNrhH2+cTjX5HtQwF4Ap8viFtRJU7Csifs1VOsHq/kAjpoVVrzA7z
GNjq2u2Nui/7LUa9Ad7pao6cKDz8bT0/W7Ss4ky5sZcqEtaNapvqVGmilzyp6zRp
/DP438vCIQKptJvP6b/iiGdXvOlPVkwzQIq/bt6tnLE3gyAJHWU1F7q9kPUshp3t
tWSxLonICPa+DR8ivKA7TlqLdNRzheTnp2nVcgpe54kAr1glV26njvcKIWE8j7XQ
UJGZtk58yjIf4IAQIty2X48bmp97+PE+ymTsKXclvqh+uubpFOtPciooUtiUfgWF
RvdHhK376NPPCyOtMyXdrpnxJte51UmbDsqYd2MPIT1BgWxpzwwG8i9JmBPhfh7I
VsgewK3olp7k/5h5mmXec8huNFp5tVClatx8ZQYChFjuPI3vfrCfLPOqPct29t/6
ah+LfdaSek7c4x/KUtqLbDOzAeGxJmIDzksqGVLlIfPvcsksebnS1gzKXztUf1FU
RWpygnZ2m5vmoX8yoWuXm3h8Dg25XOZjr1IzdS6X33dlfSKw5JYUwsHxPuojfMpv
IdCYDyKpj7MguZyYIx+tqKE+TVt/GIbomxkZCMqv1DQ28U4oASyY55NZFG8X35ew
immYrEFHHFtRGR9lMV+JbRBYdp+oKWWk+s8bpnP6bES2YS2bykGbsgO5zKJ3qH79
XrC+mg3D+3xDrvuEkM/vMDLzSr9lUirF+a2asOF3xv08Zw3Nmx5IzlE8VD8dZKgy
QDWuvZrbm30LV6KGC/Ht53TgEU1yuC8jBZoFuayX1BhrhsRrpCWicxev3O9mmWxr
5C4OhkoSuqPizwWczVBdvnI9d6dDbx7B6/G9vAx2a3fkLXkQ146GBMz9XhTvLbCS
at2qjiZTN9oS97jDmYOTS5q/laXbnuM/71JodRCz799vyCCKsqbmH2mQbj6y6ASu
zTyvOeIB2WNcdfmcM/y8VddB66eR8izaLcApgV9/K8fg5joLygthMNOw4+skbVS/
O5FQuxEPh5At0PVxD0xmfgF21foQxYG8tttyeDxduMQUfD3cCbaYWtnmyciDsXcK
fNIu97yiVQXiGip5u0+LLIScL023TD5FpbD7KeWF4Kfk6eYfTLJvlfZFVNX9Olrc
Uz/P421ZTnKeSoGZdiaKqdxwH+3T9cpL+MT8rvJjMhnjYYXaPYbREGg7kZn6Av20
CXupCMGqpF3v18KaUxBxNxy7sYOwXwxLOdT75B0KNAdcYewXxTQcz+n9RDU7yniF
YurHlbNuwf8zTkcJ09jk7CZZ8XPuVLDOj5KA4jtUZBwrKE6tBmGrAgz3rA7UAX15
ByHUb9/lGdRr0XH6umK3/UFhGPvCduA+tzz2GKFsMSl5zojpeiZZTbWRyliZkDqc
z09b4py/jDCCrMZ10vm8OYNgtAnip9r3UWIJvp5ofrcErf8VJ/0TTHGKAtQ9C3Ni
H6muqQCoJ9cHh2SNvzp09IaA+Zm/snynvA/MVmg2FjYkZG/oZpv0wzZFImWxj1sX
y5hii/UCt6zdVO+RN7O7ri2s3XqKRGEp0SjLhfbifqWL9PNJE52N3AO3v/UKyaHe
y4EHBxF78lacEpFMcJ7+Cltv2VC/GhQfbHpRJACinYjAQcF78NEtIsXlsSrOpPx1
YwYQTcR7oXaCkD3Qbqswl//RO4kAfAKuCb0bEXGOs3J0hOP6gAnLE9/N0AtUodSB
aR9HKcMdUatdcAl18/rZZjw4ZZbNaoXS7KBeqRATGL2uJoTxP9Il1lPf7vzMVlC9
PAUZC0Czhuz79L7vd7YNQ4oSxg3aBnxTUvWQQGnYjU6lCxk7y1TZ04G3CnEdbMNv
+QAVvi1vv7RGjp/PtefIVwOoOO0ff8oRo8E9Nu9rpyoD07/XfVYVoEq15WXBaqrh
5kAj/lrUZBbDjtmshVl/osFrDBxNh/CE6mgZBJqkzB+sj0UPpPctlnX2/ecz0KwL
el2voQAn5ky0QKplNnWswEqNTtahZhHXqp5oXoCrgV0RhrywanSuRE8ky5Vq2MXX
QjwtPBDVNDbfdeugwwIpmYxtOzMIZrZZLG9FFFuqYrjL50vJTpK8E+AbSkpzjbur
f/Tl7+gtS50YSdOoUJdK5VPwMeZCpIRDGKMTzH45x3jzSwRA0hwLt/sbD7MrwJJC
Bma0UWAgaRC1O0n6XWekxzyAiMRc21BwNeWQ/cjefakNt3vSAIk7BC4FXfQ/Wqaf
wE6qumb+QXKVDbh+jdQfLW8KpSgh5n8pM2uSYW8xMocBckNYX1cJkYLMp7C85DN9
4WFDxQmoS9xvFqZ50w5A+0AXJ8n3sV4XsJyoXP2HfxedJf5+bSNAHMiYGeBnJEtP
UCED+V7T+YgfOqQM+WH/yvqRnja0eJifNUbHjdDaYJHk8sjAuuvIYObC6Tfl3t/L
ycP7Wj+3xPAB4krjG4N3Ar9vdmzrUNVckC61Nwf3ViBZ5aj02WtB3hWi66RAQJBT
s9YDIkd0Wkh781qX2dWTyxiRcTiF1zEpiJ5pRNP3YvSYVgdZaxYbixV5tc0viXcx
7uizatCSRGMHBiuxfly1KUOmm6Dd2fStD4HFoS2FWJt3AU3w6qnEi6vK2oLU0AA2
EORY7v48b972+Ij6iR8ewKjEQxMjaNKeI+pwCFaV0Sx1vokNGauWetIPrR8b3YQp
CvCERHREsEqnh+FK7b+G2Ab2r51RYFcwN9iXNwFMJGMJi3HzsJiwJwLcrtEYLai8
+O2fKxs8USnGGubFjQjUZy8AAzMfmQ6IbC/tL8BlNIMDAx7fhU/2pun/D80JRy82
yMEJEqObOddKeUKwRm22eIVhGEtGk6yd18Hs8DOZrbnrBXlWprK8bDFVjtMUp2aT
NpzlkyZ5StKlzNZDeiZjt+K7tABI87ueLCO6wSzUTGL+gOapwOHAylAkxiGrCrjS
f9XSI7ai8f0ZPE2GpZuuBMk1NKCJBykey1zDlK8WNGytTIcnwR8yWxoCytb45D+C
7EFicnwV3T7qLsrmRv8SRF+tpnO4Tu6MgHmMP6DTUexqTw9BEnkwuBp6DKmIbwin
oFsJSOHB7ryek+GU+bsfx3hyBMMkgcdhe7bYPruw+K2Q32+z561sp0s8ESNNZ2qD
HJMQG04q5ZCrjrS88cyBWY4pum1Jl4d2Xzy7H1I22AJZ0T03LgGAzRf/nR04NbjS
YGkDj/ZuwxrlEdPpYVdI1nJCtrB+/m+9RG4Jjtjo6uLZCkCZVcPLwSQb30Rfgylp
U76Bp+gEBqHNIfvqdsJB1M5As1CfxeT4iU8oBKYgI1nxfUYa8GW2OED11HVDa7Z6
Z7g08H0MPFsXNLcphddTGtMz0gzEDvwM9XjFOnClWWt6P0BuvJ3muGS7QU7fU4Je
yCkAyaBpHO17Yh1TCdVLaZUcVIK07ZjwPE1VCVyuLQp5ZBuNMS73FF1xVZNa1iJ1
2rzyF7B3uHpxvvWnV/vrMccMy7JNeJ/1TG2Bhh33riHmM31a3DQEcv4HwB4x8qYb
tI9ppL5nhH5JFkaBmt+iJk5rwk4H8NLUcWxuhTtkWbMqSxR1XlEIWa5hLQglGbvu
xlKXfhl2UenUj4lFoCBx9TyG6mIkG4aFEah1SsrJIz/rvgABvkdtXE+4WkCSSJfl
62f4ME1cHcP7exI9ws5fvYbv96PM+nQpyD5ttyoJg67dLRUebHcNMYM7Qv0XvUbD
PJojNFb8ohuDsYGe7oHRqa8FTGVyaf2jooh1YEmAH5uUlRs7H+8r4x9isoGXMtLo
U9TknWbg04J2Ri7hgSFcHYVypgxMZarMzwExu5rLXOXTQFPv+sjyTYQ1MkP+v/aN
mu//K78M7lK5iUOOTri9mHdaNN2/Jn8zqNFJql8nhN5BKetiv1mc1u9/Q0kDIoUd
XeT+8DbriSn5nE9cOiGF2RmuznbtSgQKPQ2OI5rXB5VhqBb0bphz3Qw23Vnd1LNr
z62Jce4w7OWrHEMJ/FtNgrg57XSNbShjtEsiTGAHdouV6LRbyJtGDheIQQJ2ZVEB
5QE8iUoggyPq5QFwUM+GNkZ2y181NHA/Gkvses5m1NtX28O5LzI2xvTg89K4Vg6W
mqK4WVwqy0gGD8WK5XGiba+J3qu4GX0CL9gPGF1/Ya0EHs8zkjR4ZeQ5+7acf2OM
/deQYpnsCmlFclkVWvLnuvQ4kRlOOj8E5HtZpraYFAoQOFSuYkwVs4GRMMnNGhza
7AGOevdZCue4o1PqeXHyrNV4G7FLx8eEl76p1WOhYKmSsQx8d2vXl+J+vuZ5LTiT
1Hh/OoYXNs+pfAFNZIfGKAEGbM0P2A9Tme8ENLgr9rCVIm1v0VJMPySHrxfX5dgk
YC7cu1FxHe0f9/w9m7KC8Rct7WVQKK8U1VKxoPk93uLL7ASAl2nbn4G2wKsjH/bN
UrudVxRgUPuBAvqF7ibGe5alYTMBnr3bHBIZ2G+srhZHPOXzkhc/uHs6pwi4WiYR
f1cSyDq53B9B5s0iNA6hVdbelcvNS6NBdWNJAnWK9GyxXyvRxez+86yzjpUr30oN
FjccgCb2f/wEBpacgirIEVztd4Nh4FKotU978zykiyaDTo2CL9Fqf6V0ctcf3rtl
ylskHzTx2WrReMJHmpOMp1xlxbPCUDjsv75gj0qq7rXVw3DYEpJgfI/b5wYtUh7o
KfpnVsHFv2Z07Yxe7YMUYVfOKYEXNwVHO5cSMooAwzv3MB2CjDLkfvy7WNf7EGg3
cLEAl90Lz6f2g7imCiwiN5e0ehv5QyTgh6fPAeXy/oP4g924WXyLvIrE6pxDuRev
oLqFYS3m6y3yK6kafjDheq/LiAXRCrUpm6VIoPO4BVK/nwF4VttZgV6LFszRBOvl
7Qf4kyqaKT0h6UQPuyNJms9kJ5JX7lFuEoBS9jPfSXt4wsj+b5bJDrhgkU1Fl0kk
OPYJcNGT9SqdXcSoV+JamOwEw/1gfw+bOnF1aO5s/AAfVI8U9zx7rG733shxE3tf
ksRS5r+O1kyUoznijjO/+j3ZzxAv3ZK/c/QjIPahfFQhapCyAsCBm5eiy8/lAfaP
d8yVq3bjQmcZiQG9825vAJhkaHfWZlYY7/7vfTtW9WTShZoFDQHDZ7fO1ylg+lSJ
u3tugvZ0+Q01VI9mfyizZzG/DrwpZLUkVzMoG5YyLgYBtJ4fMW3tOAd638BWAspJ
sxJbkIoQIGO10PzvwrFwnudbgTkoxfdv5SJ2I6JS9LiWKm3adl4H2P6nzOv9axfa
5SlxINkrcMVtE58KHXGoP86IM6cUSt9DcgdhHFHl5bompeOWuj6BJLAFeyabFZns
uxQrY+6jnP6bVKzsxl8MQkgos3PUX8/zzEGfhGXtfDXs217oUFdVMBSJED1Km9GI
swov/ysqvd87z+d4I2skKsfQJRP3fPxO9ptB9RyJH38L+kA1v3Unmv9GE/4T1kr7
BfpLpQctsnSamA4XVFQJYForaUMm7dOpYrkeh4kHtpR0ByEwB7AwImkUre4qJpga
5rbnf/cyjzi2n4CD+aqKHblj5gTmrU6byrYDig0szA9utm1fh2UXthrusBZeZbQo
Nx1W2yejkFhF84lfkWl759tfQK2AwNjIuR9BnD6/jvUXMKPEa7TpLccZHEXOP20H
3qqmL6KkLfr4ZSdt4CZI9Q9bsiiTRRYZxLqpn36UapwUr52CSNPKBzfjR6oCqmJl
l0QkrVa3svkL/+7Y/b3y0pJauRxVAsVAPrCfOQNhXcO61mBTWf8j81u09p+Rm0Ci
vbHrDozvCfIkkqhapw7GyBuO6ps5JXY1eEY6g1VMg1IE58ZEtaS6TFDp/Kk5TyTw
/lf5nyFmnnceQ6Muyf/fEjKakIXrUgoX95ln3nTbtem7+W/y1aPBOGWeBQdB5iAN
QIHUxdwySXF8cm+qx1VY7CGzaRpynQDYu+s1jVwZ+bZxP4n7gBZpS69tN1Luv+36
KctTE68eC4XfWDUFb/yBB2fm3b1fJ3kawu0G8IieWQ+J2Wf1dg0dnV5XuTustYxs
RsEDpVsoDz4w66nxgI8EifdJ7/WG/cJNM0g+CyhDjRYLHTxFNHXqGBEODxV4pLDA
cYB1lrbn2M6AlydbtFXXZy56fCLWyGHOmbh58QdZEYpRmLCvzH9s2KB/fMxr1XOL
k8moWskbfldh/gKLTAxfM/K/hD3hzFk8y29IEHim54aw82Ysp+FL7K/q7UwUf0++
FyW5w5HQ+Jr5FUvOyjApSnvYnJxyMsHpAkrTnPkSQZLePUzkPnOlKqbn74PLcGLh
t4lGk6CVGY5FY2vM7WFshNFHzLNF4pzOpKcxq+6opIS0vnMl+43/4jRrVW991NcG
AXjWzeNWN8XAtkoA7tvuQOpW0KohtjuFoBuKokY9p2zk6vfy6ggZJgVCv/qWSbyr
S01f/hSd8n+aoM6XHkBCgfjoxGiqRVWDa5JS+f6mGaK1qJE06iaM+LBoNXfwKV6F
Zf1/qpIxhwxJXtfS3jw110d8lT/rH7mIjKIA6hzJ6swJp8/SiLO2KQbyqtIsIkQ1
VqEwgIpUXMjvCnADfyCqQMJYEhr8t7UPHy/EyFzNoqnPS29Sd5KcxWrPBoKUbiqR
xVc0/uk65IOZNwe1kXDVlB+iLRnaNzLNeDDv9UbttzDG3icd6MSi+Xc9lFLJOJGE
hw2CmYN5hOvB4Zgva7rGvY3w/syM5rePUnf+6WwuYxgC0TZxjophaNPPne2NXsMl
mh/ZNmsyxRc3o4iVfNSecTSvOZuDAfLkph1btObFYKuFWprIXVEyBrE2PY4+iFzQ
8o0WhqVwjLYaoN8CAoB50d3tizKGH4neg4JE48mfIKoTkdhD3yHJi3S9FYz30r67
vPIZ+bhauyBvLvBXaMjXSUjmkDFZSEQR9mkjE10n4Jb3nr90cbylyIhHB8KGxGAh
bOT2KwERyZUbBRN0+xbP65oE/DouL78hclISLnapX6yPZK2f5IWq/tsF+jnC2Cc8
o7wgx2g2X4g2XGRCfD8dwQg3nrPzFARhqhy7jtb3Wr3IduoqIGbmR6RSFmGxISR8
BoDiD+C8Ra85WTXrHqS8LO06Rx6MAKT8sp6mO77pyBucrcJaw5u6dIEnK5BQPYWk
vWG38wVbG7yWiosO3gWm33csQSWk2uVmusTD9bja+XFJQ6kjFExehF4gq2ja3kdp
KSp3sN7E6kUuEXIrlHc5joKSs3R1C2xVoXUctcbimSF31eQ4jMpPF1TpflKjTTfj
fVke+NkMJVa4RXpGs/Bb1YVNNlgIOoFmoc6ShxclMkBH9Wpz5XsHiBKryjxrA3L1
MxSSjtT8obCqmwhMV6FodXTGRcGqoE6tWapA5EPWm7HGP2C5GHp/qz4xDwyHjtE2
GnsLIMqY9OUsRWNI7j5OtIumgnB8/a0IiRXzJKghPyHJNEfA9Keit4vaSg5upp7H
GK8wdV4a327Mu57YF9qe2tjr0QaxbfTDCL7EVqFI1TlcpgrXxEUPcFfXIbRA2TFv
U2c5xc1xZpqZ2md7D+JeMA30QjeGrGJjwNrSbRMTV+uTMCpp3lsbzHTctV42ftMF
snbeAMjtT+MjB68ejGFBvv734BueOHu6KC1+1vEklwbD4I6tB+H06uLXdTkkNI8v
VQoubNSOFRhNk+O+JB+Z76nOS2mj+a3HtPre1BpW/1w8Dp+CnROmLZ6ujgr7XHpd
wbwOLDqNdT9JWlciS5K6QkBm5poGavfNbzPB8zZfecWQRw1R39ma8hhH8BQ/rhEi
9CIowXrsOr3rqMmoVlciPPhmCATyGpECevLY56cXWdEOFq3QrE9X3TBOadqNkUXF
vLAlpOQFG8xGM9tAIobITcTMfCns+OZJHiwylH9B3SYLXzH5btqG/VYrdt8ByKl2
UW5vHvgM1zjZ+Qv8gIVMK7qkp62jkb6whOEjuSMf6wFETnemqrga+Dv21sloSI01
0hmkgQ88i3/Mz8tdLM8f0BsH1bHBqEFQMitdGjD/a5342TzLZ+CXYor3bTAeKqck
/txZBwSkPRu3SZAzR4ac1+5Y3MVgFG7mIYknAyvkbOgLjuWr7lQ3PQnPJTpnv8/P
F13y0C+qE8A13uLBcFJumAqYowKZblVz1wiOhboPEHMTtsWOCCNwfM6odmQNjWWK
AxENtf6PMTFe1rZulxkRKUESY4sEnw0Z8l9W4uSu+nig+MAGcs+ILs6nfVhIh9U+
FLd+pzh7fU3B3PYWe84LcTotStWZi+2XLQ7CLVV8Vc7L7HThPRs0XbX+3a1O35sQ
+VQkxnHScmhZKryraMgHRe73LkOZI3SqWy5l/5CgroCgXNYCi1FS8lNChmkrgCgS
8LQPBINFidDknHpxM9OtNnbszrjoH8mknKDJLLzf5bf/MeFg9hepjeKioLp36SNh
21mk0eq7Ak/hFh2xbhU/9F+Ys1bO9tY5jGfnG+Kn/EWgayagskDkNzw4OSvLuvZf
Fii/kMuFU0IQfVcBdPnZJwmP14LVv/53tIV4NWp8TpLmojNx4QbAh1WU3NtOOT3A
KwXUqjb2o8h0MzUc9g6oSzRZbD0iJxCgGop0Atyl1gccNzNXwAmYbKGoH9oFuGoR
6/nL4XN0XAHUt3Qb96MEquYoLGVLSVRQCRgGKFUVqUzDipVs9rNlkowpt1/RIxZP
AiEY0nnpiQUbVIv2bhdLTWSYdbdivUJuAt0CpnaixLrxBzwk8z+EVeC8X3lcqFlC
B3GsVX4jOKuN3i/OWD88bcnCvV7gPHh/r+u1Yu18dkTu+6CdyT70Q+CRhWl21yEA
5JjsLcuVEif4GEwrFOJku5JY3x249t/vZuIIkuCiDl+piryeb2vePRca87JDzd9t
sGVhxB6wABepQOkfJLqwGdW/C9xYW0LzlrQB8q+v0Par/mPecUCT4d+GXb+h9Bes
goJcCoaoSvxXZ4Wdy9fV8zvFDhP5ctCzzJFp572egY28XzsSshZNUuvyGeiHr9Vn
Cqs3vyi5F12l/V/5CtAbCR/h+xuNhfDUWvT5lNQsSAkZe/uvQbh7UvjDQG6/ESkc
13emUJtk/1r7OqkC+lIdMiwhuqWGZSzhZ0BCUvpfFAlySsdHVIB3UrUW6ZBePtUM
sgGoP4gCBF4tadknh8hxTnaKjJPAbOn1cMWA0d0NJqsVWtN5QgMcGFzq8OqCZDwD
WZhENFHcIPsbrh46CqHN9IBJb6HA3O2Ca1boaK7EhGZiPDWy/SRBYTgL1aVG4m7U
lJOC4Fadi7wM1AJiKElLIlZfgvl7EmdPETQtFVn8+qxQRJ03D3Zs3eFvXH37a69H
I1vvqivpFpxzTFDTaVwAO6x1IvB6N386En81mBFqfCpvBADdOd7XzP9e0Ejtif9o
2HzUoS6NO8WWNq/+V6K3vvRwlr4LC0Djz09lKfp8yQlvRscPqcEMVJGtV9bSq/4Z
vKEybnnwpwqxYpirFCt8sr+WAq4N+daagLm2f2x7LI0KF/i0NMMIHWooIrUHOlZF
p09qYVZ5uNVBmRUUWg/iSNzyL4C2GmKY5kIQmKgvWXti+ix5cmLQV8CfUHGhqopk
3//hssWFV8w6uaCO43dvATObXDYnljUzDF7KmiYWq5v0IbpWxfKafQdW0p8AX1WP
gDktgW3eUQtbDAy6458siFlNZijDDRKchOOSG/U1UJjaeamMB5IFaLM6aHrqPixV
5FBv+IG/4N22536CswuaEfoqlInDu/oMOOWzlFYni5LyeZhMSB6PYsXikpyJtq9H
OItqTKz8x8S5M2xKBi7+ajQRKuVkTZ3w08cvC1Hc1FvHlEqCZpB3RaSPQsXNOXpZ
6vTRS2zxOvwCEYTekmNh2TNBizdmSxjI7GS7DIRQDTdqYqF3gSY8JJjl/wTvkeUy
2tAvWIqJZqv6HnaggdiymE/edlrejSqE3p4Zzc+ptTrpWvuQ/jj6JN73l8nB7bL5
BRq4jCFL5jyaH8mT1XyIhegBtVydlGCKHKIxwk/lHaUPMfENPILmEWbtuzDSyMtM
O8/3JYa7H36jVmedoHfJM4W6lXaKr53vxFYRWKHlhj6RJ7p7gsWesjujHRSPjqqB
HBMHdiXJiJq0d+OWsa38tByhVE9fHGiC2piwB+dm1jfbs6yDOvd5ZieveS5tNOuM
i9GSe1HY9BHnANmrYhgM7hmjT+X+3tbqJXU8msel3494BYdp4PLkgXUO4z6/rgEC
f57X8FQDgq4ggkAl9liOLIeo3sQJWBX/WXcJmewFrycUPr9SGI7entzrltTuK877
J9QBsKxBOLFFKCWgn2LfFxjeNfG32aRXipT4+X9y6xv/4zF+ybyv0KbE7H46Ue8t
4Jm8AgjLEvmnDfE0lMhjZfzeEOX7WQ+gI688f+tigHS7d9ttpcnG5kIjN3HAcxBw
`protect end_protected