`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlHdTNIbr5UHhlS8d66b7l8q9RUxdeonS40kTvzp5LijL
2GnDrdD3Gi3cMELmoF85KQ0l4IG1UJUC1Ilt8TLdUVohY01H+LW20mJfMgUwcevG
7txSV554zO/0gq6Wfju7MN94YQEqVlAsd/qM++SH4FQGD/Q4qSnAspYkvKJfzZKn
iRbL7e4NnEcWr0Nh69z0ZJKdOmw7zerGDNn9nwM98iZmkkCwy/PrdPpnfDvYfnWP
soy7jDCQtnXNH8lT+MPoZqHz4iciOU372BYN+p7tQ4iz40MLwmc0hfWPM1pRDpd/
6tco9FKUiCQRDB86Mq1rrS1ToZCZPhr6+4T2y3BPO05i/d7YC48USchuGePgRg1I
We067qKZFIpeavEOpvPfhFyni5GrU4MG23iZ7qATwmtTh5TWN/BPSLVJaWzS/UaO
uVvUlc/+0xwcdbmskeLd6mC9Bc4axmQCEvy8ovIx00Rr9m7nz2fxCgsSfZ3mlXyH
xKvEECX7iaiYO7eo8pJ3BZFKRjvAFJPyorBlv/r9G3cf3Q0993L6xLHsQ05kV04G
6p4f5dxyOTzKkgZvK80/5bcm7lMJmRZJb8weojLTwYQQYZ68e1RoVtHOPO6JnFZ3
CnPW/Gp/nN3BBuoSSshLD7yC2jUfxH8gMf5mf0afoeEP3+N0gP3fVqcrV0ILII5A
g8GD8WZbisGEvTnJsQwL4uZTIwdD8XIQRW8/h2RcW7paFhiOeEhOPMBJ89grvFfP
KnTJV2CFefo0zYyweMrqRbQmQOVtCOL8owe0wu/WOH7X0c8VVEXkAi5YifdmGhjs
Mj84ji3s+daQs7kLU4qV/X08pCabF0GRRHSEwCuhSQJH5TCeJK6dvIl6X8qobpff
ZBk5WVOCdAw5Th4UQuxoaEVFxBDWt0dZdkYiJbKesaFCaXlAWtXccziuhsgkppQq
YAH9SzcmHTnBFbfMDL09ufSPTgeZuWPbzA0ZNGgXeq/FS++kqZSilwPKm2lv74kW
gbRTL0NxoLb3yyHxlZT8DVppaHP//hj/F/KXIwwWyRfwXH9Fa27NA9q0Bs7wYk7d
uCqGYBBgeDixqxpaFJDI3AheHtnHOVOeVBK9Zw7/NkjbA66xXhuyBIItG3/oXfFI
sG0ONGjLeYStygTTsbFyrxUYOlYD3pIg4e6w2dnPSAv4W+pvhs4cw1hfzbS9kTWG
8i3DUhjEPMTVaMHEhTYBeEllRZhyPCI72JRDUwOzyc+5KqW86Ur1bvc639G0OCxG
p0zMWiXGmO50zbFKE4/P4HA0TE8J/DiS893hj0iYJOBHH24cZYRfJ2AKPjTN9dsJ
ZDSwgsVwv/dWxjibORnXRAI9aWiE13VcwwjyuCd3C1CMjzq820j8Qx1igCGHxQpL
hNOyRflk+2ImDkA3IZ2UGzqljSpgEdM1jwAyKkNy8Y9akw5+lgUWU00PhcK6O0qs
ZaLGIX45GTzeC3PfGJVW7oZZ4h7tTuCXe5IKjINggufcu6KXqjIwoRNx1e0MfP1H
8sFyfUZfRZ8Fz0quTkkLohQEnvm01yH1OSksSk9dXvDi02d/HKEOId5MF13LXiZg
xDT8l7j76cdUSdi6LMbbfeeVdLb1XKRtQFnJxbLs0/MAjzYrst0PdjBaGvvf/OeJ
IIBR9g47juJIXINgG5zHpT971nPeBcsSNtBFJ4OzAWW1fmF87rpqJ1aFhUf1gFm9
2QGivNCAvcz8YRwmnsKbRCb5kXbp+Yi4KIWnGHDjYQpyIBMgFNxkGH8XZAx3aqdc
WaiL+GzUyZ3IIT7XBKS0AYNSXAhypobcgVfAatutb9MSn64KCG3uHXcn2PMrE+Tf
nSmIwD994xy5oKwkC2TLvPKpu9PY5tU35cYY6+8eb+DYP9SjNA3UGyGCsbc4e3z6
Op0Hhz491uKXaX8fUyiOfcqUB89ok+wJ7zEQc5cVVCcvFIZrxMeoIo+DDfAm2OTI
VrjT34YFJ+mDoQ8HqgeoeF2j6MXFeJYS0HgmUXbhuXazYk/5u5Wy1rm3SUU4VGmi
8HMBCOtDMbQD60yRPH4DM4c5mccguXz8kL4Yn918OKc1M3++7ar4w2mqLhQu/953
5iPCPyXvWkEg4hoHgt/U0lkmtWEDWdfAorFB7OI8a6KLcZsAd1qPR+2yluSEsG/u
oqGKoKb8VMgFZIhe+S1Fmsw7ktj0fiT5AbYL6M+V1WxpDujJ/7cl6Nm5bWRZ1X16
/6HIztB2Yr6OWiBgCQwIrmrchaXEoXc2oCK7JzPFvJR5HRKh2jzoDxYiD3ZE9/BW
sS2LA5vxiepv7H9a2AA76I+C8SQJPa2FZayR9iq30CvL+KCq5LsLCn5Yx+1AmM/q
yezEPDzs9cVphRPt/ILSMrW9ACtpvFIlWWIEmuWCbVy3ru06HXngGPrIwa9kLQC5
WQz2k6X0GTPMSFtxXNAy7JWonk1ofMzcl6I43fonTEFCZAwfiT7C8ncIhXB4zaxl
QpwoLTVj3GaB4Nwvvt0NXAdNj1eVPCjESgEYLZ1ctYBJbL2lUYl25zzl6Jtmb1Pb
wvo7JovcCqPyvCgCav2tetdj7muQ654sLmnAKiWs8Ls1tSCgBQJquvx7vHMZdpFk
kj2J2PBzk/66t05y914Z8FFpz3O3XK8HLooFgC54aNe1COAqovBiZ2nkWNJEWaqE
ghqaoyW8lUVj+fDxIH33uoU3La2xFBtUVkXE6cyWOo326nDEXKb00Nh11iOpDlNq
5jZrH3sK32kzqajgtUVl2AXrvO1vCB+/Ett8X0rwdzr0HOywoV3r+ZHuvhEastLH
ZGdbBuYxg4eK04pnbU+Js+Mh51553Nj0S7koSz98tiaYhjLLtgo/VxPcXWaay3r+
ifi3PqJfvibxz7eHudgyInc0Q6vUWbCsAKf1g/B1q6aHmlbj+iywvG3wnNr70I68
lY6dS8Rc87DaYUqWkg5/wAFc8dJv24lFbIu23B/IFQ8Z/4eqo6Z9T4bOii1S2d8c
KrYjmlVd6h5FoovWc41RvOwxK9tzwejCyhu1w69w8BSyWA2l7ahz8RjMSf6/IF7E
nPY2NKEq34bx76q7i+7f2lqNNlGpCndaGk+UQCUs2T10im0Z2alA5xG5yJgklYGx
+V6rn9iUSgiRfnkPUcFd4HfsfGJ/l/iCUVzGgbjBp3P4/8VnbopsKLqFg7eLOCvl
3FUKJT81ERQvYzylZNKm39pC5aUign/X5ZNBMf/d6tj0lIrnZlXs5eQxvdwYnRij
L9yESk8MbhykubrEi0RtS2F9CJG7irUYnGE+kyKQKkajqlDhS5N0/zZ7HkI6jL0W
Hri1qT7b3dAghZhOkiybUchtA6YwJXzAQJJ7AGclQEp439I4tIT4ArSxlVC86I46
rorIKlCzDyFVH4ksBylrnfhiVv6xsdXJ8AQKgWb3GlKcLsqu/PWIOqn9MgrnIONN
2otVZlqhIwboOp1d/fXNu1av4HplHFjKpZi154dHlyKmvFGgGtltatN2xI3zN+Gb
HnhmPBsEY/Lh0lPskAT4Ls/mhrtY9t8DQQOE5LjnOwaMVHSRgZh3Yv8z3S0ApdbJ
rdW3JQfJTQm9gAe/7NGLjVbYO17fgMQ+2iAehgTTXkSXieqC6kzQzDmRy0Q872ZN
6Qf/Qd62VtbG011FPrQjGoSEuO9G6cyWTGzdRHDXZncvUA1dvFC7WA7AC4thqJRV
wS2DsLFkd1EOqZfG1EVWD9J6cnRTUvQ58Uz704sYQnphr4+0Q0mPvXmaEiqtEkR1
jaqTWzx6Ws9g6C45LV80jNuNDteqFnteq897mxYHaiKHbxeGKlQsEtIGEiCLdHpN
DW9TchTmcOIxJnFPn05wispHQNdCyHSZq1bHal9bSgiQyGD1/4nM0S/qTLukF3ld
W6gGUT9VOu5eD+hKebeC1xA/6TmV4kbIRRfaOsAogMk6GPFQNBJYn1YVv+ViQzt3
x3dJ5A0huwUA84JmI2VdXh6UxWHsj5zDQKiWD6LvCsW1IIGjrXD0kjvV6i1+SWK1
BK5OffI5o34MzkM41FG1XTt0Z+bWB9D0JHC2kDrS8NpfpgU9PYwf9o4MkrDswe9U
jBo4zoPDDiaghijYHkSoY/M3fRGJV9BY1OCR9g0uKUCMYwZ2g10+G84V3tCOzmjL
Ku9o4MfZz1fdP+3PIqEiFqcfwIeXp9jzpzr+yYC2jwUbIUNM6B/7IcchiLYstQ3J
cASyYpA6gGfGCTyRoriqhVXFtcgu7uyjZfnKrPW/ANJZz4SehndX2pEHlaI7ZGmE
iiLKYK5VUVqass6sMiZOBnXDgqB2bZJHkv/6RKHOIjmXl//UbHOfgg2eTAjC8EKB
CHwYBxXez+fvazcws13XPFu6YZ/8/eI5pprlxEivOBRW05CGAcp7T/pJM7bdgswe
gWX2mvhrEOpgjtswYNhKvAwJrzIMWnz7r7Tfgsd1W6mtxSbva1MkkzhvElIS6Ks+
IZ0Dwsn63hEbgWJfDJzVrpKgQXBdmVfUQ5uyi2qP0Siqpd+x5mPiBhu6sl9cOEKa
FJ995+Dul2Ngk4ULw8wRpRDFisvTM+/STQCc9cKNqdyUCJ/HLIb5MRw+cgUU2/OE
f+OsrJ2Sc7FmiJEaNo0V44Q0Ne3Zw72Wa9Of5sko5jrSJe9cTU/MrcpgM2lEjy3Q
zRldzPKwRrBKF7CJjEQAV+G6HFok1RYWAFQZRc1LtAW4NTG9LokQAQCYR5yW4pl2
YwNxgLnd6xDETvjVBTkZ6baAbcOs0hBqKTGSNSIOIOg3kPICH4nxBWAgQ9P2Z+By
+pA9lh/djWvGNYLNtGDcMyQcMSXRgDq6YyGyfNtmwW70OVb9DEygcEH7nd8N5h+6
dNaPFY0tlCwVDDKAqP5oxDSn/tJwoU0VGeKq7e0rJTVnvEWdMgbR1sPQ1BakURjD
AMx/l2QJXWjR17KxSss3PIqalfyHRqBTG54QpyZ6FX3dIc5B9W4TOXuJFkXFvZfX
mgG3YhGvUuwxAhwHWQq8ynMBcr/Boy7SF9aiKL5UyiXKOBO231dFRzVAorilf7/U
OMuLvGazqq9ESwIBIrKU7On33gW8c1OjOnvWve8ju+vIEZCenChPsIbaO+ZyaqGu
jZBfFrJP416/DCfdODrZ6jId4icYIQO7AVLisBqn3VNqUr4LR/4o0D1Ehi84v6y0
hPp+JNupMjeD1z5DMxMkiCHAnT0JeoNNGbGX8znN7VACjMGZK87wZV0if0HyUYTN
sM/ynmx/kG/gzLqsk8DFe9XpVJVdSazSor6WxoIJJSrMC+0mqXb1xeb7BLyuwCeg
1eFaeA4fw7PmqMyD0VHNDTkJEw9SlmAof9rj7yy76aBLWP/dKc9Hu9LXuMz1CU8i
keZiZ3dwcNwS9Osz0RL55zcdJUhA2nJaDNemiPecB52YJQM4LOxp162sMcS4cE+N
bjEvVvseDbxHzKZ17258pODBOhQwdRGLhomsxRzxqTNIjXgygXUb4sC2AkkHNc3l
8yk1zK/Qrq20rwSBC8rLKeAReQT0hWzVTluikxfHGJ2YmxCUGqWRWXG8ZIfcw3t1
y8p+4uLhOS66TNDPH9kSNq7FA2kL++jHoLxzxKPMgqLhW7MjxfEk0Wk0hhJmI6x1
XryItEVqyAMAo/aReFRqa74OdfQ+Pyr4k5E/nipeB6qxLHP/w6k31qNO88bkdjVR
3hrBXmbHr+HejJZR/JSIezD/Oha8Wpfm8BQ+gu7mJbTIstF7vsjyc7SNzu2aaFXf
WKAMEH4xUX5o2nxDfDGZ71A1rPJqhftXQ833sMdemRUNNNBaV/wGRH+Fh/7hw7g7
HxKVZv2UEzqvDPG6TyNSYYfwTYnczErO+I1laFNJUTb08Ez2x7k6Q1b355u5RUzo
SE2xDFKeOv1dLD/pOX+zS6MmEJkT0JZXfEl9asMPLyH6/mw7NrS5sJI6yYGiimmR
zzwd63u+piNDTmuUqHpvcmKMe46aBGqcVdZqqnT4+AvZnVghlmCU/ZlUvL7+6GEb
7bEHx39ynCosfxjx7j6p7c2ApIMEDkvTXcayh+fQSbHZYogz+bJktkgpUe0jleBY
omISbDqAim6tOT+seX9xUi9INkzUblAmPbbvNY0gZuT7bJwXIQp6iLBBUcZ7HB6b
cTDOmsigalwSZzbpZOe6dU1cgpGTzj457CamuBrI7kI6+7vo2hLjsBxxHi26BJRs
E9BjuqWF/PFYqaWjwP5jv9m6C320XYxtgJKDx+TnOWNdvVvB0Igbx4a9re0Zv4iI
yu2Cqlr3/FGhuOikpJmdOCYonf5TfcszixReGpFL+7CtuU+5si3U0TSm7/vNJjiV
CiIFH7gnfPVPt4jLyf6Cvz97o0rof3q05zgs5uS9+5NduCA3ebA739FaxRlcY9VF
5fksJynzcv5UG0FsskhOJdTft2ahM0lcwXPTbe5Zo/L1gVXM8zxtxC2LcKSZACGQ
qMK36M/9/xCM2Dlqmq3xQF3mOSEZrXokEaqXa6lvLHdrfuMJAh7Ef4WKzEXOmlX3
NLk+NEwO+pYc1cajRcIxH0FF7IXvDwJUuJCSbpVQMSA6OnmNYQMsTEK4ZUN9cKJz
UvySjH5Gw2JEmnI/XyzBNi5h7NPjdu15c0ZpPJXZE65NghJzcTkIFFCE42WHzbNe
ZYPa76yr+V856F29HDdSuyA9uYNPU9KAXYhCFwez2b48ztJ6fd4vKosyG+rp1rLg
uOCzkZC1X5FXRnEkZ0UkUiJfqkUqbYaSWEb41UzmD7jcolMIO7RmTUuQiKoEzsyJ
Z5ReFNkWsRzF/WhQX2T7nLZI4owNi+q+m8uJ5HPyDJNgKh5DsY7CafW2RKetgUH1
NSi4oGL58QC4kddTZHfrgeAcXpZAG0nLRXr6bu6qg5ARoHsTFlklYxzs4BZTnqq9
8dg8c3C0E7fMT5Tcx8+hxJcZ5I/JDgiu3x2Y7LMyB568Q+L6AINw3U69DR0p2UbP
lBJpoVu2xYnsx6jTs3VFufS2TF7WFWk5f+StL3kp7TcBQvIZX2EQdU2uqcJT/vJU
SiSz8vR44m1A+Sef2OH1qyPiJLlH8AajLu1qK9CZ+InT6Boyxcmj7QIJUO+w1cVE
M2o1OgBxrNPrqZniwB5Ki/iQQl/EVJnLR+/KZX5NdtV14WFZYNa2qXn7VIOUl2O8
SChMjPf0EDSzdAINjMcX4PzAsuf0HisplRvRSYPfbJ4vN7v8DGvgblM0BKI/L2P2
a8eN/GWT+9ZE8X5PUekh+QGmtkvB3hXttRjwn1s8O2Ueu763hJvE5LNEPU8V3tgl
MZ/S8Z/Gm8PJeVwi/c/ZIJaISmPoOapQmyFErM9KyM2DttUFkVALwGm1awvvx4Tp
v4taE7z3CHXTo1hnBf6j/4TDv4qGJhZcUv8iipgMvDJ2wL8X0dK8/ULNQtgPEYYo
qHriGCXAJjf57uWrsqQhiwRBNI+dTbZEP/UpGiDE8635wqBvQrbRKIztAFWOtlWx
AJ50U8fGh0DDczdQ11Anp49FKd1y+pMQzhSZpEJfEIrX6Jc7eCuDxTTta97KP1+y
wULifVe8vSyX/CDn/ftpkK/HR108AHuMUnqZyXV2gWn0BCS7PcJ7UMhZoPRPk18A
5yMZNySovINmHRQD95WcQJJKipEwY2DpM3QJP0kqvy/wZWEpC0edFAa7YL6u6j28
4ZJM77UAYfc+fsR7w9lJS9a+WOEyTJCsJFopCfkTQeslWJWeDlxLEZeIV2dRpK/z
9fdmZi0sZASszuwBrVupln/9fCj7ATq9h1zmvwP/mYCEw+UM/soCkLvuBXcaF7ZI
p5wRMYf2q9L+84afkhQnpTMZrywzGhifIM5SoL8TWaLl+075drnxYKqrEzDepavq
/vEn2roJ37ndOKXi3WmzzX/ycj9RIi8kwU+s7jPi2W28XAOrMyDkbVk9YR3T3OqA
6zCOPBikGjt9pEXkh4XLQmNvmjdteYT6Filj8+lZAgoKZJrOKYRSrpH9A/11uSBp
XMbzz5MBcONAoMzUcvfQA5k9swnsYQbLyfLLFR7yP7I7M0sC++GmC/97kJzLAXF9
j9ECzn9uUpgNc4XcC2W4DTvqztEGhvYfwMIinS2rDb95ULN9PHM2fdqCjKFc7F1d
qJ8GgC/Upo0kBc5BTGG66IOreamL7DJVG72CgLVgDwt6Vdhsv2ZxHD8KOkVGdB/a
Wiw6DeUWTpzsFPwOTGi1MMe61DuwLucLfWG9gAVqcTUXH+TmBWtTWxyvgPh4LzLm
72xsiC45yTRi7LOX9LjJKPgmpJWwCfv5g5gIP0oFl1Rym0OpyeSnGq7tpdE+dNLM
7KfAbXcCaeVptulZpj/gOgHFvbTIHJByy8iWL+SP2oCab4Bag9/dnD+li9OqanLO
nVDC/dCJYSKYtnVXFJu+IdJtMhGx2tlrgci8qC7BtqWFY6iWI0NSa3Z6zTWi3yYS
AIhLhRDgUCakUz4obQikjzD5TPJc4YPbsmKq6KlFEgU/kA3YTeIsmPAm9/y/k9hI
9x1ICM9aEGDgFmPoPHi7gY8QQVYewyZ3b7ux4h9leOATeZMeykBWFQgLnHC3NhfS
aarNWLdozVEeRyRaBGRQPxhlyGHS0E/hBpkk6KTyU10yO1JCrKnlbOBryePK1fzy
hJiSCqY7IA/IGanUT+Ik0nZ11WaUqH/TYcAUt5MLkAppofkoDuPXxgzfGITI+nkT
lKywrhHGijfz+mtDQLTivezX7u/ysNs6+6DvKXT54wtEJgi10oDeVKJgqJGZyQo3
Jlkng1ZwO+m92gsHs/Y6CGGIWdExBY+Pol/kRUafm5gdNHEwXjogZbNUdKsMAZSt
SG9txMyULrjUgghp7iW++Wkilm+Jje27Jcx8WA+uX+pj4ZmA0ybl/mJlSOHU8+Kt
Ff8cBQSQAvEGzUq14FBmhy8SB8YBsX3ErLTwjc6YIn4qrSRfhEKxFfEZjwNTeQk5
i0kLChv+heiUTKj4iCwEGHpMuNkqSk8qDUSA6D6XqSrMobVWthSTYo13s6Mu5Zgb
fv1Uv3e0jr2pmXz8GMzP59Pa2sYOlqeB1WN9arvWQx6w+Wzpbm6LIGFgKbWWM1WO
Z1HCy/PPf3PKKRJLUoiVQbsikSM+5978nHs16DsXLlTVDuKbVq2C3YHa6QjmnPXe
Zo0ncXMn8LanBzRT+LErBBhZ86vvaVvozLrIEtdSlDqOpl+6xiz4Itl7nqTSllJb
bJ2ndbBpgw6jmtF3wfYQxLA/sCqPJ+FTIRMOPMizeezZ6iuAQtICtIv9CivcbJBi
B9bPkvekorwwq50sRkzWOrlDohmQuZcnK5yBHvHFhvZxGbrs7n0gYKZN2lmy/d/T
hKjK47GMLRqWl1IcMd+Sir186LR/8PKb3Agin8Q9t13E2JZAqDLUdEWw9VbcYHHm
HvPc1kyeLNnV97ort4lwCrk+qmRTIJABylqG7GVYLWq8hy5GP+e3tc8E4LdOaC4G
TvnDzR2L/8OozVRBGKQmcYPs68YqTo/vCfAHeW4+wjBJP4VXYFsnGdA4sFBp2CWV
pRjZNLCczxRDJxhxGvi7G0hDKCUSezrROx9J+gIj6uxoL3GfvjO20WT5fbCdeQ+c
mquV0+7SQacTqglgsykF1yRFtO0f/uu+kjMU7yCfH/I1R6AfVaUU0/d+aiHhjOdF
4QpkrSelm48UdRWHomHs9+RKnrPkle1UYOmuJzlB/ffb5mHjbfxJ/9lEcvtFqxgm
9szrG/P96MSNT7hTqbY4j+WsUXalisOjUhq5MCbRQnwVx7EMRrHIyFcEQX0bazzM
rh9XngXIPkJuLaIMzAg/D8roF+BCyHYdyvtEUVgomXQMiuUSsHqr3I6WNMaVm391
BfzGWbFu22+uQPrV7OLw68O7Mpn+usK3BPy507SN6Fv0lvYJKqEt2dd1i5tTAXLL
fmuU/mQpkCpBwHvbP1Lpr/wAz4UBYHK4XynCtaMfHijVQ1lY5PrzqLMolOO5TNt9
kVV0NRr0mRkoMThGj096dW26amB+yixkzRHlpEhC6ggGyI8+DKIRFNUfNDwwQB+E
sGgucw7Nd0O/CRvmHGPUb88DavQ8saxHIXWeqZw8t1Esde8N7wW+ww6axP73aOUY
hK3NoU2EBgP9hJlZFdT7SCJwPIlwRqExm2AIR9Nrskw5FG2IZM7rCNAh/SO60MZU
py1rzmw4G0FAZHo4ejIwjDW1Le16TAOWLXAT+K1fuAJMoVxLEwXpudwG7zeqV/PX
85RoUxiWhqb4aShIPK1xDBPW9CCJgH0x67FaYXxf95c9irLffqULOVOVDsU+4fpd
McB3tOQlbXx18Vnqg1E9dU1ZXv42pW1BzBFBA1cv/6NBfXyLuff9Yt6mviU56oJ2
ZcjPIiaFt4NqqJurOVCK+45uwlVrf6rRRSJmd5XD90v7ya60Kijh1VDOYIOJXRnF
e1XaifDUPjCLj/VrBO7JtDZ1CpzhxCgKLmuVZDetLlxOdkW0aDhmWEsxwrHce7za
PLIcffgu1Q+qlhkzGIHkwDVsMovdLV5WZvXSyh6302QVgwa3Zws6Ij8jMiOyaFqO
f2WMk6lIyLr6M6+brqJLtU7ndZRr6xZFzdFKvUkerm7yWJuPPS9DjDmZn9WOLLsO
VYfLgS2I6uOU+HMDzdPjGLBBZb2MTAr1GGEfKmbsdKiCQX6Fbbi7dsMOyWL9Jp8W
s0BpKbDbi49hv2dDs7lF//Dd90RX59Yn790gGGfmgdCmOO9ivaTeWDGaEdtdk5sW
fSjdsGrhbrcpfseZalM2aCfSghtJP14J1xCcA1GSpS8Ci6tiCJ6tUU5Dprd2GtBk
R+qQfiy3U8fn5hhrIIYjBQqc5SX0+G77+qXNMNmU9oCLbjdy6P32095g8xkXyP5H
T50l6EeoUtnJeEInrBgWIIhCHr2s9GnAn/FexBy8I3e7eYHM4+JwflJOOo3HFInE
YiMML1K4sans8+8UcohINsMV6GLDGhkf9w6JLNEUDkKojWzCPqrKNgTlXA7MKrPn
XfF5f1/0j/rTxDoIh1ly4GCqOhm4OnpKUKCQj6Ukl8Y/8tRojhmHjuG9SnKvq0HY
X4o/+Zf3/Hc+ytP1qZUKQ/z5pv9j0YE0Qeo2sMFpUlWEJJQlaTw8R3ohKJbJjpjw
rv8UiI9P8e5ToGAN+j9PfN7ohHTaVyK4Cnv2idlUBZkB8RkrOMfvcNIfXnuqhyY8
ZW/mFxdrVbXhf6quuODyDQvHQz0uPDZay1KRi2I2JrfgsxsyQ+hiWFO+qayXflP7
XV05U06p/HxpxdgkMJrOS+VO3i5HEhGFkDJvXi7SFsgVTb4FSk8AzIC1DLEnnbth
TLY4gHi3auxV8B9/4+UB/szb4pKEjmgFGvcDByZUfoJ/jH53lno7qYawfqtXkOVF
tOgHDbAClx8jizCmbj44yevhT5EhkqUE9LEiFihOf2rss8mJXztjunOeF9EODGLo
Yf3MJUCpQ/W+Ohw/V4WuUCpVwEb7Qv0snoUJOy7xOG4H8KrqFv0HCT0kql+B6Aff
G0k5fJLjtiGckGsH5kZiAruE3LoAV/Q5LFtDUfo+GxKZrb7JcqhjlavvD15L8gzC
jHW4Ja5CzWxeRA0HQXFP9okxADD4RbTpXHjLDoMIFI7uhQbG7AG4oq68JEQ8Ylqb
7DzslSts9ZLO6igkUCqMltajLLcBf4mTMmZb3Q1QK5dMK+/aWwR6tO+P0TTWoX4X
14kwsY+iCPIt0Rs3Td6mz1kYxa4FEEnBaqR/iOg0B+eu+7zpVRW6naBsh8Sr6Av+
TH/Edh58MeRF/gVWhSNBPHI/cfm9QuishtwrjVN98tg4gEgW2glzea1vKizC28tm
mAuuQWBnOTcfn70llQo9jvYx8RZAMqWeKqGSxjQOiDh76zNYp0Qsw/hf7oVEZjzo
L9l1ruq9eXLX+KJ7h85pryPgPAB9QFLViE33u8Vo9F0DSh3Ug+Mqyqxp9VMsWsMj
TWIe1hEdOPR8fmFc+luM1sy/1+S9+PSrqnnSxSF6G1wVXhaXl5MlPYdia0acBDew
GJvUM5KJS7hd6YuTHAzZhGb74nbij8UGkTQ/g1RUK/s70qF7ZL59XXmrkFcrRLja
rctwbBehba+FL6AHYAVEgeWxzHE67X7SLwdPehGcQx150GsHDkiRQiNNzrX/9L8G
bvgaSuSxsc6SqxTXNb1Zrxtsc+XR6aEoa44TP1htbcScL3coN4P4aN7Ks3KphJE/
qr5WOiOdjAYZLspw/Hi4UvIwu3iT8zNx1sfb2Lzl6WDAdVUJ7eaZ+auiEoHXyorA
VReIZkt1PLyKgUm27fhSD99cSclTPepEfLHDpDa04aOFYXBqtPdjGFtZ5Ym2yWNl
ai1EW0DJbw7Nroo6HxO4+YWn/r1AqAqatOYdyIqfc99i+rf2WwkElxKvYLCqo3y6
BkK6vTkXFwd12D+eg+YyeMCmeQrx0+gqEEGQ+VKUtnKMpRQsEzarbkSCLmIhDswr
Rrj56SFyCLJevlEBNCO/QN7EM/jBWxUfkH6Bzob5bIKmMm8pyXLVv6prwwRzZni6
67AYGJvRp7wGWRMf4ha7iGAh5U5Ch34122X4D+aUL+P43RP2zH6AA8y+KLozy/1J
1k3gPMN4u6sN8q7YJgjnhHXD7E8lzTXZZG0mVs5CFOzkNL0bGzwTpXsqC3TkqbL0
/ZQngdkwg80CZ3+pC0T4ohZ+GfXjVqX6VGsji5VeVyarXh+p1KR3qt/zTNXBnjNp
hxbzVaAQ0j8gBoRvqQe14lm+fIHwWG7cnpwDmbRjqEWlM3KGnHHzZ5ymr/2pF2Sc
IXzyfTLO9UBdttDvkuinj9Hppoor4g6Z0gD61YE4ssHSgjBpnXsB/h9UeoZAWMUv
oaHZb4CS0xqLHBXjItYZzZOSEsHJ6yX4/Z77clP8RdkOBPw5DQeLcDTBEJlYXpS9
yceu7P8bFyKAws2MxqDQgWw13kvYgVRWmjBWYxITj7pkBKrwwqJOm1NQ59d8LCoY
sLUMcFCy1KQvrcnog3pqzh/sDsSnh3Wdta4s2wbDK5y6zjm20PC3u9lsuO2Z6s7A
aIZtqgGwxPLVLO4eo//gt60THcVwu7fzu+aDvviy74s5gKsUq+6MWWDhwBKMlur6
ELeqpBdUgbH2+lrFxdq2mlDlPSW86SN3g5o+UGtG9DIFTNBoUKUxW9HjVclj6aYO
mcAFJe0YzFbTbsx8Mni9VOQkSGm71xN9t5KXNmbs7VMGWE71aYdNJwOHkNvpIkg3
Jrd+iUmyO0lnabI2FtTkSEUTiqm/dc/VZJnJgIgRMtu0gkwneg6MoqQY/y7EuqZO
e9RxXU5UwrwvVAqk//ZGFf2yaSRph8g9kH+mXt2SOhQ/291PwdcJXz23bJprW/1S
vLN+4YRskXNGxSlkMw349r6NkHMVRHidxLi3cwfGtkN7ORBzV3NtSUQ1BRuFMrRp
IWgvkHjhFg8szFLjGw03xgVIMtdxorAmANzPpnYAlzt7SH2ryFOFZgLLu00Pu4uM
WF1dgpfBuWAvcfEjzOrOKUUNaRHEOUtyAqFBiWv2gOcREKuPzk12lKfA+BXSQWRF
L3U8UDA1TNLW5nNRLITftIOxgBzFfEgrfJXnsSLMGzDMX6nbqZn6OvCC8r4ammeF
9jOnprMvMurr2/UGmuwnqUZaoIhUUgfWEyMFsWL5w/qvqUOpOCg3lqP6EgLPuY08
P+6nzAbK4tb5/5x3maMHXld96E/6SUIsXJSOTq0YgKiowBT5Gkva1o/2okumIwz0
viI9sm62rqrXkaDTVLRD+fFu5YWQS6W9Ald2R6PYy+gzLuOT+7Wfe62djgZD4M10
nH5EN+ZL6YfKlJKsZ5KrPf43Lfa7uhhpHKWiBNGFDw6WPL+lQ4PmKG11K10lB21C
vAO5ETftJq9TahM2IXWdsGy+/fjDPyOA2GfbMttcm2fW+Fkh1qK1IAd0iGKLqqan
MJUT53814Bj2BrHUOquQHimIDbBynXzVt6jeAtL4FB0H3viXrQajVd1rUCaMvHz6
02+lvXGqjLd5Ns/tOWnKk8GjNgieqyflt219mrKffGCj2Yo+EeqX9JqE+QgFDW/R
ts/osHE47hpXq2ZTNLQIT6Xt6kkRbPQkRbXNNoX1qr6llemS2dKnmJ6Y6DEvBnk7
QoUnsoJeNZJQvlZdpRCQ0q+0ifexXJSDYv1hHsa5b/RLVPi1eCeR/thbOAokNN8K
yHgD2PfKtnFg4kgDV6kZmpWeXn+I0k3Z1G+Q1qt+Gq/TnNg5QQ532VWxczA103OK
LaHAL8t2e20izGbc5LmD6xA7emdjEkX5ETKDEdYO48g6k4qrLoT76EVgxKUD0svq
OApP5dejsM6SJ3alS3erSbWz/6ULG4Md5EqqaS3cBbuAk1H1kOMKWnU6Trl0S176
w/dH9vOllh/V/7u1uRgDpaOtHB4OWamm/6eGZe5eDQO5X+jepm1zzXbArMmZCXxA
rxvoOynyPaSFYC2ng7R5g+lfpd6MqWnIL4OzUpYomcSAFRMPG58qrUQikZWTEi1F
cHwoAQ4tjptMXIIlm4khbgiqdDyuImakYRXLOF3FRcisMBzN6/+rD3vJl95YKKGz
OlvqdrXj0eVgTbOmRcQrnUNHZpg3apoGQdjBLHMTXK39Vqv5YDa6CoI67wjXmbRS
CY0qlK+reh8ZQZ1VK1bLXTpyN5oedzPfWl+wRJfEUqoVLHsnxW5kXmMZjthsgv6d
nXG/B9LIZ7taNpptGHt1b93+iIRy2MZZ673MiNIkXD5/c9pqf+3HpO4dQW5O9KC2
Mhg8v+0WAm/qOt+Dg223wQno1GCgwxbihESYbb+n3LE0md9Ax8RTSJ43J6EzJWER
XIZ7v9U+7JvqWO9ETXwQRONiW5VidtsGbE7BxmCSrhOovlw/puDkKxzcSHB0Lfa9
arE3+AIK83n/ATeraf7N0Sadsjzt/9rQiWRR22QWMpsxMWm9NP4BMgT/3OZorkcm
nE2l5jugxOagKgfQcdabad4e2KIwk4iuUvM/N3C+RF71ST9vPBDBzUfhWT1DheWJ
1G3vWKuLhXSuP+i2jtkwhZ+mTlbjtDTkmJ8DhgjSHGpHtzwLYvr6dJv3aWPd4Lkx
HvRqsSKtSMUZXzyviHH0ukEtmD/sBX8CCkk4aZ/p1Ubar5H3Nr3Ocmghv9KxFzN7
QmGS7XpTwtUjET1ri9xAX12VUSIa2i1WgN2QXSZQJOOPmYMWKSrQ5EMT1lUb0GTE
nsBn4fBCd+oCKiceveSHNwr7wwmFS100cXBMnZwNC+pExLDEkdl8azo2AvLGy/pQ
MBmXk+ntCi9HRakjD7s069BVCs6bzON/c9ZsXnWP4HLWZwiU2x4PRhBkfGJubPjj
OgdbHs8wUuqBP75/Esa5CfIUbDZEcIsywJdbMlM8LXltiiYJP3/WhKQsvyYn3Q71
ZkFnqyYZfhFwjyLRKgoKZ8q+Q1y8Nt2AdigvZeO4PbpsVDffHneEDY9e8jJjDer3
wMBnb6R8yNsIhyPWJM15QIXITtWebDCbdggrCfdxnes0cLNpIzOYs1iXw3vT2yej
zFNzxttpNS6Yd28vN58MU0Lcd2GxD7AdmclAf92TpACPV2m3OKb0DYsQICir5vWt
0fA6NZETTRpUxJA94PUSEutwxU5yAmKprH53M3y9pMA1oPl1AALkmU/PB0IV48SL
1COJeMwkV66YSwoRfyCHkgyX1PTONtf9pU+G7WlE2HxrHkToNFWcVJrRrVzLExjK
ix+sKIDNi02u2BbC080GCXuF8D4iuEEr3VlK1A//JdeiGfBWhOz7nTUSdjcnL1f1
R0fDfbpMV0Nkc1lnkod5FIYDjaC4Fg9iXTOGH9iy1HRKxQ7eZqtz0tgEwNtvzMWh
JwJGMLEKmbZvfaGzX2rrh/fE5BeAyVf//aq9dvrWJ+VyukRyyzSJS31/zdNLQxf+
/dmjNp2/NXML1GxiHOgDfW5kn5ZfV6QReCm1zVZn1TAhBUvrfC7dF4Plm9Fk/Lpo
Ag0dUN+1PMEoDLKQ8QvUBdFQvIldHpFCJl0ZCObHkzQMY5RfYiSFNSlGOqsI1ftF
mNc61NJQ+bkEAifct7h0VlzbQOorENvZheDodONpQte/xaEtjpqeapemVyqWBdH1
BU5v7QlTMww6SCOijsyA9KZoy6Dl0YjZGfFXr4AHgEOUGuuE0GShxEorRdL4n4uo
VKSBC3zjTaCwibZkUeQfvy6X+i1zwZgyIzdN8SOIUxiIbxxhBbyr24sMBU7Bfc9p
yjocAaG/SlzMyJK4LUqavFwXT1NVJPptpo812/mchNnbTC4e36WD4UkXtBrT1ev1
w7M8uJEpbqzBT46fciIzauLPXNIhBRvrL4MiVoRgsDcFJ+AsX5/Co2EeaM/WkTG8
1F3MjCuII506YeBYYNQIlblHgYSqIl2aIRK4Z11r5BljSnjacb/cFFjx/rhkETXm
BTffQcza2TiFPrE+wW2N4nUKf1Nrvc3XqzhSVxmm8pEnwxqga9746N8m4HMIcxek
FKVVNjGHFk0f2GeKElhjEE5Qo66yKBzgVZ+Qde1NrQjenPyNeiVCWIulzQYnVBsT
cuzblW338IiCwjY9CsHDcGwv2z5M0iObyw2l9JkxY+9pFKSXKqGnUNVsy6KBuT2E
rHRng9QmGRdREck8goX72RtagPuxzCWCcUsskOAZJsloUkrnhFQLl9j4WAS6PG+h
aA8SaBPEHp35UohGdXgI2ErKEStRy1ZKnbXcHoqUXUUg2KmqaRXE+2g+cbl/shtp
EiG1c6NpFyeNKkLfUggnjij/cTIjKx8Bm9rXJM4HO25i3twBQtQN+ZJ3ltDRC0o2
go3+AIhqXjQNNJWtdFxHsf5FEwinTVsTAUPbUMbXYDeJAcdvVKkOCkkgjPo8mbJQ
TDC4W7ER9Wbvyd8crgVVHYrO/ngAztp/5plllsiCUdwyaNQFCOWEbODbr6T5f96k
GSpMPqJQoAxfURkTO2VyL1Wd1bQpt+b1HYTmjkThSMDE9gLPlE+S7qv8BJGl3Dhh
/OkxdbXRdWZ2gTfoNx/zBSluoUXfon6TzOrX3B7INlKkLYcCPjuv9XK/CmMKSW0I
/lAMr3e5ou0WbPyEU8DAEY0ARDxNi08psRWIzBCMmBFI6xJBHsvbf5sIoS2T8URO
/+Quc5lzLQwotR3OPEYT90fSnqUwnnehLAs3c9akzI8njlV5rfrluFCrFcJFzA0B
QVZz7wCSgpGWO/Sx5yJ6F63YwVM5lQdw3G6AK/nBq8hGt6s63adG+4UsgVku+OEz
uLG4zAtYn++IeOR6e8VDMctC0PXJFua9Oxeoh0djAMJ3NnpgcfQ+g2hQzETvEFU9
rzraVXzrDNcIoTwrX1dCA/1XgoQiQDJclVdZDeRdEoqwwOGSj6kftf9TGHX1Wj6y
baFISvFBtN77oGdgUdajQHPpi5NdZDF8EnKHdWdq7HTw7cVcr4CrCfqqaCnYWUKj
GWI6jebKoYMzT8nxcG+C1OoKegRhzAqDr1v1GWM6ivT+r47S8cBrXxttW5/UVNc+
VvdEyCe2VH6IvyMCkSgrRzTX9uwlxGEcyaLCINQvGn+wyf+jnau8C5xwCXPCG45L
HzAsmIUPFOnSjpUrM/hg7cPS1ohGHScbuogujmo+Zs3hre2ydGLhkV4otOyYulhr
mYPYdmvAHsq/XKiyf3ZshMAuE3e7qf67UDwKLeUm6nGlhDMi3S2AYl1LBqHjMbOI
pcFgqR8WWYjbGTfDh8whhTXevp9K0wt9eP2OPxLI5Vj/Y3pLXV1hSc+Vuwke7C0d
B2TZ7v2qaniCrVscpeYSculAQ1w9vaO4IPxn4iHTrVIVyTLkCCk2tDR8r1Zk1RBT
3LvxrCn91ufba4CgTKfgm1wNZn8cNCobRNxNdol4wnCYhyxePGqVcfPWPZ+NxZDc
+k1Ht/p+fb+i15xmWqOlbtP7iKH9A3vGUTl32MZvRyt57VhHF4yehLK5f3Dw34eG
CYMJSQZl7OfHyPD26Cr9jbdZQe4ZiMZRP5UE8zPtIdujyV4CkwNcKxojEl5FMTSa
hlEldRJ8/qZuC92fw0Hp/cDV4Iy6t51a2p9apJJ9I654B/+1bnp0oo84juMPNTbE
oHmxaEdStirNbtd2BgzmvRqlrfNufojVyqhsmpnoY4gsWWGHnL+9E/ZilrvWFRpc
Ts/yT5DoLx2LmNtV25Goq6f07gA7xFs7AjQb7XpEtA3I4njInIpuNHQIN0l12vml
FQkjBlRzTWdsQcgaNgp7KzQSbCo2xG/24PgcAK+nzXjNGgtpL/WPJ3KsF96AAdnf
7ZqfEZE/pbtGrvcFLvDrV0st7I21bkgH0tWeksVU40MQ1ntARuuPutk3t5R5nvSy
7d2Mzf4swV6UcwOThTHjykD96BhC/uXvMOf35DdC3GljwJ6ojoKAc39LZOgc+A6l
s8ssT/3f9Mo6AxMhX7TaGJLcUtmoZE+2++JNhfiFUsfiUWISAUXjNnhv/7wrTtuF
iVFnDv1EJQl2Vl6BfdRuJfeSrv/4cseIYZsh3CLtuVOQ4hcvjzrZ8GPd1n0hyQgY
XKEUc2EVZ85FP9bRdb90Enop3f6CVmTZJs8TCQ0GOOuuJxg/NtqPqAG94JRME9uX
gGahWj09cBM+jO1lGnfWtE1TG1ice8bgzJ8gzNsJBpKoeh0u2ApJj0WRmRkQmqIM
bQRPpXBxBW1PMn/ykTHtmqFdPf+mlGNsomfr9y7iU2oPYo4paAzDWPVyTZuDuYBl
e8NC4GRHIeo6VZf5GSdD1HxKEbQFBrUBnrbO09as5uDPq2aEW27qyUuyASG2bAxM
x8g9Aj/xs3ao8bV4hj8PQmk9/YF5CW7FdsTpH9FGe+IX790QRDrtIrWA1OW7s2uU
rMuximJCZ/DrZeHFjvMymhpotQ/QUQnAThujT6CcyYXEk5mdmI7MBGApvuZuUOV5
0mYFVNZqtfkKVo3Z6f5dZUJowVr5XrlD4dLGBLEg+Xwu5nvrmqEcnReZW/fRe8CJ
FAVC4UxLDLHxKttv1cu1dla82jWobOXTVmCFDOB3TJ2WNYiF6FKqD4lw3POO1C2O
QUtFlje7iJpgEHMh9ysNhmc6kiyUJq/hnYOxKwB10uV3s+PEm8IznJ9t+IJ4ihUx
uPyKMvJP70BJBNi/mW77zAvVNAMu0M1jMxpmXdCQcCw/+/UOIH3G0ll+sp3JVsDm
EVY9XNOKbNBaMMnF+hwxOqbpMQYeExvi22UtGoNwNzl2wbjdNh4SlAE8kfL8xrHb
NxXrrba8LPGJq2yvhGxJZHcmdjmtBycvyo3EyCrNL97AHT9ilg6YWBuiMgw5/dWe
FzTgbQV3u8xpyhXg5Odt/koIiPFOZtGvAmE/W7HgAVphwzt/HA2eZmDlMzLdK2xt
HmUpM8Q5DGn5sKeNzWEYNhUOrNYySj2kafjto86kYtxfJXAOter49I5k3Wmq1FjE
/KQ33Uau7+Cul1J5LG1OlR7MZhqRJWmtbdcNf3fZOx3fciDmcyen2qRIDVS+oH5a
QDft3Qd3s7rMfO4kxFhCcIGF4zswZWpBKvybZwI4bAI4Kmnw4K4h/ZJq80Jpd5gU
PSM2p+a9PaYk9RwXf/6tSEMSElxE7uVy1YYz7yYr7pqyYApmzg1DlgPySR9GmI73
/5GcYfIKP7J/AM4wf5U778I6QVCM4Lzk3s3uVbmtYQtU/oAq23LAME6qKcBKJhEx
SWxSsdCzqdNlgj4v04AhRFjO28ATJ2HSs6eGBBOsUFpOHTc1ye4RGIoA7sMYFXTH
mzH3YpIl1LEgnODUohzq3aR9BofEmCSA68eqQNaAOZmhCN7HEQYz5/GH5/an5fon
YKlfVVyxrumuGA65WKx1qqc/Qtc3yjmJ0deuLPm/vCcYyojUWBjDHn6gIRQ65mwM
7SKdPAyazbDX1GrHDH6vr8yqO/sKc+YABWNRl51NAYW8gEuSMCfkjELNEAwTgz76
I5I5h7QWBj6oa6RZbYDsswkG3+l//+gfaYGxm3dl1doTX5FfxddYrKqMY3fswhcg
n4RQKe6HRb2RhcVIG8UBy1qSmoweZPFIwMfaUEj24xcZZk3vco6nqt9+U5qbnh5y
oE6WLhKSKhPx1URIMZ6ZsTsuI8RxTpFkI3D6YA1qrsqICzUrTpeITb9ojBHR7QPa
+VSLomyjOCyXbFInvsZiD8vI+PMfVa425A4gxJ8bQVerqlpI11v8o4BBEl0nEF1k
6Cgcm5cOHMOSSjXu5Vq8tD7RE+WL0OMWZUpk7J0Ip+9SeFeJNWAkXjbR28XCCjLv
yTpzbLqgYNJEldV3NysrnHctauzi2wbsj19zp5MjZijalyJFjhehhmNcXSQlnBn4
3Q2Kjh9hzBtwMg0l8qQiwlpbvH4RGJO2LBuz5S565+IBfm3eZWsX8uNU9BDLRrEe
cWyK9n+87ADG/tVuGEkdfnfXQkbqFdJmRBW/yLuIkZsM3z4q7RXGP8d4xo/DRbjJ
nufppFCA/ibDuVnzkXbBOJwPSyDgQvfXnDFjoTku93Pe6/L/aROZuR2ONZ9efZ72
Oeb/oc1PAVEIeIn/yknRU2e9dzMQvjJ60FEmuKME6QgPM3qm3S+duqHQo8GWFfwL
9KXJyxBcfA1XzpIKHwC3N3rGUtBXsuaj3Hvl4Uw8TNQoiWBR7fQ4B8dshHkXXovX
SU1RF1FtPeGJkO02hXUa4h1OWeea0ZSDaydknjLJzFdc3y3wyJ2/OKBC40R8xv5U
4V1Lzuf1s5TnFIqTwC0qcmDD/VHDnHowkbqXnbxsjkpYHa7E4xr6nba0zAeeHSAO
mNMyZndasip1dN/4e9bRYaffVkPt1pOr9T0CzyUTIjO2X/UNRS7MKKeGcFbWNwer
IjWJUUqxlocICPdCRABd2S5LY3yGn9tGSe1g24peC5a1RQ1dUqr0gd2LaA7aC90r
myhqgVlQTplGUJ9nQBKbaOhGIFWOgsPqblDUtiPXDeIw85niKz4nSzZdl9+4CJh2
AWsWfDZk5gWwun2lOxT4Ou0YiU8yDCfJSE5AZ2CJzE4XlQ7G6N6OYsYFq6r17gTu
Y7zwOePdKn9Gflw7gf6RZPb+B7AamQ+dIbH7iO2RrO7lv55CfdPPMnMArVe+bPwQ
zto8frHGAilAUj8j8+ytj68WuQRCy7pCjhXxkwluMMRfbEE1LlF08BHeNfrcGK+c
BrHPFvu8XUPBAyM03a82gloDI9TaqlJMn7CEocdFVpGOLoHdZFftvI7rIEpQsPf9
zG5uXmb605vurgpxnLBhheCJty+hPXlVFG42Gb9eAC6nIrTLB6gSGf58KbdhXILR
lNP+DQTqo8/2MZD1gHl0ixZRk52HYlUEjh1SU2cRqTS0A3W2rtKiGYgJxwGX+PCW
fb+K809t3gDnQAjZdMI63zP0ORoNQMBWR77/Puv407wefUNa0cXXpmsFQT/46Eya
aAvDaujtvUYP/CyNQ/R512lBFV+iP5aTYZYQGd+SPqwVEPlJpsrIjOZhNuU7/Jwb
HCr/yHw2+8FUas3aN+7Qj2H7MCBFn32UvI+rGzsMh+f0FBVsPwav1QiMBLhgILDg
RClxI0pd3BCKfwci4x0coEBCynFeXdSMPXTbnP/tZpGcQ+/rQ0J2/IfR25IaDd+B
0ATQxzvKTPTp0qETz2jftZPICf9TW+GYb3ZKo3LL00mZj12PhXxq/MJh2exISFJj
gc8BIUhmR7eA6Vx2FkxpV8aSfy/v7owhVoTA7rPGFtXAd5dVyJp4w8j8p6pHyqSc
gLBs/ftlOOZt9wwXYIA/bSv/aJjqy+OAhWwaBy4RVVgTFUmsadhAMSy6MS16PGet
Q8lts+GzO85KdF9v5OnKa+Ev2nQSorMfmz0XZb86ajRl/vsE6f5z62/wGA9HoRF/
qa7yDKZoL/5O+HLe4VG7F8nUu522hNQHxx6IQ78SexKss1kHZjH7FVFJCzExMU4u
NWQ+Wgm9awAVcCXPumvReWAvnvFcNLXX3t/mbrJ+fVttlZ+PM10fK5I+G5peu7Un
9AogEdASQM80re2Vd1R3Q/e8opSmHPoZSuPJPJOcBpF5b1lMJplnZm825J0iaI04
6FVZekC8vClDWeas09gAud2hrv8+OTIlUy3xnjw4/0M5Y3GDkYn0Czavwjff9C8W
hyu0YU6kzjgM8cBC5RR/94qq+W+tlS8h5D5DFfzfT6gkA4Cm2NNBdPBiPzEH5/yy
oHfp5F8lSaeYaLVBGcNV6Kw5kh0y1nyN6CvW0tJNKyPFU+y6HXjJ7V6ec67mCq9n
/S5TaJi68ZQRiD+Y9FRs+Fu3zBNtET/PZfpdJu0KbxsjXYSxSHYKZ7A2v2LJg6oN
4wByQl/py1qPG+G57j9lCyb21e6tpGMeMZyWPvbI0V6wMMf6eeMu3RE5jrTzQFy2
+bDBtByhi70OztdXybuBzG2nsMqgJE74hJEPDxAeJ8azmCWML8zptGFiwrGE4SG/
6rO6va0VIHn4v+1vmAdtZK0D4RylNpqB7efFEzfQqaVa0SncG2xwjb4+uHx2z4Lp
y2yo4JPPnLMH66aq4eQfXV7fnzS6ixJUTx519qr7bcQYiE8WPiZTDIdbT93eYM0A
1rKiEe0iTYOloQ9ZiYyGmoul+790wZyYHzAngtEqs6OOFUjexdAnl190cONdsoDR
tsy9besOzERlvjasD/Ig8iDKEpvGeR3yT84w6Nd+rAW7Y+V632STzRXrauaDyZeU
zuVc/hf/XOqM+29u57b/2FC0IzpomsLcozkSV1YAqWhGS5Q4rwEk5d4ugzyLpSl8
CT3/gpc+AcRSMjzsBMgl/6MM+zAWJzvCk1SY6OK9MHPBk4o9IaOjwSjW/5ys94Uq
qyMdASBS2N4amI00oA0AhuUu3KzxxwiAFr5FgaVCpZCLlbbVZfO/ZXW9WMmrwyAH
tWXwIeiZ30JUOzrjSAsWkLM9k5V38Ffu0yrAjLOSHXOnCAs5rURVtAq3xc0IhExh
3/V/prF/HmkZ0FOPg+dnTXglhNQX0BkSaqY9pdvnpgZW7c7prTWhB0Mxt55BsAmw
vUDYM3qles7Zj2INpkWf2NIkRaQ12rCGGRGVJY75epKT8tr+nOC/+P+dxUPI8aR4
SnAPx+fo9Sy75DdXdWSQ5RWrpBrRaAM1i7WzYPdVel0iPvfgxbN1go3sdqv4G5CV
O+lbPeJNYZyUVQhlmWU2g8b5OglPLenbCrBKG2hXi+oLH95RnjpH2W8CseiYwVsW
Es3l0LCwT8zMFeEQmUIfvzRetvgoEZjbFJL14cfJRhVCaAbCgFq9muMG4VH9L6k4
ECZh3HHRKKoYBjbv6UoHXR4r+giLnZv/Ng60sMTP0I5GKAYTEEqTty3BvCKbgLyU
grQEYQB2+9lKehLzD5KXETdYeJUloL8sVrfiAEDJu9FCO6oPiGDz40009gl/XAU+
QI4taHfZEyKzMIW57ofULEC+N5dlXHst0CghtAVIfRJnaGrf1ebAfHgJfj3a7pYC
WinA2Gt+wfsS42trJa7bL5WNSyJ/r5y+ghpTTMfQDjXTqnXHUTa2GoQcW6mM/cMx
y0q9qn6nULGI2gCM2mltLX0Qk8OuiGGSJIE3XLQc4bVQhqmbpfjnFfkUIikyakP+
7wO0o4eeRuLPGytXVKI2X7tUR3ZHP6Fd2JGFPQtF1JApC80W6IVbYMoJOu6Q2HiV
ry4ZXJfop+V1u8VoAegyeXZFvrs+S8VZSsC52X4l1hH8vdXbGKDmu+9cUam5KYMT
MT9/wJodkzTZzYFDNyXDwzElZ1n0/OW86XVxCEpi+pwGBAi5HwOdb25eA/QFEK9b
WJA1mR0bOGeSy8NhQv9/M5iVvBWUO3Kwo2anlfC+cBDRlGdRNVjeRInQpBdfVTWv
ODDRxIl2yxIV4dW70cUM+tvb99cL02P6z4qAAOihuqI6gTzOrg5BNSUQd+VXwKaB
WkbhcZhiyU6+90sYa32fMTC9Ul/2cWZ6Wcl0MtmetjuTVnjK03SPO3qOSf01XK9U
JARJyfMMy0HNXyqsIFqfVo0Z7aJ57cxceJa/L9A+Bde0hEmKyvxGoyYm05xX8OwM
9AvkqyWemEZQqZHLtbiF9AFgvMrnNAvwccvbTsHkiKJLSlkKfhHcXv9WAFdczmZf
Qsb4jl6PqzNtwzVqEbjifS4yBmSvVMvTxemMKEMJFPucpqtcSwhdyN0dcKt52qiz
952Yt0E3AbhWlKjeV17qy3GvzXXBYhzevfSyzIEgiGpni1CqNOyMXQB07+1sk9hd
z+RqyZrGa9hQNkh57ZUwAVnSezVu6JLWWVTYbDXCFBFjkhin+T4o3n4f8QXt/JnK
JiMr4NlYdhlESpP1rKb953mPogEyuzGNSqlA00AoVBtwcLyCoKcxmjkLQ1io35zq
b4XsTU8pRc88guaizaxeiKlfdulPOkk2ZzczDk7hiapuXMjG8rWWh4PLjc4rr/cX
L9dYbYv+ciTRoKDSNk8kZFhbJV1FrtmvIrVTzpISgxmh82JNuwDbiVzYyDo/Kwv7
ZYAsem8ptHFpHnIN1ppiYcRy6qSL+SLEOGLhkC6MO0FXrx8XWjUXaxO+p2KJW+8l
FEpkyz5U34JVn8T3Dz+vVZnpLzx2q+OnWJuHe2rvxaF+ui6NqjsbFCOQPt7TU/fX
2nlfN4bWWbnZfAJIAUn77Yp0l7gTw9fYwEyyNQoUpXm5JJ4pTCxG4T7Rxr6i57y2
IRiDMGDETAOZOtYWoqcrTVB7KzlYDc2qrfxO0iR71PFc8+TLHJQaqR03M1jWJ2I+
Wfq17/VlxliCDGulaYJX4h9VaMRFVFAKziChkwaUhhv8uwfLbRGJss22mnJhY1zz
6jM5rDennh1eCPRlE3c0+ElJ9+Xzha/+8EWlTA3FWBY4a/JYvXZ1jLNTqXEPECpu
V8/xps15QC6X87KBZ689i2tJjEfZYbL8eWwH0kEA3EJPsGLlmobgg3dihYkajHW7
aVcCcfmtBwSAHdk0JOo2VWK8DHHvo0l53A2QGS9DjQxR8Op+t95AyvSNaLj3tUq2
EeLCqnfbnxpv4tql6BBady1yYJm5lmYJl3gKaPNmpj4Eh+DSzcaL5LvxGCk9N/Bb
BuMvSWhO4AODS8JOUBMWinI5SPhCVyzR6z+ua5uCVKx5hhuN4YZemiVyF2DaXWQf
Xf+bXnFeSfM3fcjMjGijEA4CkulQqfsKrWOAOkJUNBdrmPJqUfm62s0ccH9/K7eZ
rAYJ4fNFeHp1FKvQmKVChhU6iujkinnAB+hLkNP/b2uA6Z/3zU8FfEcAoH6reiZq
7TEueUDA4aUXMcJ12HAANN+jubK0kwCsJpEHLEGT6gHztL+mV3ap/Gt3qC7ScjYT
A66owIcy/AXujH+zX8m2iWaSLC4kTXsU1MSmSyeKXGUJZTeDlu3j/0lUC5IKqRGA
J/LWOz+xk/AUieIa4p8nW6jMziwzd9DXnYc0rfDyW2GZZHBL1NtR1kacsMnxKkIB
ZXu5JxL7p3xEu8adO6+mDhiBwiLVb476iP2hCW5EdWwQnhShu/BpWWGWDHh8IvlU
woCREZCO4xOc72+gQg4z9/6gw24UBTuQ2SLv4kB/ZQ7eAQbp7xWETcfV4xDdtxc5
t4rYk05F2+8f4wedGhv5c3sI1rfmfSz14saa01jUSeKuSX/utlcty2fwPR8kZFA+
wAstng1kPfa01tHGCo4maM6Q6Tm2jZVaA9IMU2YA4JicvabI0X0RSC4ibYdHASU/
i/GnoQ6lzev0BrI9OODmLNddAcFVZFZ4NT51KLTVdJ0F7abOdSaaajd03Q3PuziH
gex9jAEmbkKqLYsYoOZWdKf7EApBo1661HN9OstRV4hRaQgJhdbSmmm+SckQT38g
jlLE8iC0Q85NT4jQWkkirKRGLyCftOOJgYWPTbXgEC6swZEZZWn5zDEfp0dNPyU7
Aj55SnmlYR07CWT6qexAEcCYY3gc6Vsri7Wr6stLNT531uEVsKI3TTpsi9JZ7stT
CEV8uxfBLdojO7rzh/UpVDeSWWt/nFF4i2xvVlDazVwUI1g0sftj1bTOwuL4D7it
xJwopTIQmo1DH0Fq6ZLSgyEW17YuSL7zsRGluJvUeou0Eynz5IKff84HPtWFSp+Z
/pewQNVy8ZisWJzFuJy9Dru2cvngGH80JueXO1cUfhkTd8hJBa6NsNvVcMcrFC+m
dZNhulEJdJO48MxlWzKHFe6QY5LCZ+DFXrW120099Jdn7lUV8H2oI9xrK8y+5jXP
gDw3Rvsm2DlNbIr+8vb8j4qYupj0yL3rX8Z4O8o/L5diwAwzcpIPFW3R5Gpvpn/z
pMYwTIhrkw3Ar18o7DhziYZPQOKWEX4XJ7VvtGdjZtEpCu2vsRcPSLN6dO1i8D15
uwsOApCu5iToS0BBNAYKmn17vG3YGTxM4trO5b0EziFePzDDlz9BM9xGFvwniD3I
UZoprh+4YNtRPaLgh/z+GrxQPfag+HzDKJBYgykX78mZXCu1hmd2F22YaRhpl0GA
bpMTJRV2H7qYZeZ0nV+yECoZDn97VfcopbSMdqPTQGFpMmNFsOBpgoOkROu5tt+c
4N86IMLUY7OwAAwdROICgds3XBKQGwm4H5d/GWEcWCLy2z5GIvKSd/gdXOvodZFX
55QmqTLQZL4+zN9ouxcRb/OpM8pfOc8P9hnEciTDC4BEqPM5rq0elanAVq8eFVOD
HvK6TvdCd4TDr2lFcUYX0eyzYejxhWNL0JaH4n9yXilh7IZnajKO+bitrM/Qld3R
yK0gj+zGkNmuQmhUMzdZtUhNZI7Ox4RPEtpRxRrNta15McMCxZDcFwyCu/bSx5Or
6J6kFdBGMmZKn8A5MgEzQRGpB8txxxjWgj60KJUSITEcFbdP9YYgW4HfHAhKczEe
Fk4QoeYmOa/pEoN8SMjo38EBO4DrnjUNo47UjEvw/DkXLcAskSbcseNTBCOmfl2F
+DiuNiFu4nWFw5xb4Hdxl+3OgOLl2NPU1V5b01tDt6T1VY0vZT8dKMlpSBcgs3Ri
2/kucf2nTFDRfNr/a3KiGwwSEuI09NVhS/5qXV5dNi7cYeUrd94Uz1qVzu1LC9ys
vmm/V+0M+p7GGIa5SZZyp8ipu3crDBkG/7G4xoHXDbdTuAHC8krvWkOiXqKKRXW6
XN35XWm2mDMkXpxmAIPXdNX62g+Bl/3yTGDllmF47Wanq10bD9pymfWpRx0Tmn1j
WA46LO2hknzd5z4OzOp/k6diNTsxV3c3VHT5tMj+O1QYsIt/OszyDEOBCrrngUgO
XXVam62ryHPdQijsGseiMJhYnjTeUgV40WD6l4HhYrHCtvlkIz6FusNQdiKzFPNk
+y8W1moLn8Frb6sqM6l0LDC771sAp8Y1ZHejDrGGvRNi2GPrB3X5o8dhfEgSKBRT
y+ePre8rzWiKCivFAqOQI5K9fajOcp0aSO/NTUgrgJOfbZ86/1NSS4geCd1CmCtc
05SFQn07gYdI5RdWh1yAuOjRDXDlso5OrX//NHxLJYylt6bXfU9NWahGzoW39N+M
eMTGovik8mq7TyHI4tXJO6QytjVOZ/LPiftl5XCicMD7qhD79Zm1IT6g5qQYjDbu
yAmTViqC0ad2QeVWruLbWPjA8Pt1lSpg8sgsj9D5lHbSLda4yE1ynD++nm9+o3uz
9++I424LE90Cl4KAMo/EYnYY8Bt1JGpo+1cI6wGzGqk9jRjR37+dOhnyY2/5Oa9t
jeJ7U+Fxhxd1N8eVRDHDxiH+RF+mvBLG79tqdTJ3B7DfT/xYHax7nLE3K5NRjFmz
xFcOpG4mDERG3jahL6V8g+s/duRvvr1IxPAZjRAJPf75Nwq/hAJ1Znr5e5Jl3Z0o
i95IZgqZdvUfG9waieck/IT8w7wHSzRFstB7jghJd1X9O8PO2mnJb59q123uUIar
06YRHaySblGAJNaCS7ZXnxkZ9d/C0FMp1/6NmXqLeOirkH0BL9Z7SNw/adqIwiDu
WOJjJ+MSlCqK7KvBZhUqjj3OEHAMCJLkYTcEr4/axzaFviN/fykFmEiUBGtYDbyw
QcLK53YrOuAO56BdPOFPUU/phMjSVx5/AS02L3lZb/wWfGWS0dKB2ci/HV1Sx9YA
DaGAa48R2yT1Te3pdFX9fvLSC2BcubSq4GtGbhZbZj7onzQ1iYqXt9Ph23mr3Z4i
btJB51m+5Eve3fbceUNyQ3unHMZi93+/Xrcxh6ixjQ0/cH09zC/IDD5cN1l5rxuR
ix4+x5LOUjH9qmqsKKE5v7/T8iV/WCRKjlnZ+ZBnqe+lexOfUyctTdDlTvufi1uc
7Q/0qknFk2Hl96G+X+w/S+j0qTCUvxJAw8Su0b0pf3V/0UTI+qXw4vjJk/L72+wQ
MLyf0I60zOvuPOhMjBbS98sdIhgsYgdoTtLPTlhdDposO2nSDGlp4OpYKEOhEh7e
xBLL4m7C5YDvc//JoAlK5qRxPZbt8vCK5kkGMbqR5OTkPQlZwpN3fzJD5Xh8qZwE
yZ536tExRakUnwAKRJfS54WbXGNU7vjowo53fzmn2TuumhMs0mYcvfICAWrMx7JW
XiSLEMvH23sO9m6ciTeLvSbt98ZrhDYAvlYdp8vGaT8FAuwFQa8XJBLYN0Sz1Vpp
9YdMTDgNAQuTn9W0ObLTqnu+zTRWnIrU1ckXVOZRqKPj/93HIoz0v48IPJkUCwur
YkjW4OPFVZ6us2CZJuokeT2cXgIOfJquQ0SD4yypBPSeJtrlkwiFLWGBEijFSNbJ
8q3QdVtpd70qd20Ry7CncxlFmsFq5AnS08LicV5CSMpgPbR7vJ/vuLLccRYy9DVP
qE8kAA/b+iQqZuuJIbO/h9PKuMtSgxfLlr7TmSt1wYrgI8QWaqlw1rApOxqomfpR
NELyHJVaDi1Mq5no3uz5A+XD/K0eAHAYOaOTYxMJAtuvcZ4bUrdJH7ejyLmoOM3v
VUUq9P+uz/KvVKuRqounG0Kl8rNI5GBjMKqg9YhZQg5tb8n0e0VYSwFE4p52Bexs
Gg1mETALPqP9Efdz6Vz/+Scd2BEmKVgOoV1aIoJTLlHvgJTkGuNHutdZ3Kfa5YgD
Y09nt6pCQkd110R7R80uv0GkryPHbZO8sx2UbKDj7N/qCBtXIot85WKnd4uPfYZ3
43+GemunYAClmAuhtFkupCYgl///GF7nDcE+85hwAVsabCA3DIUqzehpamifeQVB
cTBhQXpm711sozj0cTVtumS1n+dDYqDxvBAwMKss/XJ0DkZSuJCkRZMWT546rood
+RyUO1Ih8kZ0LsV5RIyYC3zCkw2EvTLCWOb6XWnm8E/hwwvhJ5/9rv9aTZkwHDZm
QvzaYugvq7bTobSpj+W7sHLzXs5TQbpFFdYXZO39yGXvllyrdxhqpaxvur0+WQye
Q740JXm2u7JRnHfpdwin/QxL/NCSivlT0KGtTMpmYHC+6H5nmqr6DQeTGgLIdkud
ct0GHzRhR4AyiMwXce0GbZBtn26X4cNMJ45WY+B7URkldLVjGbhtZ4a4PwO38ChV
U+UbSbTTHeJmpRbA04cDE7XBNkH4kRd01KRxjYNAeJHk7EXrreB+PJ93d0T0J7Rh
XhZviy3k1WKhDseJnlhFTcLuw/P3NHj3fdl55yN/wDXWuVWY7tpXWF/DK2HUcxHX
OKwrKzSH+KPfMAlR+MR/3Rm5XKQAaYG28gG4CKpLN64r9zVaE7zOSxL7RdhZAVm2
AtFuGa7E5/eytcYWO6jKCbTqZc082bqzTDQp7zA2OXRXOZ8uFeEEbN+gNzFIJdD+
HIUA5e5YONoLVOYp8NfFgeblemtah7xF672BjTbC0g/1l1KxLIwCaJEHTSDMkZPU
ykWi79xPiRBWa1QzYfPOUg1hjPnwKbjhyotKcZTCTrpFWTZt+42Vpkql5srBj89d
FvQ5Oak1xmCYEtgoaBWuLhKCLeB5Zr23Le/riIoUSGyy+P0q4ZJ2YOCKeEE0q07w
Gq9Ly5EgGiG0JTdA9gtAwfhh3gGU5q+gyB5vnS2GhDDg7WlC7Z6nU/KTizTT6pGp
YdX1WtgeQO10lCC401bcJSLTY+rhp3l2++x+grn7kxp68iutOkhc4gOZ1NcflyEs
vNznzC6FG9IAHLMRnXOs0aySHibsa+cSqkfxYFcrx+809ZxlvyXuNn/nAzWnAJCh
Ii29S85cNOFHWUNPaAdnJxh3uE0FXUsDao/p7xYqwcmB503IX6y1cba3fNEuS+Cp
FWqTmjIN5p9QwyCjnk4m6wo1dNyfVVFlL9Kxet0O3/R63jMhrFN04mVKQiHxyDjy
R9LqnyBbgD6rHnnoLAoX/TZjuf+s+6xJI7ffZexBXnD0lUz7ziM6jA/RPInNlUGo
NR0E6xp8XsN6nus8Q7HdD8dOBHZE4vUOm1S3TXfvK17wQqu/dnnj4VgWE6bNz2HE
buugHRKFQ//A2+Pl+XJhnCofQ5qAYQ9z1Kka4BJvwfUyJKqdf1lJTPjilA6b2NMD
0yiUiU5oWL4OWf2v5+sw6BqJ71ZOGZm380QbpcSwCAGQzryiKJ4Xe4yRm+tnaoJj
qizEw+/wcq0+IZyo6TO09vMNr1yzjktenlaEnUgNQGwaTdYub5DbHuTIkQi9xizd
1ckMtQ/chdyQnbL/+z4CFehFJEnHCUiMw4GAk0LzKLicuJyu/wLWJa6dBcqrhr4Q
kvCLmUkR8axFphHMh1vIufRtYBEtmZKS1FIZRVdnhaInFKmY4v4GgUwgxGvcV24Z
GVTnXJ4ZmKeBgXfbdriWgyPRtQep2hPT0LYafuM83AFyxcJHf9qgnpxbn1fOI4Ck
8KRzKwvhDqVyZjask2b3NlX6MC14sA9gv1vNkaZqh8Ixr/sgyb9t5PONNtoD3TiM
w9a01GEh+XgNzhztLm6zcXrufSGHAj6Y7njxRUnO+DNQm7XqaxWL//aa2wvQG0Tw
b2Lmh2peQjClecrFCxpJedg5vYBY3skZvcVM9P3UI9ryIwcY+MhRdsxSzHIyBmKv
jSwrpHyiO3EqknpTQXO4CDdfna3vZcQkcIQsokm3vgutTTJErsMANir8ac12wplA
bQCYt5PKnEy8uoW5NQbwG05d/n/kKvqxmbSYJxSg/wZz8xPE22d0/a162ox7qNlM
ybaRL/HUPf1TqDB+hX7K7242getChJbWz8cvEZ1yMdFSsb7Dv3fzzmS7SgUopvqy
7gpa4B+ih+qPwzCBdiT6UqRkmC1ekclyjJolluKWBrk4pz44+9Zmr6e22jzOJJm4
8YKLeyZvRBcRWRNvxhK933cvsA4keQxsvJQfyFp/GMPRfZmc6Z+Es6Ehawt7uMTB
lZBOg1v7EjjL6VVrVzvFrT9GuLaz3AVM4Ejw7cEbBQC2iOsSyr6cOG1vmjnyJV2z
ngfnwioMyCBkyQ78LI5MU+uk214r3f4GdtN8RE9owdtIV8t2QIcLieEenHjhYW6i
DEz39FuEqg1igwp7I0irc6SWU7UKXa5U9tbMCHsRYrmQZQQJFERw4I3d0AieVsCO
8HfCpOeNZIMNkWU4lRDgyqdzXQz7pBUcRNjfIzlwgARGm2cfxubMkqevfc1G870r
VA4gzZGjZMIhaFqF02Kq8Pcxf9A3evTE5SFrnlvUvvMgLU1zdm68Bc06HNIgJ6pW
b7kBBAeydIMbsCeywobBoIQ8ZJ/dWaPnVU5zshSVIp04uf2ld1P/w4UOeqBwdDoD
sGLMpuRrGQQ2JZLjRFHRy4jyHLTW+1wV46b2ufjGa70V3KmgZbUFlP3+dbZVddl2
tqW5OklReaCkRpkeR76MEsV+c68Ngt4ASZTGJca7JvxOd5zj3iizIh2NCOln8AMD
TY35hFfHNBYTmkTGK0Y2IwcCAN8NsBEXbeqGMtMwHjO8sk+k8plCzPWb2/v2Db6t
7dNrNoxy8eNJpqvZvI5+SZWLKEBpoZovAOrIT1eT6DDkBBaWlrhci3WVkPZiJzfR
39LojwaE85bRhJsZjIlwcpJArC4aBpFDRmCbXiuseKOnVpaPEzpyojN10m1onjxP
G+0T1HUcKlfGo5u0fxql9aD0k8kExMhTGTUpdpPIxdTQ37QJCLeXkIAYGJAs+lll
A9b0oZpGoenyEbySwvy4sxIdxG/e/TsrLarx2+6ErnRRzoPgWMs8wcr3byO9TRvr
ThSkrGYPSqYhrG83fFfm5qrOaUlNU75ACoUKomeAm1bakX9Ma9NmY5pq9QZvyQpn
D0gB/iXeMv1HCkoD1IAOpKioxnz1xhmDeYBn4WQjcejleGytRPm1FVNzhleO496/
LxSxdq8VwUWyg74QQxd406sJ5yjvf5T47+wn/3rvSzFzf+wtdZ1uvke+/RXKxwpl
AHEn7IHtLgkT7DHLweVl5IMQ3ivkkleB5bcGYN2E3nF1ggIp5KGjfsrgfkHAy5lL
pIe2/49HM6euA7DokU3F65S6h7e9cMSDAaWikMVVDGWO6gKKcFmsOcJKnR3Wq8GG
zAzWTI3HV2UFGQ7smg3N7nbHvEDpYDwFzV9yLlBoyCi0ZDfr/p2TVEgHplTugeFl
ikyFBUN6kVtwQ2va41piZurWYeLHSUhlPoCxC105rnILgl3muMWJ5cTBTv65pZEu
GQ8hZhuR+unxnZQf/QQyPJQz/YPUgQPWpZtDyRV8vBJZVK+Acw6W/Rcm2xgI+oEE
xPR6t2i5YtW5d5oIcLk6FSNqqT+2icANetsaWp5ZTGIGBWXuITuUvS+zqNbkwDRF
1siI7SqUc9uHkvgprlbASnIaCRBYNuc/ry4+gAvmpYa++wuY0WPjXuE+gtFNKT4/
AFgTSvuyAOuhxsFSxVNRfABYzpS6RMaRzmLDkq2iRGLu0mZvuXajXBuT1Rn89YDs
d8uG0Crw3s74KSJo7pyxmV6JYhNBu90azsF2ce1UwpzotJo08PZbtFY/OOhN+11Q
sy71FP06eZ7D5SFcw97KgnnRwugglsOfaHGDi/Q+q+NoSSynsYwezLFCg7YdvBca
Hfw67CInkxNDF/BgZ9VYci/C+uBMeutIISCdmmm9uv5kxHQAsxl+Gf8mFl2Nw4sn
4sSEiqCfuaNuX/rmFz7J+Bt4jm+X2CrJFSf1kvivZXv9IdVwYDL0nclSiHrBuagD
Gkyfaqoy+vGUT8XI2KXilX+nTVJE6ZZ03xM/dS/OHQMGDRzoOhlx9o/ZlGJlxHir
bHA2BUiZnrfErM9D5EppX7ubMDsWYEFl5Mlr4IpqZyN7asDMBJptqo87La8h+OOs
Cuxiwdoxts2iBJbU4Jwvh7V1q6O4JHbSNY6/OBSZcCMVHMo8OHkgxGe9PDRXfsz+
t2Tyu/APNPE9fb/Lvz3ig/KLZyiWtxbgaZV+fHKG5IEQmkocUYbSgf9yaHnGlHRm
zYrjeg1AOOIGZja2E406JLuNZLPuHCQKj0tAUsU5+B/iFsfmEkv9iHlaBarT2mio
QdsfIzSrxcQqxHCiV2HVDJCuq2vvzkUjTY1RAWf0G1cwIjGUJhcHrlkjOINYN13v
00qQzT6s8KSkWSoNNEM0G8JLANdUOzZaVnlWR1T135uKeCZnwyC8mf/USaryByAY
LzxtQ+DxDOq87Pe4Q2A3njKEtVHso6BeSKopLyEc/pzUBiY0U9yxVNk/pe7xS1Ly
D4nsP/zgIurtvOYDF/GMNUk2IMC8kRpajZBFTXV4VWR73U/RxbXFNBLLGciwkVMn
r4BzQqWCKDqxJuSDoYplKkn/0JfHgm/DbRDUDW8umlkm6Lp2h+76PTjdm2H661Oz
G58aD2iGZkGxlt+ynSYGwOKR/vTq2VaKrjeuejPThJiHyTuNnlBvtTaufgCGFbH6
uaCXU8CRCfavXyNhKygqKF2Qs8l+vKvPjDVWsqi8zv0Bppme6mzkUcoqIIIBGRwR
GCc9BR0Zq4E+Mp3JkCiT/ya0M925i1oQs3w+djZvK2iWehpSkYGupTC9RwtgDCB+
AEQrm+uoKyk7wmHZaxTgxDQWpzBQ2/UOmdNInbNcfwrKCIvLQdA3InmXf0KyyGTu
7g7CNsx67TXJWtfm8QVGlOttuwN5t74NwFCU5bB+61vtmcKXsnW6NUwdk7fwgbhF
7r5dCheTi4scHnRSCuQqv1JHa4Fmdc8dGVLi/P/oTH1vm/NQeugHK9qWG1OwIXxh
9jLprOAU5BLVKO47niWExP0Y/QliSHWWqhcTqYoXuKWyTBVvub541g7uTyagxDiC
R/LNyZJ8NnZQTezYvY3b7sqgZPWhk+IPoYqEEB3IgukqMJOA9RKzJjLiS6BicNT1
pntNee1fD77xRm8+ZeTL7Ojp6GzMM756g7ralslGXOP1qTsWxuGu4XolaSzIySgE
EIL/gioTQqeNeyD71yigxsTiKBXPrvqcIe5per6NzqzEl9zWx/Ba4i8STRbXAQbV
uCz0ahd8X7O4C73M6ZZlODstqAMYffQIi7orjwXY5CQdvl5ajxvlXyYiu7thKFi1
tzWy/Q6B94FymaS3T1vqE9wGX9r+eTeoX5fJ9CZ2lbilmrQ4adJqJEp7aMcfYgIq
Z5HREMO4qcnNvHA/e8dVe4QZQYHCYH1YLfkoJQxszQep9wiXvqmrkSyiiSlfXdKp
COayigvTm2EUpnJmCpSKR0eOFoHnLUrWr+2Mpq1AOtY6H21bjOZKJhs0iaA4hxjR
PDrF1B5e6Rq3kBhTmZlpmk/26aQLbLFJ5FmYvdOBLBCuRN2HihjUJyc9KkDumBXD
yVgFO4RZ4XDf4YGLBRGGE1+VOOXVTw3L/tMeSO566549oWNXKe3qLi0vb21Vub5B
70ZFQ3Ig9m7xlZ8q9fn8yZSqzd8Z3acn80H8ugJRKRwqyQHVsj9jSglQzjYd5ium
B5zeJtabJ56rmUoXt8LN+oFbdietm9SSyXWJafHJEOAGm/Jh14J6fehVdpRGYYT3
gZ54gH4MbEnOyGIt7G9UsMf+bD7CmpYD3pNdwjLiX5oApVYrphMOG2qfT3OEqCZ3
e4nUMpZNJdcN89bRdN6LB7cRnlp3KHRIHw/ndNDfuTRqx2VpsvyLeYOPyirVz0wl
7mlZ0Gc7gJWq85GCAoyv9aC9zg7zx5/OjojVfHGiDu9hnmfDv3M5K1fztHCoaguZ
WRzDpgzsQ0A29QjeNOinxnSuI346NnTHQ76z7WbqKSiu4GTs1Amh3B+6QKN/0H41
y4IrpWI9nu+CcMW/Ur3glzgmMLDsN7F3swSRY0IdKBXFo+LvBzHYqmEvRXafdd9J
PYhw6ZkBrhVeFUtTEgpOvSODfI07S7etO6Ad/1hk82mc/J505YbJz/Io127LYVg8
Ny2PnOiYUbzpruJyn9SHtsEr1WVQSe4ug7/cFUA2hHRHz/AXOYmJfq3AE6XKFjCR
sHEZAgfbhylzCn0tYfziii9I7WxDcms6hjCTJgdzIP4oQVHK9fiknxxW9LNktIj4
AcL5hqLkB8u5uv6co38tIHI3kSHH/5WXoYHYvdhcRLUqFGqCXY+6GmZ/BVt3kPZg
Of+Kla7Zy2yTeyGMeJ82XqNPR04ZqxqdzojdUvUiwuESOuF4z+cXQoTNO9wpEFQQ
z1XHUbG3pxSdCYLPMRCNUJTtB5+bIpfTwq6pNXHwzVFL4nJ8DtjpV9T+ntYo8iOH
7A+ZSitvpCPSZkZGLusb7sTnIDZpKhmuUrbfKMxKLceE/wkBEE2YdnmY188PUJGm
exFb52JEB7zyO2jK1Hd3pqARMIy4BlABoys2TRArPs+q5wTRSGbq0zhSHx8B251I
+4MVCGvATZkAyCv7a9y0GY/FjX/kWHkd4486bBVex5n/Y7eNzaC7eVyRq9dsIgvi
pYWLaDUa7qkJSXljYZkvnFqUAN32caIGxzxN8Y9jVPiXlwaYCtaB1KD47Lkzv6VQ
VXQWADUeTDZ1zEECFxxun2U/sWh8v3/EN8r8+DpEdmC+lne0upZ4gAM8PqsXC7BT
o/4wgLj5kq4yRu1DTMweEeGObpwHhEYzPp5TXFVu16plGFWxrwFk4GXVbRqf7dxy
HfKr44OticPfzR3BrM5S4hK7SLq4h+TrLkqjZ8LU7ErIFcDRoDWFlhqPjaIrTH35
fbkhfNhLu/icZg9ZZDqGuWlZuc3ssNIYdd7kExGSzk/EUKAnB8RxrvMlDXmM4krv
Sqgy2+M2OCDBLNwx984RB0hyyLgwOQeK3m5GlA+IkmF6OxIC/81jvKzckdHxGXN5
uMRn5Lks0fR73+pPoYmsnQ0j+C16cDnvRKDGjdn+I2Dg6bj/8C+N1/dgTogen2SI
UtHrciAQpIUARyeYNRhQ7Br1xzNfmDUudUl6iE2gaofyqkrGf84zRy0jvob+xGhJ
0b0Z9ZynuQR/6FREb8Rak69wiSk5g2UbgVazl1ZHzMh9z0LkT/UgBxzRtMURAx7y
ck1G/e7dS9XcLnm0PpgROWuMjAyn1gq85eS+SOKn+6nVTxdZH+1A+e+cBLCCEaZq
L1KX8WE/rTPsTgecdJJFmqY4uWco4WQOwR7GzEdv8PB5VTK9/gi1NshqKqwVK7wo
p1fcnbB4Wqf1LCgRdphbBDrYAx70xed4UCi1jPlq4z40Lzf0AAoONbzmveQDIf4k
lOj6bsdpzQRJUmExm7FAiEKgm0mdDniTswqgNlO0hB3rcdzI6zSAyDZue6uuGbj4
7CgxaJSFBlWC7gY+Tl8cR6GbfzqmmkH+JNjF25+wAQHbvLOh6EA1dZacMM2j5Y3m
o8jiaEeYqyJow1njkwJAeGFRGPDsl4JFcMPiKvPGXaelxl99sebR/meICcvcZSkt
f5pAwDTLisaBXUelCQ8LkTdmje/oDR9Zx3xxUt+tWUbAvXpkXmD/JdHr1R630IZg
DOlHcgfm5IIGR6efCCGJaHstEXLghPNvuyIqWuFGy1Powu/4fXzJFMNOXv3RlsME
a0pimSAYjY7eRaXweNJ+u3npPQHJXdun6cqrPWs7zpnNYQPjkQB7GtzJ3yxsSQzM
MfNtyNLVfjCd7B5yKL2VoNtNmGIyD7wddl9i02+BB1FE5WjQW1Ri7QsQpDgxzv/H
V9TcMC4YNNE4imrlcfjeJjyaPa4HbL3WXEdo8psid3Hz+WuD3JVZ5BYzyXLSpfm0
3jbCwg/+n+eBeKpxx8/Txnty8IlWsBpSuw6sgDjA4E1McbzwoQnrNTLQ92Re/Gvz
wTFexgUg459LrxYSqPurLEP1+uyiPZF+6WEVI5FeH8sqIIq3n83e1c7Xs6rLg7lw
OHPIHdP8MAqZ45HQPE8K3pu00R8vvN8iT6f1yLetZ6AANzdc5iwg9HjN9/V8EwAJ
IYkOMauKCe+BJvlW36Pnekhg26LWjioofgmZ8h3lTvT5VZWOLNk9g8dY/V4foANZ
3Z2uxEFTOzL7gJqO4Bm2+YuRhBcT9L+1VbSgzwuDcj5gbBPGhvQNKS1H+XpCR+bx
mcQGN15E+kfTWCwVoicE0KEiFu8jdSm+4eNp0Km0MHDUItA53XmQgFqkezBWfxst
kTXydyVts0wLBEmZULodvrL3MlkL2CsLOZFKMxGVVWABG2cjNknhgh9H2HWp+CQn
tqdIRRwFbofAv467z1tVf3wMBdC8GluhyUGGwwRKETxMliTpXN1Hqmp6ikbhXj8r
ekOTMHPUNu3GrNQIY9jBVRu+6TnCzVB1j9AzRhrlQmIJGADIVq3laKYxbmginGr7
TKjEuTMq+NoP3Bl3n33wtEHAXDRbFHShxUO6Xv+Hs1FKNinVuTTQRjmRjoaeuzWW
iMiEV04Kj3nWfRJMzb5m/Be7vQJAQjjWbQPaK1TmLHLrASqIWhKtzPJKyYO47P2I
1PnMi3792YojUKF9V9llCjgz/qEDBpyXAFUyabgBMcfk26I48EZOaOwQY23pZUIH
idlNmbZjRLm9FLLwyL1u/r+n5LoXcae43k1tpNHSsjDszNiHA457X6z8TSDkU7ou
/cPVYoZxjU20cU2aYBMizauch09TnnTeReKlQQWZl0OzeQAmXKKPai006D/rXZqk
zdbQfGdfqn2V2J6SteXG7Q2kclcXdGom1yQbu2fd/sqGD62UIBBRABVfuv9xyZhp
2bhtLDS0WjJuQUA2UgsKFo+TueFezGrtr22xcc8K9vOxfxnqSRoOPNXTb06MxcyG
a/jfIvmlw3mYSY9bTDl5zMO0drC0asRdSsIkYPqZlTZPPXRGRShbOaQ2/ZLkgdZL
EMpgot9So9arStoKWNFHX4qbjP5KDbShGC4S5fShnT6FpPOkLnZ7NWqcM+g/Ghcd
v0CwXwRw/VEcmIB1KfNMTCyi60fVTf7DXBHy7JVk8uVmiNRj1A0mg1XNrVKE6pAV
inpsF3d0LDpFfsijVnMUocB5NpB4Ef8JVml8IVSwWF0LAoZ0PSIGaqwkgRpuIBcX
l/SaMBLK96IkaU0m10tu4I/kckS2X1ncm88b0fqVG6TVUReeshjWyUusjSfUDej+
j4kzoh9s7WQS6lFwaiolLpLrsCacrcgni433yW9AKTUx8jPKYG4/2/qDp3cWP+s/
/LBx/dlZSMFygA1njHlSJ/75TnM2MjUdoxrpIcvlzo32P8NhjyZcxvQyMr7doZhw
T8YzmdU1FIl6IhQURbbDlqN4SvL6vJf6ZJthMcXFHJWDj08MURpY8D1nxenO6q1h
tIlfzPa2r715cIUgJ2rm5nNWPMhQqjrsxutjCZ0RJF1+oE8DF1dB688N/nyqVe1S
ej91Dla/PH9I/IyyaxwHIJWInkJqLirU4+0UdEjHdzgFAV6T/isVDufDX6uQXrO8
nK5BheVmHFUnXhWyEXdO9EHjCXWQ7omguiPbkAv6sV1jTQyoCf4J6fVFQt7VoIy6
7ktj9hGq+V/YlLSg6utRX/zUBFkDgR9qeEzhhCA9gEgu4sMDlyVKl3fh61H4x6Kt
LVPRG3FM8rBU3SDvUqWZ55+1gzW1D1iztRBVmcaPBXRM8RB9LGa7ikJ2vS0aNiKZ
ZWNPcR+LclEzItX4moL1ZcdDk8/n+3N5lYWjO2YLn2UzJxt79aOeDcA/ekKZp58d
97ahXTO2+il9HHx8K+Km4nOzsjLPdYLDxjcLfXXt30Yosl9ZMqBoLyy62eyED6TT
2hSrnD5M8VVHyUAv402IhjHrAEnrkt5SsX3ZQvwQGKW47cnVxWNzCblPQTGLwE8P
k9oXKy4sa8jEBmeaz10nym0C3s1QJOuYhiNxO3/qb1N92o4Xb/pN6tNogup7MOOa
Mbkd0duH7754ABXQpd6uPJOdgr6Uf1nT0M2bRTCvxfHZg+ECGRb0YieLQeptmkGE
+MD+1mHUjXOKTHW44VFC7bk5A6P2XtvfKvJj0kutROE4+XOpA7lgBqHJRuxM8Jd1
KQ2ZCHg9UskE0fisH+KgW6smBJf/9VL2LmW1mdcrwQ7F8n6Y0iBSdW4FRou2L0I5
Qh3tE8NxVWYguC5qv0yhwUa4PmrPzWjQim1jLqeJG345gzVybta+r8Lhzi2mBelT
XCEE2tuM+YTNSdBh/bjTXZGDsDkP7huH5I2fBR/IU8JVCSqGwDHJlOa23enToa4W
PrfC5fU8M+boVYAjA6hS0rfBuPU57GZRZAY+Ag12Z/BB1jzO7L2CuqC5Stu+/HRH
nrfZM/CIUp69Qt0QcFP6xzT9Yn8mAGNDrRYlfw2wBPaFmm7fzkZXHAzKz5t7tzL6
q+1AxseRbTVPyC0dUCCpKapKNp5ovEkcrJyXtCDoqxASBLwuGe5+EzlJgDcom473
3rs6AoYcc9zfj3fBk9kYf/Cd0pXFg47BP4vVzrFvgZj5f+Pm6Szw2qJe0tX6HzDa
RW6S+3kjTCCFwNeTvFfM0k0VsFLY/PL5WHXyKqhwHk8sZoDk2tCcwPNcOKaHtC/a
MJbXGmKV3YXbKjtL0C1BI0rapkKt5k5yuxu4UfCJAwfghA7+IoOR/N9KvwFQQIE4
t7r0HjjfwetFedr8V/8bZKmdagYritGoq6bYHd612DTRaTeJ8OIOJcLd3Ey4z2It
prpsYgLSXZg5BlxkUUTOHPpPxH8hiIA4nqu+yvKhl4/cDt1nsTL1WscbDKiR+rKt
XPyPUZYAsumTWhTEusP2s32bwGWNtaQx2OyfC6bzdBwKU7bdPVBtuM6rertQ5s2w
XodPUrg84MZ+D8z/urGfQjUhD2PjlOlCQ8BBKHzGRoZaTNnaHnTvx9AFwv0027xO
w4aGHnLQ12tNEd8+/57SIgU8zPusVcsYQKJDv33akeeuXWp5jKDCld+qqTTnvyXm
FquiDnQAJ9LL1eiSzo/Aa6mJ99n7vvPfV1dq8+8MdBZ7lK1ZV8BhZW+Du++XHjzO
TsaFOSTw7hoYKSizFkYwyIcaS1cA1kKW+ZPY9Zsmx8KKfzRGr/qwh+JJL/clLzv8
aauy0I69f2AASM/3BlFucxDCeNordqJUMQdD5ZAl+SFvMeylgfrv2mVNMJ11w0xu
DOH+KXJA+44sui+ClB6LmmmuD4sOMIqY5OnrwbkbUH3x8jTENkmIFXD87j1N1DrV
55vH30Q2otnJtRnHmdPeJtdVAR8ryUuWcCpmiMeGnM13zf3Wa6hMnXJehQBWrJwH
OpgRbP9jR/mdek8R1nFH23UcRwpJplBh3yMDDcfyOsfLZsbeTgQAfotKLXncR9gO
bNIU26wc0od0Pcj0XmhDvgtpD8/IA7mE8mg1Qez2/QMwzTykexPqu4swnlDiqOoJ
xhV4gTGsz7Ts6xSOHppzucINRnnx8YBKK7K8KP2NI7gr8SENgDlUa6hhMWmg/Afm
TtKw9uVUz3JpaojrjQSW5iwOHCW3cJh1cOumtbmzAZE/3K9c+QwtqTJjYBDNPp1B
wI/V2vmLKF7OJavC1DQinvbdp+2xm/hwQsbk25UVIxpCNipKl6FE5YH2GJtSes1h
urXGx7W9CKpAf0LwQClU2uE5oJ5Q1sxUvK6CRSiRzljSS7EQOvKCg1ku3XfWnIDt
fbAq/X3dkz4m0hd7bHpGAK73lTOz0fxeq2RzhCSf5/Heqlh4pWaZQWYIGcTwBL9X
+iExpryuMheYkZALyktMvQ+AWLUg33yRMnlBLQpV1FwvP5JfoufzLSYpjr0nR5bu
0jG7LwOs6tWid7pUw7IFw9BSp3pPiPu37VImKWNqoRbeKwin09vLYSGKbYkZUYM8
DyQHmJQFyKCByduFRQWZ9ene5ZZ+1epPevxZ6cowXDYS1l9/Aq5HiH9ioN1zgCXy
vTto2gf7+EMXkSkDRvZgwYwrrqCWHycFlHnaRZGNtaWe0erU9pWH8SUhIhGvQqre
1Mp0nK8gchCKTvkRoemH0+Gc4Bztqasnm8z4d4KO9EZUei3yeNO9j9AEpSh+ij/n
NiSxBElnG0MG+4acBsE/tI6I8VYjpiEirWVEapPUuYbcndy2O3IHU8/f2E9rpSoy
blXVnPBxy/+Cbm1K5uFsKXj+xhG9YYTSOSeSwWqHpakpy4/HaOMi+t657Tf8MhQl
JZWsaziv8k/vNYVcs7dR4p+i7AG4VYM91G7ZO0wKHN9Dv5JDcUi5+NTEd0clmFnf
amFH8o04LrXPtcMwU3Wdx1OjFEAGaBsTFN+aZsCPYtQDhAY+ADyy0dHQP5vLYhAa
lEiPxdfAAhyLd12KmfXTttpqzSat5PuSvkerMxR/Zptw2peZJugPf/QV1Zpl3qYY
9AzV5pxvQY7ptbYzpBfHSwj9T2C8nLNGK/DpfeXHFUVDFVMPxZzcNEQ69oaaNRQp
uEgv74373seJKR3To9wYP0WxMp8L/XFjvAaec9kNkxsHbQqd9p5J4yLUnjdfrPyN
abcUpz6LyL6ikHuH4lDhpgg7abn4UawN2xNonVbVgWKPBia25E8lpNs8WcCzZSq1
43KlvoZej7KcIZ9XOABGWClUBXbrG+oTQ266S8nZX8wcSy0HmbQ75vig+pbAMOXv
IRs1qoKEO8dOnh1TohxJZanS36csvtrQgnqo0llwtt41N+hCdB0XOIfSoOuIhxcz
X5ocG/Kf47q+ZtW1T5VE5QqgIUsxJ+TwCdXTMR2KDLWVEXRbzScta2tL58ZFDuY0
RdadgDUnvnSqgUSgJ5ACmE7fxHcBU6HJDaZlrEmLtMyG9W94QVlkIRb4gXWYsZ6v
c58Cg1Y6daY0e9A2p0z8uIGMNUQQRzJ/o/LUutneFMTKQCuUa67qFE/s0w9HV9N/
HlvGeH6fWAr6gmvuxz48EO74IXhJuyPm1e/k6u4L7hQBYY6G333FqITTC9Ia6BD4
CWLARaA8n5W2qKVHK5Zxo7wl3UrJhuc64QBhwMKGhBSWTQHnu8myJxyciN/LLOzG
Y2ns1LDvu9ofPjvgks83pRoptOV71Kxz9ZqJwenXazszJCA9lf3zEeoyHr87nb1E
6QHFSxKi3kXXBhliZ1zEx6MiCnm2RB6kY6YKKw+CeiF+3DHSNMj6E6bAXS3gyUwF
3rJ7m5I/MTYikjEa9qPxtfUajV47sPToQngv14HKuqv4l79ENAq3gOe/6dJZjapk
XnHk5zlP7QuBTjG3G4qFJCGMOJEaqqY05y/kbQWbHizQs+Lr/Yqi0E9VqTmBlv7H
1dRrW2DLxVt4bah1R2Qb058SJgb2LUbK+d6AwV5OC0qwKqPI5+5Qwu8Q6un5rQOc
Hoh34+rBgm5xEetdchJLKcYURtZIEWYtppkEG9jcDcmaFDRT4BV8ZmJ1FHAcCWUN
7JP5hUG6b6KfL17zynQBX9qQjoDmVQM5eJFDuv9lsOb6xzewBlK9T6ItnIQuFZWo
G+6xbl/ZJRvYZb84cKhT3F2OInkN8xPhydFo1TbgYg8/h6yLvTm7T+dT8pTKVPaA
JgsRXPfocBnPaEUjvtZCYQ9pG9YO9V6YmHS1M347d5jZ/jCMPt1oJ5H5Pyu06gMZ
MkaC9nFDQ21Id1NagwFkf8tfwKvb9IQjBJHe+eVliMXiCo13/uBtoZzbv7YLaGx8
fRurbNXrxGTb8CWT/fT3h7trVoi8ygjrgGbKdqfeV4ZuVOKGFy9sJMc/jLe48Zk1
qm9C2/ifnh4SGxK2sfvK/sSGkQmrMqNK9ijz4R3HAvl062d7Blg8pxd29ix2lSk4
B8QevDSiw4RRTgoXVgxVH46y5Cl2MvHZAYaGqXUVhrXDuNKmco2s60scYLE+ZlNi
LFCjOlqdDS2DhXduBzX9qVe7yMY6clNjZHnhheEq4rQU5bdTid7al5i6G6eOQhrn
c9LgmeoRI3XuHmO0TiX9f/m6RkfQDlvG+D9IyV0uQSWeUOeKkXTxdiQjalP/aozw
gaYT3xBzE/7N50HJXe8EGQj1A6V+RaYzmxdfMrdHNZcKXVNgCXoxtuRXO6nNtuXo
t6bDY69Ht42a/6rAg0cd2N03VbhLKefbrY2nTAsq7oZTvcx3aqaZw/LZui0xpJuY
BHf/jPJhPQVy8IsL1y8ZWKk6gVaSQgU7ZK2SEWUL8cJ6XuNy2ovCgvqOfQ1f8q0I
CwbQgIgjzFMHTI9UiS1d0c2Ldc4iAQ+arUxu0F8A9sKmA79ytKkMl7fT+HXv+FgF
sOiFPoRk9q1ZLVHRUcnViyd7YRGTAolhR/n5bxVbElKoczcASfdP48Wfb/4avEdb
lMsxBYeZkQVKC77j4i3HuSAaXV3/fCTyX5xADJ+wcQv9gqwdGRt7B8jvGXY0JD31
lH1s6Navb87acyA2XqDozeph1r7smme9Fl5IrHV49Fbm5YlGJcggVML2ScybFw0w
gYzDnTwylJh2anwYLo6nIlKSbWJ3V9XoEXHfRhEDxs6w+fEzoU6IskT6D9Y9wQZ+
IRjoS/HWaCre2Nadg6OKBwnHBfya6ipAhMc4V4p9TvOXXAJuyWxdf6//3xfA+7Dt
WFiIdATG5OTc2Sqa8I9+Vfyi5aUFO2CmKRAYqMgnfCPcm3uVvHdrSWaDJxYZ06eK
EsSobJTkmSzuR0CDH5+efs64Ioqmew4tPJ4BES5z2usfKmhkW/KAFnUCX75hagL+
m6NNH3WGhSPMYWK5+aDBIOtlcBBhG83X3SgxFeRY2Nt8z90qa7NvasS5sroEvvrz
xY5ohHmx5iAd6qXrFVneUkZQ+xKntajVU7L7F9fLlliVtZwVbazdlmP/vWi0PCzn
5L7qFvtG1r4xWrM3Nc8e5oYejxAiFpjucwaVHdUr5onXXVrdtRjpODcePD3hrlYG
Rgn1+Hrd9XyqQrLWGJEv+mGicxrDZCFRHEg9/lTHk41Zks6DuS9Kr/UJXBtNkbPQ
NmKLr6OHM/RrlVH3h57Jw6LL0qnv95h84DdX0a0FUObqOZzbriVjL8Va81vlFoy/
NkUQBMXNUxPnd6kf06oScSj3NAkM/oWAfRknU8TeZyhpRvVIiuCZMvgwEll4LWIT
Xx/t6nYSordgPp0yVNSml3jQJMekTQipjnuu0Hk8gqcdNM1qenwK9WMK9TXcXfuA
gP1CTSxXmwpsWLDqq4WQZsZFYff5Fsiz0nIkNARfPxW5NrydixGtNwR1ij/LxSyO
BQnSUrNul0bfP4q9oekH+OmquepUhgj78cM7Ulj+wSIN+wwPyQKUJDnHUK+kKBc+
if+STg1PnCZvczDbtxaQH3JlfOYgFyGcUFobEB3mxxcAVvk/Qq+vHRF4o7lWx2yR
os1AO0bbr162iAqJHxnRSu7xB5BX+orsfRg0QaIRLtRMOAreE+10YePkgxhl3pqJ
eWRCsuZ6sSOVJKTMkD2mNdlSnj5r8I0u8R6jikqH9pOVjr11q2IdR9c1KtXZXElk
dSqpedOICtXNSrGopthPpx8h4VloSJjW6lMvc6mFI0cYqALQkJG0/X6FqHda9Wu+
8vscK+DoDPh/WZfnoLt+lDtWJ/TixPwd+gRAqrGXr3LNoAkYF6Gv2FkY9yIA6b8A
9QuW40thBzhzX2B1T2wsV0wDeFKvbftBAEosoAI4f+EVOkvqSunkmdcGnCqTYCK6
0wIHuuad0y4AXDQ57gca5Gbj9hMKhgxSFEsKjf9xLYKuAA+Hk2s5iFR8Bxtwwor7
wpJ2u9OU/3agaUiw2FxFUfXOh/nrEUvdW9BVCNcpSfTAzvqAd/zAlfF/tOZgbeiE
tATBb1Hwrrzlfp1y4ET8VC+nX87P3MLiXaGxOX42UVWc8FUSw9MtVKIHxNbQMQ+E
WDj5mW9C/xTMb50QoEqkU4m1jqizx7FHaaNkANXwHCNTXlQ7DAya+SBM+JpvusY3
8fdcKdM04hdk7/E4s/b+5dx+JBwDrFy2kZzcPg2Lq7z6DIHZmRaAsh9j2y6QvYIb
K4EWzkkbBhzeWlPgKFLy3p3w0/Sr3ESR7q2NA0nj7KLs4BlohKz4xiGASKsHgFmY
4eyakprEZYvh1gJq0/8DtN16AGYExPYktFBBm95qW2pN/8+4zkFyHIvAN1C1cu3r
pUCQ+d+2Zf5aOHn3r7MCktyeoYRpTtodQxiS0tZRQPgOBU9RnzWu8aWToU7AmzdF
HuLzJkzSgcP2BmbikqepwV3Ju/B7yo79q+AI8nkWLs9KbSEdlIiptPLHoV1Nuf41
/g55G2M2VB8mdRsnCuoZboAjkWneSPX5lpgFSXK/6RC85OZQkbWYGkpgZlsIRd79
7awQInFiY095cjxWeyQJtzBzTr2pCtuiovZs+xqm5B2fbXrXzKMTCWFwEJuFIHQO
LRlkf/dg8Ckj14VauImXUM+YI57ySk4qSYYAO3sSTgcJh6B+oc6Gy+s7CVajKwIv
S1x2ssjX9EeMgoV0UEkHM0U8pKjWb39Y+/j6bgK6u1LOCJXhjZjUSOamryHFosT/
dabKVbgyUwzTHH5Oe5p5L1zVBqSZTykhO5Ryqq8g+0YUSma9w4Wvd1aim5TuNLDf
y5hge9sVvEfQzWTX8+79dKscMlICLTMREVeE3LRNkmiVWOem3tbffEfWxk8dI5Q6
6wabjevYmLOFY0FTCV3immXilPdAPwR3SxcxXMkaDgrCUfUErAezyYBDzDuTwxQ7
floxIp1iCDY52B0jv24cEZJa8oWUfSPq1Hc1q1OaWcIbn3gawEY32OK6qiQ7hiGG
4+fdWkFCcdfC4wmIpVUpylB/5RcylWDEG7HPhOu+MbpUDbSMbPNBe4bFGU/eUMK/
JSHY1BkMvNM8BveH4yD0GeXLmqq1LOg/eUwx74cbVxSGG2x8ohbUy656FZQBscpL
QLtaBnuDHXFjJkKsrb9/KDzh42FkRiQPrTNPalFjI/L/97Uknt/DJys16V+oBtwR
pqSdjuJeSwpJpqHQxDoSw6maOtBbb7gX9onw4iHp4NYnHRodW9w8bJtfQVae7Yuz
shWZppdDOFGs9gz8cj93YL2WcGmfv/q6xPrYBwUAPDQMvpJnjgZvS0/MIwxsDom1
UZ4K4al7RjvMXkKHxDFdALiaShBrkrVP/oBbTOV8bFW5jp30nq7jWXs1wyxNdeUj
0N4qsltV2iz8uUwLThfTq+OPr6/gf3EO1/HB8CDo8gUrIJpJERpUapdjvCs9Yru9
FbxAIKnkvmBUrwm3O4ttr3WNPCjUhgK1iOk00/QbYYvvsXSnUjUGDoFnBugrF7Re
V0Rc+bxBcc87VWjAwnDelLzEPBcJt2pr0tPdpYiUIZeVwBlfqO+VJPLwAat6GbNy
PKqwPMD+AzNuCP1B7fzq4DkLAikGWeRGi+m5VT8IpGnbgPba2eLn1c27TmJYXRjJ
LNc0tYpS7O+z3KvNUwNoMnUyZ4rDDIObJRHyEfut9RrxkRTuarKfnPcXjpKbLd0Y
CEuN4zSgcCcZKLRFM/53SDOkd123hMR2D3t5zv90lN04X01g9h3s6lXsw3XwgSIr
WsbnhWbe6GPEjzTsXPTqi8OaMQiAGapBj+oI8erhbctyub9h39PifFJ4LOL+eY7f
oVPO2Aan1EyjuA6zh5nktmsuQZC442j00rNk3Q9wWhh6ljliSEsSTwiO575j2rer
sBjp6i71Ico9l6yAgTT2TwsgCKWXL/55P/GgP0nw85yJL8aDpZ3GS3k1SoLDXZCT
I9tCT/MuKAezUiDGt91/gxuogvUTOKhf3Afyq4zRsXK1TI9K/9xeyG292H+qJHMK
+A3NFiQz1R71IM/sI/X7dg==
`protect end_protected