`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
CRVGrXj3LNIgA7Z8dvGgacR37c75aQt9423YJL1xAplupVIlSo+VLjTm3puwEqWC
MmkyEdK3y3RoU3ns17dnUSXzlFbq6HAN6JQEssqdV2p9uP0QxaCqD6XNDhalTOmO
HPPHMKrwxrqYJ14GNeAYXkRrHly2Onzeq4FkVwLDw5nGbrSNaaaPkfyvKfT+iCB6
lclm6J1ykJS0lgZ92qe0ZTG40tgazon9Pm586jJVus91/oUX0SlR+lrwQ0eYsTJn
ZouYG5Yxjaihk7Ruls5jIoIPtV/uo0FccskcZkJy+w3ERzjqH4JzF9qACktT9OKy
9bmDKUEj4Rz1xMBW0naOuESxvuc4hf00Wq2PF/Cgl9uYss1KmAJshZ8+wJ4MP6dk
s7D0TwehFHVEApgzvJ9HKihAO1piCAm1leMfmG3LHgVGFb05oZ28M6Lt4nu4T7bi
G4bYqVTAnztGerHxlqecYd5xNOWgkNi8M6h1Bc+DlqX30omy+MLcLb2XB7SOnDDy
4AgIC4EimpTy9IByd0eDift6y4kZUCpOcF3e7Hxpv5g8iGxAZ/BZF4Wp5gerMph1
3l80+Q5XTGVv6Im8rUErAb/n1LSho7cMP3xw0WSRrvxdTYEPhNbZOWWPq7rXFUgd
6W0YkDF12IqZur4Hup4wwo0jqCUEcgStYAPdm9xb+hm/kWP++JUmSeeGDVTEgWwf
SYYD47shjdONfbpImMQ+1KcHL2dREshj9E7jU+OtuF2F/MA12T+ofyAMjHmZq/Yz
tk1cQm9Jtl+t39btkzagf3VAtMEUutelvBkXr5DaCl1fJWl01yZmMntaDRf5F+Tj
NDRxP+8LolzfiiNoLbAxbkD8tknAL1ktAjIIEKijxpNKYw8IVqP0JiIcDl04J03C
hbWA7aGldX4TbBu8g85iiq5+GmEe4UwYydaXpO1YpNFIaSTvGcsviG84Pi1rzNaF
jG/5u4w2YAhAb4FEqxJhYhAnpEv57ryUi29jLLFMPbiUc9x3oHewdFjVkxBt43sz
TmMEmYIdsMjj0mgxxRZGLwloYbB3SwYiHHrwnRVRTZn18+qRJNlROx73CxxbgPYb
gJ4XSpAhcO9kSxgjNBw8QGD8L7aJrG8aviVP/FOJqeFzcjymsd1Ir8o1QxERQUG3
B2RNk9zOzC+gRjqUO8QNDR1di7WeM7jsRq+U2oPmzjPfbGb0emNZYGORfFlI7LuA
Z5MsnX/4GNe7zJFA20DHO/ctiBjoYb8ydp60aadFCU9Wx5LxWFbKZxNiOvDvqFCy
rYQHEVPCVV4zRcLEpNKGJS1h5dGc2GobUHfbefH9xq4P4DbiF6pfip6fMPHqvmlj
FI/QDeL/XT1ZAY2QQYnLe0mk2y82obyENaKPa8WW0osqFYO85RUZbTj1o/R/UOeX
kGkn67VsUZ4BGH29xarq5uns5021K7VPTpe2w6oD5vED6ODVARd1ct/MeIlzMaGb
umL4NlDqmsdR0LkuWOCGDEJ+/uRVSp34HeoFHG//y3jh6+Jk5CRS7MZYQelBlTVz
stbh7GJe0rxQsycn8iGlC3rjD2gTZNISl2h6MV4BXwYKEHxGy5wL5f0v3rj5f6LB
AlofRByVBMRlgdK6J4wjnpu4OLETSRGcZKNF8kcoOluJMmPkR1tmp+t5X1KaNCH7
FzZ2XHZBNvfDOudfcISgGTdx0YGNICpmlxJ29mC5xCL3oPYQYDFy5cbJZ8MMDLAY
tYZiSvRLPlRq3T+2TwybX+cJrqrKAtKByMEGnfvf2xW1TiuSaEQItnKO/+Lxf+m2
baptIQX6JXIS9lptfDbrbsuN7r509YQSpXtegePz+kOEOvOQz72bfr4PHs/p6Hjm
ohNix4ytT0i3SW1OtrwcvT7S9wcWrnt4ExsS+hXYbQNvjblfHa/VomEQOn3wXFEV
yRvx8ooB8u+tRLY8kWNmigXeUFlgPGK8YfraI+R9tMpZUbnQ2zq42TQY0pQ77/31
YOb1w9a4ra5f8OwN4RNtTBDuITUS8DkGV8i0uwJj/04NA/YHQvwF97BexE4owS+y
yE9AVqzOa10fv0k7IQlt8MGvOIfMyqjWGk9KC8fMh4vvw3gkMO66BxoAalbEISEz
QpZvitcH/cDMzrxRuFvzks0o0v6SIFrBL4C6II3XMUm9j2WV1Vdt8GCkqzTq4fM7
f3Tb3E6gGZ0a7LL2i6MoL6o9C4SzZtXfiGLXL49LsL9jFdhrYQSJIpnYwvPAr8u8
MqWd8hPEhmAxiyeItq+tU6SIoqLjD0vCjfVzSYESVIs9YudS5CMGa5ZIhyPQXjky
v8fvlw5D532GbkL+4U2jYSn6jQ1UA2h5zv8VfYuKc67/5o3toJjjKyuSCZCdNeCs
za3OPnUpOXx+GJ6VfSTxrZS1nn63RMMEtdGo8ztSBkjEBlY8ICVfUJF5jkGcQPIm
1x8IjWLU+ITSvlnTUlFC3kOsDE7Vx3wjya4HCQ2jFs/+tZwA5cZ4y+tykCmGB/6O
2WY5DgYx6v1zDMtQ05aqfd6FRFPGkX3h7AgO6dOyCF7ckGohsA7+pA5Tf+v6rMrQ
Ix3naszSNyc/sJ58vydsTuMse+G0OwcuiIEsLspVRrfGa+GwNI9BKF1+JSWAXUj/
wOI3TE5ku6RIua//0j38LOy2D8fIfNsXgFCSMRKRNh/aPbRyzdN0g0eifkMzv7SV
KXf3eh8yF/NJP77vdkZj9Znjdn6BudO0NaNy8j7KbE90eWJroVYjw37ytaDGtw00
j5281ZqbMv/s8+ffYYuWZWLpq5+wdTFB9iGH150nwr5z6bFTWU+gZUTXHBh2MfKZ
ulpjGFpRTdIQ+vf8xHJ49+aSVtwP1wj5NaVMvQ+bhf8Rscek973XkRg4NbNZ8FX2
Zv1Jsas7pDj/MU45YbA/tyJ6XmdT8ztkUUUqrnAulxUKO59AT+zHPImW6xiyj7rQ
r/PP4Slaj4f2nQNLCdYEbc5pb61rSf0Gu0Si2hI4Ikum6yltekiJzR2AtoxxPj91
yTiDFda6fpKcG+d37aOs5T7kLcUGzzVCwHvnp3Ic+92YhC9paryjE8zcSm7IpiGh
TXVTa9R9/DUQGTSn9l/JQuWtctnDjjft1G0e0YFCvs5++zDhyaEY9OqTXT39u2gO
/Cu8zdboGvhb3EdVbHdhFiHCf9eDb2dNWPdjXB12o/TSmG5haOHFUbxAMLOVCKhs
NS36JGT3iRcO3vA8PevPTXdHTgRj9r0o+WVE7mXRQalnTPARXnbG/+Md53rUk5xW
oPtxlfiicvw2BTkldLH4ssVZE6/hEaZ9Kj61KNxCl7Oiy/Av0xbwi9+/TWo81OR5
IONZSdcFuDvvRe+CjocJ2jjtwEJcXvtpiANvTlpyNuAag2Zlo45PsVL1z6zRm08D
n5YPoeyHnTmvbwBPlKicOwzydZhTB8edIjElax4uPzWSUMdbmSh9y6NoTqc5EEil
1u5h1Y7ACFA4DXpiXVCMJbSP4OTugFVuveinnWz5KBrjViwI9+VeAalWKyHctgqk
I8nHBcftkpUsMRIMQB3cO9s3NJIWEsgoukI8j4VK8veXnMK9nnWN2PwhCpdDcAah
ee6vAS14fQNoDo5e1rATmJX5bcnBRI3Tk5LZJG18PFDG47hi7LUdhSXz2OhjUU4+
kW+H+TYYSP4R7VBxhGBxXSI7U4iHSVGR01lRlwnbaAUdd+TEMEeWLRWrYitKg7o6
tNTEREs7wnKO5o+tGlB19rzEvNYXsvtzA/eksk76VH7q5oxaD54rj+/ZlEnHM+bv
V6T14luyQDcPQeRt9uLfiPCbad+zP3oLDK48AaZXakPFHjOC+p2/T+X6yedtyJpM
3H5UlNjuHK7CQiVu/1rCXdaNjv2bh0i9QEpg0V7dCoCBlZiNB+R39MW+Sm7xpvWz
Kfgp5l/BGWFyryyvzi3HIWjyAHCCEa3EXGnOwMWNJznVLiKFQv4CkS6vh3xl/JvX
XmGe4Svowi9/inK4YJhyGCxpNGKraHyf3WWw3VMXrhGu+8usLSsjRHhk3XI/yDBV
5wjvfoUZ2HWkWSqQ0uNoRq5ntaqdGq0yMYrKIUSEXZ6m8/syGfuAuBHpILPYjCE5
UYnAQEjwZmTUZNNuqc6TBofuLSY/Q4qSmwBa0ODYC6lf7nzeu1evN1k4JGlNYvG1
z9wAvHDaD7mHO/ivUQeNWU2orqi2ksARrkppLnvDxSqkJJNrxd9fjXDt09/4dLZS
YcPFBO5byVk6CNvDkD71gfITt3Vnv1O/ZzqCkpGYEMtJ3rHQJ6lUA3mys9Uvmj90
m3Mu3GlNGfuvbjuzb210r+9JwjdfPI2WTV4lUcnDzIDVrLk01gg6dgeL4POPho8x
P+85zb1k06owUUoiOIY1rmMfmIOn620Hq9QLkSJgkDi1kxqNsISa4Mi8i56TmBQg
W9RjEwwHO9ZmpHJpT2VTkw36V3qZhrhBb/rJqvx+OgMwvkXfRfWpOIxv438MiuCJ
JVee5AD3JqSUeyklCLjM2TfjjKro5h4lsggmijq47B8tZI0m1ManmelLBlZnW5o4
Ny1aqqqLEHkti0AiaMIdaAUXfV1d+qCvtn3X8ii9GdJj/TFDhvnLfRPMPR98QDDM
gkaf5PNFhyJaqnT59gyj3NDGa8501vuUrRbdwmJ/T1Yqa5d+1eDeG97ReszozGq/
4tDpMjcEjToGKAJwtVlBv/aciZ1WAWOzOpiGmFhVV2k1Q1mRpT3eY6CBoA3jmtCj
uW3m0s2+oR9GXUqgBAq0UsVOe+mUI0vgU3lC9U3v8uETnEK9qWFV36uM7MXVEt7p
SWTfCV2zW32cV/pArKqb2K0culCfGAmji8xuRbFPhGSzjMR7rxuSld26r9uBv4KQ
yKt4iUoGYFYeyHltE43ZYUmrJCxL+HUXpxP8C8YBTQij/buzQv5tVRoRcsKLc5tg
Yv1AlDxkgbQZ7Gj4+hfjYVZUwcaeNanEphAF7H68BMLm5aZzMw4eCcbmYORzJuG0
VpNW/KaMvzwaG/xN4B4h4SrL6uJH5F+vvRpm5CewBzZNv1lIdIGWIr+gzZteioXm
4M+l06HsZLfORiTkoobCsBWuuxC7fBoSap77V+E+MG2zhuei7qd7yQplMWEhwa9C
VpD7p81uox68AyCgHwi7WredJI6SgxGP5CeyyiNqzRMT396gOASbEvS8+40kxiDW
ijdDc3T3gINiiU29w+hDTwGTxMSoaorpQSnOiaAwnoy074pi0xDOvEz97+xPfkBQ
0TbBWg+3sq956NTggXCZTDTj0T4A73Kx2NMLxfIbmHhIDXb7azqeOkVarxukuMae
jEaupDeA8h5DN0PJLlg+z8OWnYeiehsdc+cjRn/JtxsMImQXYikVjexAEAg/jfj8
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
+N7VAUwNNLS98R8HB/Ki85zMR3ePj9mNsNuXsy3aAP5ME/EnDdFqLtbvIHdsq2HD
ZVaO9RBQy41kBPiSfNjv67WtH2iVo06UsGkUpjY+p6zhmy0lVOztZ0u2WBCUsEzp
KjYbTHOgT3cvWVjZbS+iStJKK2fU8taEp+E1xRzRkDCrQGwle3xtbteLJ1G7aOC/
L5zPM4dxoG3LzRodSg7Ta0CIOSbyAPuBN5gZOZnPzT9TDMxDOpJvnq8m32ZXuOzu
gD78pzMk9U0Cdy0yRgdN2MGIrj9PIx/Fl98nsrqHpxTLPw8Kaq4lzC5Mz02bgk9s
pCgLglJhRhQslYmZuB3+O7AtT65d/PTZJjvvq2b3psRz0SGvtYq8S8W21oTA1eYN
38gCeaML/WNG4tmoVsMMcmxG0jTaDpPAO6a7b9wa32c3LnMPruVkJ8tD2BA16LB8
M6T0egAAz1uUTxTcp39pKbnLBMGs2DmdRrAd7p57TImFEA+k/aO0MJKiNkkPjFej
WxxK1CpjiRbvbs585pWC89lGbHIPFJrgv3p3NwSG0VsEkvp8S6V71pFaZHFi6N4B
BCvoIPXtv2jjVEH1B1HN4AcGS4LEUPvWlZe3Jaaus5qim5tjqob3rtXsifW1/DBo
NBrZ1YOCXNTScfa5O0GfaM4X5YQoPSqVkFb6MccUgeFP2xMYWpqtClymedTknnqZ
DU1IVKys/8k5rokkBCyV/ee+Tz2RBjSybkmKwIfq3Gsa9HK/L93cA6zv3FJWCOqc
8Y1FQDu+bkAlYlq8VEhNtxlHXfOYvWdHfmDoT8wiBnyNzZFmNAisnTLW276NHfvi
mgwSPRIf+hcHGF4U3reMmkCYddMG1vSCNscqgJnNV5AlTM09NBJrL0BeAcfHliGf
dGznqKgOEmCcXJaQq845E/SlYdqCWAEWTtOryWwUrGcOAw9pBICXKqTpbvGRsSVI
at6c4IT1ctydGIv2oLTHPC6KTxb7TqUC/m+Ws/UdT11R0fJ5m4gms9ctDRRHI0tX
fcUXa/14VzGiO7dmw6HWiLc75XHKpb49Ndx7o7v5uHD3xokQcxfCaxrJVfFMI9Ts
/nzf1vOXOx7ts8FH4XjQgGP+zaMjAzGcThBvGIovOGSLERXWMCwTGyu77BkCCCWV
BUIVGuwOTGnp8mcXzh6xWDiu2yVZiw1PHmwdNyiFeG7mLSFDDW8wC0YLVQ/0DjTR
tBkTgn4FJLHBduNZFOq5y+gVfkZf80qUR7SdfoD8pAg97hq3Q+rdT4QWZsdNWKfF
BEUjxt0G5/JDXhCLdDbRBHFkmiKGTkqt9yH0vKAvEf9i67peXcU8ucvcv4NtN49k
Y0nHtuBp250EzaNvNE/7IuMlWskisXONA0jSytDcM1KmemNSjfInOfyWB0+DXK8G
B1WKcJFblUSKtZafo1bwIMUSuuqeDHw6CaN+DPRKoXa1nbVOocoquAKgfS5VVudN
vGF1nu2R4z8pRDo5YEgxHhNff3zCbiGNUeF0IiAPBBM0+3EtT+kCSfN3TS76pgJ7
QWhfC+YslKz1+uYLONmV03mRzbsp2W/H1MgM/yyCFrugYzYpv98flW0bPa0QFffw
6sVlC0f+gOdL55CLw1d5vNjOJJ1vkQesAgrVlskg0l95INz9aMHQeLdFqrKp0CzE
BXerMRKCvnGec31CdL1H4DGKpbo0omJ27sdP58fFpGdguBT427TjpzOMGSJB4SWN
BtLwYExF/zDcX1SgEh4hsG+qBdPCv4ASAyWc82oEegqCg8JHgbegXYW6n3HKgqFg
H/7uHsuYyU9VA5MmVvEP9arcmX7+sjXkXpIAu754TUF4kKVD6HSJFHfyK/3M7MAU
RUO8wbtYpmyIchVG9bW2Eykc6gbK0Zwam/4Jv+BiglbM7VZC1Kl628evolQTTH7M
PwPC6q4It/m2E2YMUiJ2CTpI1vr/MLoizetLZFcCILF0fXPMQy1kYKW/xafuc1Bk
XCrv/O26ZNTorSo5nWOFuh3xqDeOGRs5+joPP1uF0b4IwC8PkEhddyAkZ39zk++a
hnI7WUbSEUcszI+8vi/ueifog4I11TgmcCgvHUzNHAyFo10csLdQtIQE4F6F8TJv
EzwR1iD6NoTZrvJu/b+JIVgh1bto7b6AGLqW1Ow1a4WBCEU0MC8jV+EBboZm4t5k
4SNfZHwq90OfQz8T/5yNXMp38pewgEehFnAI0uvwXyfvVvPWCTwpXZWxcEOjKKm2
bWE1Z+xwK+Xx8GNa9Am981bXVixUVJi760bXON4qlqNlXhmvS+ToZboI/eJ2dq0o
nGeOmZZnAwmleVXTm96eAxlr/6TyfM5WBePYtIzog9A9atY1QUDTRvo5nEjjD1eh
eT+U0+8iDRjbaTusQ0d4EvDJzxTb/h+lQIq/2IkLjlfg9emJDVl+g3iO/fSXiDlJ
DK6tIkjfhxYbJhaTQ70WX9RLL2y3UImlYFRKXFER3QUWma8egHWD0UUyqDLriDsI
kNsYcDSKPEDkzdrBQ8/9lxngZZmQSIkzVCdxb1F9V3MNyF+6WdMyIut3mOelqZ71
OBhnKEwI8yCD2MC5mz2GVtXSPNcLeQkFt8y3JrLGATDjRbS0TNha02F4Xr1qbGqy
6rc9z3cz2tvZvTEomIyPqGHrCK7oMyXafFBc6GM/qGTr2Hvark3pCag280Vu2mdj
MPU6a4AI27fhrIqcJl8w1O5PAX1pDfxWK+VsTpJzdmJXk4Oa39AD+iGHjFd9gY+O
KyE7YeS8sy0/qsP/2AEaxdJML/TqhCGb2pZ+JL59S+249TTGeomjSfnEd9L89clu
ZvFB+eDt07/ovg0iIOcf7j5vNcn0RT7vovYi+QZ2vgHs89xTvySAlkRZ3AzEq20I
uC2msEEowH13moS5AcsFE9MiPpke7U4lL5C20PbSX6VNGqs6mvZmQJ2wc3BcKuxp
Lb3bf0inrlX6F/i8kg/QwVgZ2eFtFyP7Kk25fJ7EDdD4w1Rn2egv8aeN7nJHJRqv
EruOWHhj9LfjCVTN3+Jrw3s4VQ9kP/fJ24uvVu+GEKSN+pvrZKE7HRTE5WYlyFa8
Np5Dg/6CtDy157+cMuVwmmROAn3hEzqWymn97sj8jxBAP+ujMGM+ZSq3qGuu/zzI
2HaUiFFq6gl0pZZ04JZB9H1/gA4iRXoYSabn6RRhP5W1fyqx3DhiFIzCy6VPyTzp
ffpmTz55UnaISjV788Y2Fu8+rCWsl396Di3RTnvi/9Rz/msfb0nHFeyPq3m3XO9y
QSxE0yuKNJ/Pqifh9dpVrUCqAcavdQOy1kEbpK5CzmSTjC/1jVNys96W6m5g1LT8
WzOPwQrQ1ZrsckvIKnuDKaQ4LjVHiutbAk8FX/kEH7oN/mIPG4b637+bGiAWEK0D
kFErbYezIY2MwAX6PSPpvYAduCb3VV/VEHo+GRyOTmtUoiXilkO7SZlzhNxV6DPY
B2/uqMFinQ9sExYg/twVsqBcat2twxOxJQDFO2F942ArYRd+Q2i2Ky8j2PaIfMe2
uzoSj8Mg03fcUCMRHRbZWDZwlB+JC9+wlvFmc/D/UlcErKd/HRv+c9CgFpIhQnKv
jDAzxoRHLjlMlrRt+hHiBPNLKCcqVPkZxPTbp3G0swfbhwD7k4p29I34XHsLW/dl
Q40tcZ87bf3pyNG60NVenrv+Gup0s/6/AQC7l8ZFWnUWwrgz8QZnzCubuX56LySh
d2jIDofGn6aEdh/LzBv7eMXcRChHYKed3/W22WXiJvZJJiQAjDhjKGSG1SZNSy4f
WzwXCsxElbI1TXg+qfH/fdWoeR8pAV+X7c/4gghbyvI7G6zk/0v4SahmWbRDWc+g
ldRZW0RNHm7wirbGHUskAW/eqHmZTggHD7mLn7xZ34xFEp8R2zTr38oPlP7Y+Elk
yf2CxhCDqkgM9Y9TLS8mUj7pYm6r/QJXe6mD7dxYh+kvSndCLQNlJQI3AoD+C34f
4Mvn7AEr6AON2EBxRJjf16EBfOamUlw3d/grZkr0CmptcIM5JcC2sNsqkAhuMs7f
HTHr5vgQ4U8bGRVJwzF5wPeE/xyPf6PCllgm4IlYsDCPOHgInLNH9xtMJ/VTVIhx
mAKohqv9yVT4N25k3jkyYgWAyZ1RAoT+E55Gx43PQzazUqdA/HmAbVOAywesxMaS
5HZu1kWDtusZUAoQtydoKAU68pALo3C7DF6djoi+2JYft75rmx6O9BJCXjxqWtXj
isV0t+9e1j7NsRINRfrKSudDol8xO/5kDWaxB4e8w649zz0ACG+yBNbnQ5haVvnx
6kmQATfcBT+tKlUKpFWBBBYayhlU0LqQpBx+2t8AJXwJme1f1M4CkKV2eIWSDjQA
PVPwdC2Eb6Z+yBuO9kI6RxInpF0lNnQ8ZfTLZFLhPU6wxRGWfRjXFZFockVMMChc
1NMLFceHLrjTEZLMddxQBDd6l2pZzyjzm1SnsVjtCxFjfzJl2dDOdDhNymeSPbfS
sySArenyinNeOyWmOCSzohZ4AuWY4wyy/n4UO4sjBjl4bLq1q2GNl+EcOPH4qk5I
C3/jwdMqHUefnR2ea8Pi2nTQ6B50b2PjlogY2gb105+D+r1DpbCCeoMVXWuWtYi7
+c14BkGaFE/ktBbLp3I+AQ7JQBJlgyLQqi0OeKELE0zwKForPNGR/03y/UuC1wjU
sHJc0+oRvp6A3GOhTttMePOc7QHSNndQEzKUT3y7i0b5/JBv2b0if13GWBaurUSW
W4018zU8zkWKZi4W8sEALOT/vAdACdFQbZWJUxiZWPsZfwQ+f+FwRm3wPo6Eg+QY
UroGVgDUGivYRWU1D1aWhuZw49FRXFDLT20a76JlyD+Rbgj+h8Wtj0QBOL+AWyxw
z3GTa8e9zc9aA4lApZ2FuBnCDx2D5vjWU3ESCKbl4am0iManmS4fVJ6ZP9ycIHoY
I8jk/AolNHxkjyEqvqIsE26zj9pj487yq5+wMbypcDKJ7VzzG3WaVp8d4n6vbqhX
x9DMDmDhZBOFFNVFWmVrcLRsziw5cH9IJasmSO0fD8PHEA9ThGN/7xvLrNMy81wJ
2egORYhuzhbE6yJ6Js9NcP3vREmI1M3/LFfVitzvalOwgu6F6IvTRROugeEuTsbs
Lgngu04eS8Zul5/zLCfjj+PYXpqTpH72FGXklQIAQwR3VH5T15BMdLASd3TCsoER
sPtd+QyAiLK71DX6B25nmKztKjnY7EkmblRT4Z6etzkcu5AZYe+5XxjKacf/VJiZ
QjyVy1dAcwh7Aq/b8V6rGtR4GtMvhK8Y/NYgkVtfUtNVk7CcU80jU5xAz7a/AFD1
iIFWQyX0IZyg5kbxdLOp/oauENu6paMiptdSqaXgV8cfuQE/hSvvZUvFx7RxyvWB
>>>>>>> main
`protect end_protected