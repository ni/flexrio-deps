`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
qPJokL5dgHaoxHhpf4hHtoBJVA0/nU3sQXlTmFUOcN7PoXIv1DKxaYdieMCREjax
8RMuAGktyrd3OKCIDCgMsh9FI9uSSs1+A2lfUbpA4AORSM3A7bw8Bwg5W6PtZirK
s1KvCOSob+mPo+H2S2C8K1fY/s9fm/514qsOsqLUXjFtH4aawAn7qxrI3qyC2b/X
f+axWrRX5Icx8JtwDooWyGFUPNzZUwWWIMaLTCk/sH5RYUI+Y9IZ8zFHoRRhcM2C
tPjJO4xIEJtkZLVLsoWsTI6J/V4Ae+AXrCtBZsE3XaTiSReipXvxRU0XZCM+nw8X
TMf/K+qvByaFbQeAJcE/1V0yiOKF8WSXpZaifTgvELhiIHrCli8m8ksNRsxTfm3/
uWdfC9GSabXJxwWxAXNCTfoSqEqxDDFWot+FPJlrcXQd8MwUPIT0emFU7hcWslJq
UhiMAM0+P+OklObHb3GMex7aU7MukRBINW7PpRGZHP6zGWvlm223eFgrYUAceCaW
WdHKEB/XKvo7ythLSXBFLyjWcbsJ9ekI+zmSHN+EuSPo5NBOYsNpzOKDHRJLc1w0
y+XyFgIUeGoCri5IK3+JxhtSQBMNbcZmM+Z05vjVsEDIQCbsqkW0IriE+tdFAHYg
hmzgxI6EZQRGzzQZnzGQ0Jev2URZj5a4Ay6iLX6gZa5XDewrQbxgUcvDZWlsWwGb
wUjCaf/TJLznNXfhDWt8IDAvWx23N1Nd9xeHaXYtLRgd9/oKC7w5vEAjkLnmsD8I
VmbZzbXlmnt1f/FMVLq2l6OThYyUZt+StplpkdnhVg8P9jBLUUH128c4D78us96R
UOTrd5/rRWdo2mhQAaPaumqQOPaqOLNS4VCh0iJYo0QzKmRu5JvM0c9Jh5CcAsfC
wkGI/RiwezQJhIGFSOf7IM+9AINUSXHNjJTXmTxepvEeVKplCVNWELoTLkoa4L8F
62jcun98yM6/bhKM1JGj1Jb2RqtEV4hbIjAqMlU70pizyWrl6asdQ7t5H3nq8e2+
tpg/Qtue9Lsl3stx+82AbXJuRKH+I90l9vj/xL6DHy1dUPF/MXzkBnsI7VR2oQsw
vfnjoq618GujUwkAEVPKAn24oALpmO/PgWX1mNCTCGEJWWcI1VyNuEFTBhlfxbRS
6bG+HvjBaod+pytiBtOgIDSsW12bdj5qi1GuD7/SjNahpMGmDyFKrUa2wbFEx1/s
hixbh3eZkwbD0uhi3TN4LcDYRUJt1CWFGuXskCGT1b805o+DTd3QrULGbbr6wcX/
tNVkPOtBc+qMkIBjvTrsYFkcN65roUDaxSauL1eZ3N4NkUxYebXTdAtUn3kyQU94
MsCwr2GHGh+x3annwcPNCt8xxoTuepF0Xp5eYdVt/kgsTE83LQGS6hly8PAo8qmt
KoSN0njLrnRjQVFUO6ktCAYjsLtkYjnGQt15ox40CtQt8bcdDAR7rhM6nzETh4HY
KUEt4t3Q/MZ2AeMA5icbuYiu74sGxy3Fv8aFuNuNdBId0Ni3Zapa4EahUnY2i7TR
GlKM44VohcSXKfsjDjbPRCMGOU7wTA+wHuE4CLDHMqMun+fh16h4l4Id3JxwmWAA
K1PX5RUxo41vDmX9fqSXBT/KcpaTJ5D1zG8ncI4DQm1LljEyPzsdJSgp73SJhhjF
9kg+ZL8fGAAVmCM145dVq6XFEU3De+kfnRzpWgnbhL7laTYy0o3PlASKQszlxcJY
Uim+H3Y6EFSSwrZoNKvbAAnBPuLg9C+r/85PJQC8kWzki6H8D8q1nMH50nF/ZibS
GJWn14mVJG8qvAuRoIcqLTpNi6A70NOSLpv3g7BUfY5QnsbDneD6uXihrKqzM692
6G8Le7o7bqsamLHrrGzPc86XvY/+hvzHumGvRTm71VMPWJ15HpefI2g3GVA3bOK5
FiKJBntkfScjDxsqqd+cetXQbQ5uTjB/vyf0CpMXIDfDeQZpbha20xJF5NgHFlI4
bjTkVfUc9ukg958FF5WKjX0TlO1ofaCvk/La5bAcj0x5Gdzi3WzJBmiAZlZZ9blU
qkxn3REQ/6E1RTJrCd7ARcuVdpIRnGv5owbw30gFqmK4fLxoNTTF7GQv9A01l4nf
iLHhtVtjaLEAhIMqVo8P6evLDI1UkQgPMMfSzM2xcLHjapkBwtnCNnmHO2sXWWYG
LVWT1wBqTn2HFgsq8k8qVwlbRw7x6cj8RncV3rEj8EV11HMLlI8SHd9o33vGrIcq
iyPKU/91CzSwCBY9YSnxjt7vdoz408oPbe8pwjXW7YqqWUoEUjojJFq//DPNlX4K
KfiDghq3mU57s9xXtgmd+N/NiNWl6BM2gQMjD8uKWLXu2sH8LIoHMMGJJAPaWgf2
iNaBPSwYsWA+t1Wvk94I48oSeeYn4ujkFnlYVl/tL+DgkX47IIEBwZMqG/qTXh2L
PWMfRPvqU/rs4Sk8XWWg7o203A7i/yPjgpBl6EzmjA0U0ReItakj1aOegW+JxLvP
pXUpzn1lmCU6IZffE/jhAC69SD43T4v2hiF4e228iEmtNJ1C0S2QQckAaFcwsakt
Th8GCIs5h/miqGGVoyh/mF/+ejlEodbtqPtnLD5Zcooja/lcWxUd/xvBf8ZvWAGg
fGD8MZ1UoNb785WM6W83+Kw7VeIkVs7bOhB0rEUvy0pdz0PaRyMRTIYSGAHI5Qe7
kCKrV4HMgvw44z5AJ9lS9Lf8llTvnBG71AVcgUqMbgGWOm7Thm1kn/SL+vRYQcyE
cQW3hxHMsD9rXpq3HT+y8ivcsZ288sTrRSgBmXr/15jlCWxO9o2JoD1GkyMivYca
At9lo8qG2W4LBSCdhzgwGhKWabrlX6n6mANrG4NgHhR5pN88WebfspKk8WraKNrD
FMUQrPE+BhFxa4R0TINpmHu9dKxkDtvvr6TpDav6bY0kN/USep9/DdRhVKy/RCLn
ecZPx1L/Mle7TTIc+4JpCANcpcA3mL4nxBgLeyN811REdl0Iucc/jnoCrhiI4pmA
+S/SzTzst8rJ+XGAJCCjsaZ1A8/o60xQg/i8ZX5A7/F5/Vu3ivil3oPfz12OIjxo
2GyT9RS2zgSADrLFUzkR21JbZLrkhmiKszY8yN/cfqJkdGtAbBNo3JN48e6VAl/Y
VC3S5WY8BDqEEu1Pe9ZUNjNydGn1yRLgyVgqX8TFcYbEYv0+ctQ9uZPfBpwTATsb
5mrtYRAj+5PgNbdVItaHtYJIt6cQvlGjKEzjLAkYTHH8G8Sbr6+6W1RJkUTUc3AY
wx3MXyh/47F4WNBEin1d3HQ14E2B4DNvUHHuvZVDH+vCH7NxCMyJxDJOQnn8F3Mk
U01ryHO5Gy/PWbPgiSJnyus7I4EEoPIC2dCSBYje/zOwdPSQSgKzMMbATzidaMbU
gHeyRJMn6D9qRXVIGDN0QvtTVqZgCQGk0h1P4N4ia1WnAzxv9h1wOPbzBnSrIOCB
ZC7xQl64Fkj0G5tBeRJ2DWHFGFTBtWdL7+8M64m89joa2CFwKom+mYicHdaGwMqN
BPzXMp0nPeDHlKKAq8AGySkBvIFD3N+OoH6e2dOEnowdd2D444FiBYUOj10fur5Q
msuoAHAD1lB1lbzq4DeUuTeOc5pbGf+6qHlTtqC9goJYKR73jwxVi1nvPy08K0Yd
BrdVSN0CKUxCSwY4xAVYUaDITTccn213SFDf9zbqErrYV/HMWJojuxwyPaCZMH4O
XlHS321WLQfKS78fTr6KUjuDVB1QXWrK886vA6LdOEnsUpZvUwXlhMbJDhow/YaD
Vzo4xLi/aZ2BXftsrnNFXo7IZcfJQkxKjTgxV+nRC2LPXym+Ek+5KnKRsdB+fAbi
+ae6cRQooNQ95kUSIdWskEHvh/zHWvMUKEbwK2ZnWTXXEk9cv3/BYXHjV02kv1Rk
mUanK7WeD7E2wGha1XWYhgQLB/JSDMPgONYNBeTuXZpttVCSRCQD0WFnuOsmbiuv
MQopygnRKV19BJH3ekdxzNeqxI0UJnnZ5U44d5Pt0m3cr9hpB3r+Enjdr71pypDb
Qf+758/MxHwe3FWGv92H6e5sk3nHrQ3VqVnLjswCUvWZMrEh1i6EdktqBS9F69XL
amZ8yuPgAHb8CcDTbJq83szf0FdsB/W5ImMua7sommQYKvCsyzIPI1UMtkSt4Kdc
ZES1qcGuhumiciqjSeNJ/mHy2bWz82TrSxAtLXKDXL4B8CW7AQBMqCpoqS/FEouo
zSpsZDySX4pir3PUJZQTcUV1nydfgxgO4xrZFZDpOyXkknhbm0kYgRkWmFgK3+or
LeF0tZr+sfNROrujCS5SVRw9xWyg6U52/LL4Jk07iVMQwG4HJDpdrx5vCiW6QDqk
HQ2QsrZv8tdKI7wFnnkvwe5TP+Qn6sqqfJtU4x2H0X1ZrxnAA9AJ3wIgYUw4Vn/L
GTTrSYB58/zNGqnOhDUNSLXFk8+7/kbxTNmCPpP3PLo5XiZpufON2bmtV85uE+l9
OJcXwEuHAdREXz6Cjani3izW8D7xQ7HH+zkbnh7tN1Uip+gTjhoI6/GyLjd95x57
St3MH97EiTtms4YlsKaxiWDkZDhirI2C5HghEsl1fKaiNkaIzAJIx4tRnZ84pQm6
ynwtCqz9yMnbhw2Szbw6hmh/z68O2NZPS/KqStBOkLeKHW7VXZPcbRWs9LYpL5Aj
Md3muUIvN8fGWs91g/0ee+k1wgQTrhXRs6mnDuN79ay62X6eDIVQVrxZ6DjliyTP
1nEVRfmyfMianEG2WfTkdoqXw/e+gLtDU7HUExITNFSz2Rmfm2wC6LAMCd8oguPg
t0Aurnls9jL4ub4IyaroK671zd1KpyGO9ItQrjbpPbznKw9BcFzQWLkb+oJisP1h
ZDNsPuhCINdyP+D8+kcNBymAnHbMfaphgMxzTNeE4KjM7wn2SBx1TY12B5DNjsSu
6coHAlb2wxgmWw0PA7sPIAJsBL65VDp7Gk10MaDe/VNNfILztUXZC/4e4JVtrOBV
bfcT7sZj8qyKunVd/P+xE9KUbUo/cXYkJ+dax/PcCcHw+ygWAOU7+qELU2gTkG0u
MKFEIyoe9djs0woqj94kHteLxeLHaiL/Yvep2IiuI6s6bvFmasfXpMJlcWTzcRku
y77i+ce8R8ZeFLB+P2EMoctgieJzzL4u08+5whAaTbmVutWuhrn7M3AjLWkzUEok
ilFBi6VlOiL07vSk0krPTTt659FfxkKXKIcBSL85ww9d4Jk9XdZn+jBkpwFNMhep
1rtNwisP39S6l+KBB8SHEoarDA/HL6KH9N2ruNkU/FJZw+fDnHdMzkId6hFCLCEv
tvphBwVj7CrAmNPogd9jE/Q5HBW92sPc6gvzfFAWwQUQYIeqx9QE/8EXxeUov1/F
Q2QZWU6MNGXRLO6crbxueHnOe5dkCN7+X8XEmmbblevne66vugrpXnkCX5xhadvx
msphNmvVP85LPppqjmjxuoEP0+Q35eagJPxW5s26MNxdkf9xKfyc5l4HzweSaARx
dnTprPsSJr6eBstLOduFYr2VM2mx/gMRbSmxLD9IxQyC24Oph8yoXWZD+CpZlq7p
HDDSdiF9k3Wf9sFiU7hVW8IaLc1wVIuwniSq/Wij/QaxXf0pVb6sc3tD5r7tLdRC
reNkVCFzUK0aLudNFEX6tzZOeLY5beYk3K/EhgzAmfFww6Mk3GQ3OhDbPN5hN2KZ
gnAJhEkeVsIeZQYWB4thoaXQ0m4t3Y+lWAUiegiMeR8ECEDlgGMET/7XGcpiECPS
FjzJfrl6YWqbDFXKRQTyvcAKf0P+EpgUZazT7MJsRxHaVfl27APa0IFtzXkmWmQA
Sz9l4i/z882/s9o5rSMNvbLsnVywmh4KQY/O1X9bMpbvTDQGWpkEjkzmFkgL8dqh
esKL+SKVJ690xmfYVnYh/BJEyn55jIxmJbAKV1YJYUkM2ZLCoCpdU1n7lKOl9CMA
JMdBk5KLWaUSDmMH4Z3yU3hvo71gAxaPH9euvSmo/vdPT5v90Si3UA8cwhxWB3Yi
CjcqYKTPUlQOCe4SKwb2qNKoCIdCQY/LY85QCL5kQuweBQDB14BWkHzZDvxs0qWE
xAGeUYAeXraEJHKub2PHWdJ4jflcpM9sq1yxdwMjJy99rkCLHBX3zfPHC3lJE+wd
wi5//2LriIlhSPDP6d7xH7LVjcw3CKVFm9mBiXXWB/BmLS18EWj3QsVL9IK8O29s
AT3Y0aTw6dJ7/aUHd4lBbsT43xeVaqL5ULe5o8fpeCIifU/yIeep7tD6qa8ajgOA
Uek/K1FQnQXyFQBw2RKWKv22EnuIuvjhJcKwAuJr/6/ZEDEnqISiDw3f0JeAUGoL
M8fdI5oKmt1cGV30WmudZxePGxt1zF2ex5vTnqmckux6aBHYjgzqQjIhNMvkj4jW
u6/sV5cBXXDjgs9HAf6nzKoABVmlV6kQdT7lVi5b7u2s0oFZLFTtjo0nozfMMdEQ
uFwlzRBqej66lKA1CgyQftSzq1Jqtf7S2UJq1D7SE7kvP1vXnp8CRuvfkeN9bxga
O1x+jJkfq5xJGWdePc17PxiKgOSs7Fvn+q4BMJB+YAgjZzfkvL3Suak1BU+6N5Bk
pCyCiCc0nuEirhXcJeGuxUXyLAP45+W6JUY35xyluNLfI1wT/BfX5xJpOqCH+pXR
bH1zXe5REt2qrLzrECqewidNIqFdOxiLtZ2iGYjYK1R8BrQQavac4zb7y/1dV27V
4AXtX0icfzB00jXWU2gzAlSGJyYkc9He+Umb0/khf/OsM3w18QjpvnBXPjVz//RA
ZiGlGeGbGqgmBL890VvyH2dHIqjadVQ08mz1u6Mdp/wCkCBmQM+cZoLwO5N1Lmdd
G2Cgu+rq856xuG7Q3NDTQpxHW8kgU0sf6x2HV6cXsoz410SrTCFsYV+ghjQnUkNl
ciyvl10dySQ7cZrWxC8LGinGgMyGv+RqZ5KbXMTt6drRUUj3Y1Gunhuug0Sg+fYt
EptqZsxpAC5hHJeJ3B2oCx1EGhb5yhWSAl/3ZthhOma8dJi+fizOWz96Uluof9tv
6a6LyRtq1PdNqGUpWG8KQzH8J19XSL3p8V+OraCXc50cTa+GzTAI5BDUP5fMCwIB
Wzt5VE/+cHIzf1IuVlKSegXPz5MWiaz32ONMppW9qDaIEzLlADD+GHpr8Uzv1lt2
okjdUexThKwUH0V0CnQ2XLj4FhBb+pZCmMvNuLzqZW2lROa8ylSgZWou0LI7BNDE
U6gMY8GLQcKCJCOztfEzaYL8en9ol986LReRkATpm/tCI908XXZhB54ZIISbB7eZ
rQGm+w81rif34OXi8qcMi+VDzK0/vFbHXNmO/OcBIuOXgxuCqU3BLt4vH1K7YDiz
AsrKiHBcj3qVnWwm2A9YA1Q7IADApGYIuWIA+WnmsEFEpiiy09IxG1ndFmjVtWP7
AVHz97r+PAk1T982iZJGE4jwbxXh/OCKgk/2mHEnB/I56CDmKqVTdRuBBbxtthnU
B5Sv/Fnx2ZEEVZYnAd8gQnh7qR79iUdRbdtYecfXhN/itop1gCoLEWFwKwTt5y96
EREHyCRuVADqRFc/ZagEV8Xnos82YJ+BJqcYkl5TjFu8NF6BiDa83osxA8lnD2ue
7wQMKbKRax6tZfMA+w7BIkJpdZxHK06DgSWvwNcwri7ajv3ZOtRSMwNSnTwwBz1I
OldWmEI7Iz2B5VGYVGDBiv0VV23ptR8qKyu89amxRhjTBtzsDuig+OZXsJVgX1yH
2krvcBnZu0QQeMHnaeb4WlMjCVP738JYJKwcPM/BFK09aCXmDkiWiSiQ84DCoHCX
8Xk7Ql7Kgyll2JEp4xYr5QWS/iTBZ+/mzXpR1KA4ZG8fa+pmlppxnBtOM2WHY0lV
dUdUTKVrxJKsyyHxX5vFn9YspSNkNKZivVbjanVD0EQZlUzZpbCK7pS9KYTiCv+4
wJW42jdqFXZCJNmrz2Rq+ShCvtdYC4AevRlj75ykFhH0cmVPj3zJIQ9e09ab2oHm
IjEjwaGv4cf05Kheh/NGXn3at2DxJo3Sf2mPZRYtmzSzZYjE6JSHWAQZHuzb1Ugd
03NGtL3tWplxYgBLiQgrRhzFYmBKFa8aq8N7HMpwL4api6Zx0CIU58VGiaGWTKvc
MFAUhYD85LJvSwyJa8899y+fC8kzvsou5kWZrDAuXEy06RVi4yNF+Jj3Q+GQ+Dpa
pj+xRa7jzvc70HHN52LSFG33vnG0Ymhy1pmkp1x8y7nRmKauEzCIJqyyEEJFlkOe
uE2pZ4op9Pv7dYnHHalDRbZLaFVrG7T/4ctSbL0IFJtDuDRmFB4WLx4/qt7kgBCU
V382fO/d/V+GdbfetirEW143myYUFqfI+vmUgjMwWkLpy/eEZHSLepLCe8mfjvS3
oqZ9ZlMaN17IOw1wjhaE51c52kXY0qaUqWU+DZXPz+gfIPnLY3TsLL3/NEQ6jHg2
B5RgHrCr5FQ9uoRuEP1AaWVXYwkKedtsGuEgPWyxcBMt59LM6YdvEf2cR24rWUtI
wNlcAwBhdTFu7JZtqjTRq6EyUYJDFvTbZc9+WZ72lImZ64BDXXQSbjW+MdOhhFfy
V4/n3SwuEsMPMGlu0xGADYxQAYypKjfDVmCO1HnKYL/2LcPjKF31FxUOu6W4gxOd
lDRt56mQtKml4HVtltEaql+zswKAXdy3Ez52AGfinGD0eExJu/5MzneMWD/782p7
MGrevn0UWM6AIbvR/xjQrk0QChctbXE1Z8ZSvRdzCx7xlgfx4F8mWG6IyTGkPCoC
ECGxdlHeaL1LbHDS9sLkmBuTQzi0MM+cQzSou2zgc95zsaV+92JE7wK8TtJt5rt7
aX8Cfmu8SQ1exjI/+omTNcT3ounMRTqSgJNQmc5K6hdSIdF7w5mC7FCMOSvRTeDr
mHHkwaGyQ/X6GcCHAjXhVJWf+5HcjY+ZMaoNtblmjs/jDKlI9pzGxbBUmWNiLp1R
OUE/DcfqIK0293GdvKg96UJQyolZ493V9k9MJVI+cRC2E9FsiFHDutEt0AmCHEos
0c9aUybNlu10mHg6DEWlUP0B+XUdv7LypuaJa92YUDrfI4EZMYjiS5d2WAEo4PGZ
qUzWYj2avDPi2bHAkkXkUEefkLN6E3EpzhUALlYicDsEfDjXvma0vThL8m9jGGgq
HmxCR7ge/8spNn1Sg8+4dx8x+6BPjqQySPP3w7jwmwFjvwhU+msr1NPotH2Bn5hM
lgLZaMTvx0DlHR9u799fCHXyklS9RcXIi+34N2yTXblNCVdP9cE54Xjf/41YBnup
HgZNKp1tcMzBTM98c83M1X5WgA/WorU1MBHV/laV2/hV1qpp1VqzuKRU+8Or+YIl
ip1K4xka9Rn/nBpzRKvbGnk7S+kA/v26Z3c2M+BB1KS8zDLjPCDP0o4HVeILMtIG
/t4BsSGyzM0ujUsflxQh3Qi+v9FHCJY39qtKfPQMx3tfOW8R4qQugWY2+3weOLXf
NbYGreOUCxyWRx86f2F9uacqQViRVQ6MEtMmm+OjpuHGkDboD676AKqN7jhR4jsn
Ieoc9ayvVSQh/X9Menz3XDw/oNqhkPOfGEutLzh1QVxu5s7msjvkV0YSMsP5NjR/
TbKY36ZVBo9Xwwyz2KnjQ9iwnFh1oJ7Jy6278pm6XX+si1X3+yKP18pz+5mO5eqK
sDjVGgSXRH7K668a0rdCNdIfdIZcvMAmqlRR58wfQEptrWvYCtrworQFx95cEaXL
s8nx8PsWpw6ANH6lZ1l+kmyTQWHN6TQXEcABRS5p55Z8f3B1ncj+cFypNZrTMNIa
el+OICP3XKi0mUQndwfy37ZhAtmtXqQa7xkIwXEeB6aiIKpJJwijRcJNeIH4kqsp
VHaX2tzwToqmbSGF4zxRJerfuK6adpG9MEmGG9gH8QGkpT649v7V0tDNjvit7z1j
cMeP/FCRPbwHhQqrwCYTGvyWHWzIrufj1j1TM7pTmWtzWAk01pzzUB7Oy30vhsiF
ZAZPXUKGDgaCLt7g5mPj6laGS/P541vYwVadp0NbtaxiC1GPeNfDZ9fTxkP3XbR3
xFdMq/eI8je5F5CZ/Snvq1xweqHlSBIwUOzSkPwJCvMImt7sjlx6QKnHkrt9Vp1z
2bYiMZe21JBf4zy2xfQq5FhsXpNAQ6FrAToFyx8QR7km9g0/+v71mbtJ4p9Lu17p
rfWaVABSWtPhHD/Izlwf8SKrvcXlMuAkSCVjOdHSUHT3j4avfId6En2QHZEbhbxI
uNtbgKodc0uPzuYfF/bW7cHi47N9HRUu743je6TA9B3jePd4mitlegkMdw9q2MXT
83px8CmV9Ikh57B86sAofjE/FBu/HlbytxuW4BlKj04Y++cIyhS46nz0S/XJKV04
rU4WVRXzjD3HKpvEYxe+Y2atwxP1MT18nPpNe1KK5dzyGXAPMS21koAjDhjcw69r
tllpvPN3ByaLUorWHo0A6/4gsPkOHE30lu2BONEEBZ/XwA/Vy7qyyEhNjyWAtlAf
K5jEJE0K5zurjJOdd8IgsxbDxxRqBnDD/AoRbi/qq2WlZCj98r2BtqXwYq9cNqJc
JHQcgMSD4u1j2PMzEJsSkVVPkHVNhjH243IR0As30heSDCIBP/lyG5W+jFUMjddJ
SyvJbMpuqijkPuDu5BEzu7kw9KBf6LPN4DdxpwXg8Z/RajWMvpXEJXCII/qW/Idt
dxXTqD28cyeSu+wb0TgEtM8KDIi52cZ1+qxCj/Pg+eo+pOWHXnmERBpoZVdv6DYR
+TQe8hPVrXgWhprA85yhvm5hxTRjJfa7db7aWnr+lYQDI2x2GAN+YtusVpvDqoon
OMOzx1JYzHYFi/X/5G0B5QKcmJjNclPS67iQeRXPd8EJ70SHnVVKfvnqtUqG7Xt5
naas4yO5fSaju8ARNotpve9Ql9OdwQZJQcGIcsIrOCg3zvYtpKAv1N5GSDDGN1ar
NVNJx0Ro+Pdx1o/Gj++zQuMMa2WQ9CjlnpQfb66i9Q6d6SE8SPlWTxfwj37bmNlV
PJf1dQ8eHPFY569mp36eTIscwvA+Qpn3GEtnm9K0CttKfSwU32N3YS4xsn3ikmF3
MvxH7wRelqPyBNqn/lSe4HEKMKkYGSUu5sGS3TamxCzJ2U4BGoXz3VkSw8NiY+cb
Dfln7tvldjDs9RPRDkCXHzAJ7L+EyVgPSskw/NVmmOvlGLzrRVWiHWjq7oAoF76k
5ukDHbuzhyO+j2/2zoEaXUEuJoqtlrdVTx13ratBfi6k+WIuYKUw9M1JNf3lisvU
p1ZM/sHCayw64rKHpOQjxNA/cmvZ3Bu1hkUw75TbKzV+B1ptbla2rYA6v0E0ebWv
fzhqxePPYhOSTVRasNejzGJYaprNQhjQ9R/0LzALzFbsUr+yf1G72n9kkJ58g8zR
bTbKoMP0HbYrxmwJOd1LJeKZG0mCeIOW6zwg8zacCixrkNnEAGMITS6DME7xpRc3
3TAkWE2GEzv259WIDgcMW5MzD3BAji1pwLGzWsf1kUTN3qg2jcnKMYMKYcRAcFeI
/QexFsV3GRGra/lr8KmRrJqNPV1d9nNsen/E/e8MH9odP+cY5nr9uByODg6oAGEU
lSqhVbHF2HX7hQEs/y5Czjg+Ac1Tw/8j2gvP3Dcqdy8JgvKCHFiw9zBVVYPbdKoR
Ajs81nfc19htGvO0RcYKbBkS+EzB0wVX9mejKkcK2M1ogUCa8+n4tWPwC0qG0TGR
2/EYz+UZNmr5K7DtilQ5ZUPwx7EJWCF0Vp/bnH30MpEu8pamv2gHFycGhTWVbSg8
CFAT6D+j0C7o9eaqvx3tYCnxT0FGuiEV4shCJkj1XMYPT2xlAR88XwJ3al6B3bwS
Hnq3wyPC8+BI8IILVW8wwWNMbPgKahjqsvitk6eFMXWoMxN/NfXjSa8B6tDIcE+v
xz4jahIeTvP6k79kar0K0KxShjpf08OhMg+ZYY66B3ednEuM1mxT+N32bLJt+Qv7
+QD5Bg93Tdo4gw+RkaxrIRdU2XlBlV5uYBW1kfvUxfUXJ83f/AYT0c8rS87zkd1G
wnX5gaooVEJUVixLtyplGr4D58knynCUh8hhGI4hYngZVnus0CrOSUVg7g+Ivktu
+U06qyAurM3lCelTtZLcQ9ZB72GdHUnF3vM+B2rgExv2Api2IOarWfRGBMDn/bzU
2xzCQjYB2SPH42wJlFEaxT0kqa9zht0HLT6AmwuYmWvvIz7HKgey5F0uMBzQKtxQ
zLFpZH2lGwZIMgO4rt7gSFlw86cVRYyHhENA/dKpjCuDS5sIbVpt+WuNunWEwF+U
Oym3nDd55kmcsSWtn4ZndlDC9LSYIi7LHFqvdO88D3KswQKuass2ay+2fZ2HKPOM
bOsbcxTba+ujK7KOfwRypuzq1/9ZjXYUpCwtkH1V8ZDH8ZrdUes8JSoVj/rEiHpA
h9Obhr9DoXP8ZMK8a+fayzCvwyU/WZ7/KNAH29WP2aSi5lyT61E2219xsRYHWkU7
UP6cMPeracMO+i3QUmVlOcw+1FlnUXOwNpfiQpteP0wgUsi1nhoRwQjniivBaCDb
pS8aAduYPwWqJmcvUblzHMy5/fvmW/ZY4boS9IGpsg1oPbnqTl25tuC6vNfdcGFr
wlQI+Nphx6UIf3brTYJhrmeanBV7yDqTeNyR3Dua4Z1EWjrx8TtKYoJbsDhi23w9
Pr1gP9OSrYJYhmMamXVYBQEaZI77zssiPITTv3Fcus98sbJkr71CmuwAvLKleFsN
VN+VfH7+gXt0tQCIK/YwsPMOsQ/RiorsUmdzLrRdFzb5PwcixGm/C97DS9RfdHyl
aau1rOLuls405IQ4uyhsZU2vQDFLY9S+Ju/iCVqQ03cp+qcap/Yd3NEwT9rrn5nt
8LzaM945OAE0ZznrcHKaJuZFoh2VHnPyq3CdqL3Fz6Ko8VvNovrmtjdlyw4BKNm4
0WZGJQLulZCDp1E1Bp5TBQpFZoCTOqcPcMgD1kAuWXL5VckRobOGVAWW/8yvgEOC
aeEcjd3vtRFyrZa2ESvjEJhKoaiGCwDniaMXZ5vxbgUkBUmFD4qGoz+GHF5Y+eOd
N4ADQmzRzQHEXf5f7H8+MALtXDDUq+6Ii3KAZaMpIsX0J659U/i5sqwLAaRN5a0V
ZPxAlTmoCbD4L6EHoWw1W+mEvPdGYhDC93C6Cp2Az+3EcHbSmHkuOJV4mup9VyWT
Gf1fp2JpGmhrPRe3ZP3F1lkGJ6GoBQlLKZHhkj+jxQWavAGUo7U1mF3CSxjZhKWP
hZZzQPIW/A7+yJvKoQzjE70eak+oA/JLDoN7cwi0ZgIKAXekIXRbaYKAGcDnv20O
bedxc5a+ACYeiSN1huHB/GCiXGfwLtL4dEKnNDD2yKmP0arIpK9dcLkkSDzlD0zG
DQsuL12H6Kh++EShkmK5/NZH8B62HSQBSnklcA0rNjRmHIoBqPEvGyivdXHfvLdp
wzx+o3nUD7EMjr/XWgeL2TbbmUeHwcSdUEs1X3PX9OaXZGjIt23bv2quz0WcIYbQ
9lDvPDmh46tH4T90FlSQ6AwedfWa5T4k+vCBuB4aWOzHpz6IMJm/xfxwyX/n00OG
eoUXprnLYn2KLhO8iy+mRiALOJ133sR0phVi4K3Okn/zjKh1M0WegWbauwPbrNnT
YLOJJHpFG9UqNABdPYIUsdvCkTrGrUBiti2zAvTXireZZIT3/lhrtEiOzQQ69HA6
CXC3uaVIcreorYHpC/m5NbPVxbLoYJVcL1i8a1C3BrZR3usvaIaGtsoSvHfZKe0G
6hbgQS3+Uo1b4RbT47bpuHGhBXnhesHWjB8CSUgCuTiMfbVXlXDO2FBchFl1jURb
+oNOd7U4LRMxsZoOyuT0Kz8KSRT3/RkTBZBaHOhJcV2B49ZYg7WnYTYUKqe2h11e
4qpbad/YMZjk/n6QGggEpcYzaWDIet+Ci+Dc/LI+HHyGaPd9zbNC7j5Fr+EVSRCg
D89DhCm8Gs0LslzIPwSaVYYaGhi0XQZdryYI4SVr2PfBfyRy0cvgkOPHZyuumgBf
/x4Jw5s6Ng0s7Lvi/RXezMcK7yCjL/xEBdyTTPn9cjeol0XRYgaC4U6rWF2aGNOK
jXR14UIN/UO/GdvO/2gnmN9ASPXAKmMshuoeag+G76RziNShP6I9bl5/sptkVaYa
dmIMo7y8ySlrBSyZ9H2yQ+tQPHQeSos3MMrIc9jXn4Rg9pb1Re7vAGen3JxlGM3a
EQWao67WGv/35ll4QQF344zKnU+O0rwGWExe/pt04UhcUHLHukE3z6g/u+ccCaVb
NPEwhEdTUlrhrp39KRprm/vntGqfBJRgPW/Bg7piPBVqr4PqNrVVygsshWZLIqdm
Znf5P1YDX98ZtFRFKFtH/l7OlrWoALVFD7okPbTBZNeETK8l4pYm1o3UtNRgg40U
HPKox7q51a52IUP3r0wwr/g7UYfMZK2Pxhmv1FtQ8p881x167jcwtLGk9t7YOJ5Y
6zUey3zBYjYq0CZ63AtSMysdlo5yd7Mu/RrWlmRSb4mZTMiGARTdSIBM+c5ht77i
dpjChQbAo8AXWTaMT0vvoYCao6rbk8smoX8OkKo2a9va5SjPdHwjuCroudahJFr0
NnV80Efo0jFZ8cnl1WQbCofeJU0tBnOvb91jdESyUeX0ytoo6W4RRmGU0wkQdKU5
rR6v1V5XHeTKVu/o3vkDtGS2Jk9CisIjssPkWHZ/44agtkH8jCnK5d8iSGXvUuyI
Ntywm9i+0Hjew6PcXj6C+0DuZkqEvxWNBjHmfmRg9h5p8S/yID+fTDPn0fqHd5Gw
rK2ZNvPW7FEG2K8N2lbY9MdR8kaegKrcVkAu7PmayfHnChSqkDSraRzv5/OXpr7T
PumF443mhDITPEPoYvaV1vgnKdb0x1P5HjMZzrPheOHVbHvb8YKgPKnpGC7GKnUO
7vLb6aLikHrCjSE6BbKCFP28wh98pfmXCahIHsSGrZxVWTrRjosu8YiLs08rt+0X
V39ay5SH4EbZgIif5CU0KmPRgFu7t6brJpM1ATdIPahflCaJtTdfJpTiNIajlUQu
WDs3jXbEY0J/FcOk+e4BoLDxajYuaXRZVUn/o4WDif1I1Y2orVaoWLVsaBqb1LXQ
o6OHheSEry/xZ7yjobGyKv8qmzsR0J5t+AqttRt2NDETtm5zslqx0zSdezUJJ7zu
LELiEO/euy2fvGbIRVpnnqOxlnur51QZiSlJEWs7wIwzWOxEbecYgSXUpdzNzMGb
mq0V8JaNq/AmTb7QzDUvmqZvUhz+cLqN/TNHk5zptNlBonwpu/Qm9ay9lalAQHZn
O8P32nZJcWXrKl2Wl9Z+qyJMVqZFFTxypCS1Nnj+EziDhLcg5///Rr5YI+KVE8LD
Vh9AIwZFiXk2BcO/lJjfhEVMpl0uf6OP1bR5XzGWdQojr1vyUdaLDyuavg0LGhjD
s/bjDzhAa+hMkycrSwTQ/H7dsp8WfCVXlWWemXEzv1vuxHLlNnVeMXudXIWXtcG3
6MEpCO8HeowLJYVM5PA9mwpcwqdrB2n/+cq73UY3yxacPPckEkmMSBILEwZDB29t
TwCcegcbFusA2hvienCpN6nxvxYOLU/vOYXwkVUAIyzTYHI+A8WwaOdV/MFu0A2z
3+lbIr0Ofxd2ta9TusqbhOsrBCSVm0cPcZloYcURCzGK8NNaTeuTrB/0QkN0+apt
CbPi8yqRaIEMU1MyVRA9kfdkrzOFRHd3BHd2qVLNPsUFdDn2ijbBubmRkaDE2Ak6
UpkOnQXuPIT4zubulcZVFA+02QvSymyDqBDOLOBlN3Ce9UvkR2fmRsgoshH5moHu
6mpHo7wTvcRDLCa5XpbP0NVSEXiIvgQQlt7uL8eiBJs8Okt3b3KAtMIc56aKp41q
NEqwjQABZn13iNHM/GQXM7s3q6LIDm4Mmuv175KtqdH9Dwmrm7haWcbj3CjqIDOW
/KdvTSxxkHOadeVqcUaOALN4ceOTNFf0YiB5pBD5MZGHHxYpqWdcaiOZDpoXw4uy
uxbfxhYHasgXXtHfBWH/vUDaWUrPFc5QVw+TGHi9dYzUvRbI3a7qiDQLfEnw0eO6
wtnkb7aB102oLHPCkMgszA/AaIZ12CnBo346Fpmg2Y07kZrCztP/3vvvPVFAlHcM
kl6p8GlDE7EGYokhAlLXGLOMH3qQ8usTgz+0BK9a+ZZCTA3pZqxEotbPMpEG5/vF
Hjf3da34p4geer22bGhQCcHPv7c26otMLxO7Wa97s2U40zkNFWgveQjLLp9PUh+3
fSGTJLgh7yEVWQNigUHChPabQnGIyguMs+domRp0+d1/CkGbcwH4VPM9QWgIGW5V
96OlDZvuY2TPjdGkBZixHUmbwLCVLxRZd00LgG/BcC2MsgIHRc5rChbgUQN+mYPr
t0/xlSkgxTWDsgotnYrRIXtzlT0i+VTSoel1NydcGTtEdjq8qEY/OhCHb2F8SPfz
KYpQCeL4m/coe+UPbKV2W+pDwH7PERWu5ebr1zc00r4ytNp3m5cXbl6ut5owUp2R
IcevcbQaEZEOMXErmkoEl4jx7pYDFCfkNklDpLX+MXN0rxCuIYYHqhEuo6zv9yoG
ReZOCE+H77ylzFBfgVL21hhfAdLYjiW14FYb5a8OB0uQuC8IYu/EgLgqaLx8KoUH
tCmbQKZKa7jdXcKabu0caPBTv0wBMYHCIVXKb7luqJIP3HtAMx6gRm87XJmynRwV
5TDuPfn02R5RtyX7I2susbPKcXPr3NPhi9lrHoJwXZA7QlV9vt919JqRLZcycsIQ
Zfj7zYk17vS2YdzyNTUIi36W8qm4DGTZSQ33D2nQDdV3V4l6+rRuGWsJAStBWTY5
lkXzx7t5nQ4QCfNpo2cVVe1pN+OuGPbMe846aOMK1296sXPDR4lDYLHLzoF8zRR8
N6FwR5XDLAnqI5d4oGvMMwzdNsQz4Gy0Urjjj/rGQj9mV++pKUCsv6NE+YYs8l40
+ZDtnPwo95H1ZplsQ7BA/CeGY5yqNTc6hkIj8UnanuR8QaKgFr9OzshMwnBem1JW
I63qS7X9/ryIuI1v9s5VNhiEwGhR0peu+Dy3PzPICfvoW8R6bIIH7fPfHTyh4XHe
aZzxXyT6CGG9booiusWO1pNmzOb7tuHsIMHb1w8h+mQpy9jPw8pIuVIWZTkow2ji
6bAwRTQNuYK3FNkCp0n2f+LuyB6g0soM4zXJYd7UoOMCTWhSjQrg41nD1vWIVRw/
yjrbYnaWHjapidIDnMlbTEflFtm+HoEL/gyo6Q5nalJ3LOp01Jsa71PChU5vaz2W
9/pi/zjJsfAREDoG3AK3NQfHzp0Q3lXKsvSePodQlWpzimgRxazkycmuOWFMxHqw
vg+IV2w5fVQvg8mSY0eq3JXBxDLtCz/WHdinC6fKK6e9ZfSc8gXPg7GJ4n6D9Y3V
5DarlMct1Y+W0H8pNJUfwJO8G6SYHckApPWj5UipdFu/+q+bPaApL9I1lM3vmN0X
Ux5oS8mma960XsAaQOUwbNcIV6dsKOzt/LNhT6pJ5RyR7jHUCtxqRhYq35124/FS
IEKqJzKIPdzChSjf3gjT9mc/KPf36yYm4JKAu61lQhWB1c6t3wI2y3d1KtjEN/Hi
iT8wYprQWI4xmOSsvjqrjhergDTRg8jj7OTdW1qjVng5rWzbJVMDT2mPPcWP86hm
ir0RGcdyV7xhIY5NSXRWws5EYwY2gvAZUAOiT2XLIVQtggAbZO2f1UENfqP9JL4T
a/d7K5EPKvdQS5D0StbbtBe7NqLDuL2JxiureeE0/Os2QmMjS3lF3o8d13RnvHgC
sqIWc1Bua7oWoBFBp1LqNZDW3hcxDU2C6zjiCEkpEALQkNOcLSIAJo5MOeVLWbNd
fCHzHYkz/tGMrdWW1v6MT4RIdzWjj26WdlwynRykv5RsrbnWdOjVMhZlV7dC6NT1
n/U2iMMTnyR8bieGFLhNsHXfQkFoVYKOy5lCa/9LJhnd1O4vFXRtmmNSoh76t6Xy
5s7JO1MUI11+BDEL+TyhbVc08WJH8eD1+hxLdkP7NAeOkptQQU8g/E/l/LDEnU99
3pDvqhgjtuFdx937JbCDxztWzu+Z2l7InLZkvKi65C50UxXbMQ/R/Pl4Dvn7MaTK
wCaoSpJTbscQeg6TjrTwbGEcch0o+LzkpYCZaqOVilWumKhYX8EXQ0oekwjHOlp2
bWTJ2w8NlJmsqxcd/BmcEj2K6GDOuWMDVh49oMbaPU92sInw6dfGoJaKroftxn0C
2WNbGs27ZX+gmsztKGYn8shvYSCc+AcBBNfXVL17SRHLk3TPT7sZweGJD756d/iE
63pX8/fG/w24VyB4hvtzz60XW434AVBPhWBASwtqnu0/Ih5MZJySKMn1Ei//kP6e
89B6+jmxXAp15P5ZdaJfD5txQ37P85pmCZDiKHUsCsRGVW9pCoaq9n+POw2icGhH
pcvWnd6InZsxf5p25b1KoI8LkqFuNcUKQ5Vi9KAQbiLqkb6mhj+gRcVTDXkq4qg1
gDlzzHacu2jKaAPM/OyvIw5XtuEF3HYwtXmxJTKhpeJ/a4M5zUFDMDVQgVtt24n2
uewYQTVoJAt4zzaLxcy9CX4iz7ySye21LPLStMOK+MpWGk8sqB4oZorczzvXurwb
cK9Ijn+7KFfDe7M9Pd5Wrgd5j+R6zLJZGXQ4iuRFgY+R0ToFpdvxUlhgy/NqFkzr
D7pNc4bXuyeygL9XVslRi7rmiDuXp5iRmygFOMP60hKuf5q128bgv7K3xw5HQFAc
4omqH1G+QWhedTULBubs7N9a50poWeKaryeUJoU1kNQ++43VyYeFYeq0zk5cXfsV
HRK4MqgHIpw6cs+o4nD002ugPS+5riQOaQHARNSM/r6gwxpfHxV1g5KSeRriI2HW
3LUKt1shBp/UBPAgnsuQPmQXAzSH3oaxx9T7faHMFBqxYyI7DMC7rTCS26+wvKWg
baGWyVle1D04ckOMKcXVPoIWSB1pKh0cFiqtrAsF2nhWixxwtNRFC29Tv40XwhoA
4MoTnPIdiMFcfpKq8qc9iaVSZly6b+oj41L3Z3W5wVmfxuDr9X+F1a85JUvL5LP/
Y2f8y40fGiAYPxiCXuJNjrBjMbznen9VH4PrAsz+ylGspMgjrBAV5CnUKuzrMrE5
6JtAbV+0v2yN0R2IrvJLAzDihcF+H8TBLkE+g8SNhgOfh4Q4ORbKwudlD7PXuaam
AsLGSMnD4CK6Et4Ev8R2DsWtdQEtXIt+HVWv+LfgI37ziCQEog2Jzal2G2YjuH7r
b137CxmBnjB3AlR9x7THrL4M5z2sJw5krioTCneMzMKIxVhYCC02OEQWW4qpoV3i
OxnOIGfo4mNssYxvVC7eA1pd54jL85dVTuGhnjWXESa8bydNvx+F6G3LBx6dS0EH
CBxWtzamZKJKacIkN9R6rJgBIwES/1S3tiwks21RlRJaPYysKG4pn/Y1xTjSI7bJ
AqoRQp1g+uvqepBjTWzIFO/nzMs8xIH7UVfl/d+aLuDyFKMrcn33gOjgD+hkmtbT
UwXE4Tsss/J7UpuUOTTTV8gthtdY7wpkAUZ9TwEkfEk6s3vffTMBIr3XhGT/wkpa
+F075ofMZ3xB9nJMnz3d3kHgVPkjbws8nyyqdQJucXh3hvNDBNDFGNNtFKA8p7+h
07nq930JDySFf3azTNti53r5vFG2HuC92dH2Rdopo8SGdtNori/aptGshl0AyBKQ
pPDiit8BPkDehVWInFOvEgkfW9okiDrWO3Xw96OEt5w1FDDl9cWKLBKMATqcnwUJ
TTSStmZ69eZrUVtoh4uzpIBWYvLVy33cBxz0gWlgStCT0V5SkPSYqlHf4zQmqPH9
FdSI8OohgeVY8gmxzDq0BmQnmjXs8WcGZc3JSYUqO2ceeQhN+zQ3vOxnauiUgLVB
wfzSOe//OwLqr4QvCiYk19vg5isUkxqfmVXIvAOnInhneJY+YUBDmeqVRZ9VfRnr
PyImjwOfrIuxPMcG7BvwQM2735zhbiL5sUQVPReKAL50aq1CFdMISJJ7dWvd139B
GGouKotD8orrJxd4aucrV7MgmN0ExHWWg5UTLdtMVZBDXeH+MiaeGCcscLQXLojI
NtBSMebuuWAoEYu3QGQw3hSX/m5Ks2tciHioUYngQnoGEhX5f5s4eOKN1oMAwkB/
kiLHZzqpwSNO1WMErcWpP155TxBVYht+v/i0Z7J/Ns5dHlC4fAisZPBu4EYjqPXZ
WUFjTPt9MjbgVV/T2M3t4KQ/rPgSKxzhweaUeYZ0/d/LNa/kDv6Aj6ugNjx9QkWa
pvqRPJL8a4kVRcLb+kPHkWt0jRm6RO7qi3zLA2zwmTeN2xRbNTJmgLfR8f/gZhk6
Z2SXb/Akz5S5++w+AeUTrzIls+EhLha64VTU06TkVmIQ5pkEAB8nujjSx+/G2zXZ
dMX4bhR2l+OHXZCfcrBEw9yVnk5xbdc7gTirke/KFaGQTUAIxyD9Z1lnU71VXHBG
FgUr8elXHiPtqAlpO9Y86poOi6H2LrV+eYlTsl2DXkDe+MnHd2iZJyHtRqLrKsSL
NN8uHnf+cqWQbX/oDrHp0PB2CcvpXfUOH0GmnNayoPrIFGcB2OgSr8qdFFMcyyFW
ygpZkhB58yEDmYAF9DAe1rXmcjK8yMe0y0bufkuhVLD9Lt4Ag1K/FTRRldsRcnAl
VgH+qblgibhDpFnywivjMjq8FFpEqfNFvpeLl0rb4yZCaGGvdg7LOnyUHYm+LWvm
O3dR//4rtnwom1Ztm61Ba/PRQ6t8dgwdXIk+xTL57xGdvKwGxwTlYjCbYAWzhHb6
/rlm/Fm7fNaVBRn9MumdB12H1yBKfXEvApN8h4iyb90xj694Ns9EIXbbxbcgNnt0
+Ly6uJPKzNQhNGWXXVCureMVIEd9PdwXuNghILU5zkCYchWs8W3jyKCTQGk/CArZ
113d5ZaIei3mWsW/Ka/V2GO1RGnv4bIf4TSrZ5DbEGN6iXnKrPnIF1taoqbLYHWR
1NQPSkshfu0cqyZP5Wov7p1b6IXHQb5stC7ADAXtPHoJufNsWeecp/KQlI0l+FJL
ur78e7Eij29R9Y4f30PDjSqXQglk86trCVFs4JBNLENeGJCdPruyaMi4QakpmY2u
tQzRAqxgdcjoALqK/5MHuxaL6+zPMHuJDuHzVIHYpNraZDx33ZzZ92QBvZSbiO7+
1d9ZlPZvIixTsLOtaoq8mzIjyF7mkbhiumlywaqeqGHuiRE3oa4FiQatyiDABzPz
PQUtEZVkpgVqIG73N4kBbo03YKLbBulJpQoIDLH09B1mgRUyy2JxZQ/hJ19TTHSK
D1l1bhNiu65abT1Lnlac9QaGfFkc/nOdTBgD1TyeB2ofIiSSBXug8EQi59H3LJRj
iyZOY99D1y/3hDVGsf37xJdjmpND40KcwSbzL7d1HE6DSwrvv9iUBMgYadlJKdkc
0Md6rNfKCCxZ2mSIMHkOBJutfu3I6F24TLzHbqlUL65xVSEghI9w+PwzZ7C/KFLw
bMRfHgf+jxwFjKQLM82g6Pd5iwjsnvB8c9sV6HIypwaIXvaT+FZvUjbSOXPo8f3a
wfcrhc3LGZDZHC++j2w3GGeMZoY6J7x9CuCUG7CABFeiu7xid3nqi/6q1YJDOyO5
azVZwADNILA0m4fSsbefSO9cDJyIWQab432eiKfYrgua0I8peeEPWx0wih623bKz
1EbLN3sSCHSogkYjZQ8B0oojtWStQErXrvqwx5xJ98dgYorT5deIAY1ezLUFa2BO
nly+lp+mldj+h3t1iNp7zq74g3Pnpa1zptfM0VbloYWAmmLE7j+G9wI4IXj0QuzD
gSl6PdEaSBBDYt5dGJnsUFzEilTzNf+Bj6m35CSnhCa+X7OkJugLkU1Md5c9mUVm
bEOiWK4+FeYdu3a9FF9De8gl+2G6gBAKtYpEJmeyzncZRULwzYKV6sovWEmHtBhJ
z/7PrxsapITw7ML1ZGX4/zxyQXzKkG4RC28jhxzvm2E6odWZ6uElsWSi7I5PA/hp
IPoilJereIkVRYZpnNxwUVnanlPBj+TmfwCWx213zi6deAOf7qTTLYXBJBC5mH3b
zCjaE2oU2zmYoac2mM8ExG7Z0qaS7z2ToxiHJeeYbsHCPDx2ZUg7ucHmZ5OwVgJ/
Yj218ZOtzNU8192yya/3tVPEY+ohsmuZDDP5wnQpm+36ziOf8jzwhI5ynv4lbP8F
cHVwG2/zLSjzOS1JQ/k6nF7Nejo1Dh6q2rCjj+0XlyTEec/5RXNUwadV1MEg6wJA
QaTSbp//yXtp+ykT/fBIFgVf1CF26pJta+ItM2InUXEKmmLV9mZkxSBOUQ3xrkny
9Mf6lEykmPi2z5eVHB7NwJPq9JoJKdQITT8DsZiQpWGev3OxQP+VQYqN1F9QKwUe
Ck0gUgYWH/oUHhg1acOlvFoEks8684uuiuer4k2u1X2JdXDpspDMpuI2bjBJR6OC
3DePFpw2l5l9w68oxZnbahFCIlYHOb1Nmqmtx77slcniVNiCdynR5H7AbCh+2lzE
MJRH/ikrmqatYtnFhCWvyqejnZBh7DhBPpbGzyDgi7kff7DDLFRTmboGMVegeWdV
VWK9k+4Sz+zQtQTECZPqV59nspAdeWG40gGuxOYbwyWvuaxXtc16aBnE+/fvcZfh
KkstRMP+VYAzOPdagl88GcJmGSoMYLvE04HxubPhV9mOVwswPeBUGlhTQEv/BquE
9sR7yQT1lsb1VZYJ1Py7gouJHQvCOwjvMldmh4Qm6u4LXL3VVBBghfVXP7yk79pF
DRrPZTeNZDAVHK6BPC75u4ysEaGx+csbIdD8QgIcBzJ0qptZiFjMgYV2yOxFnp0P
xq09gBakFJIUEbmLHa/W75LV7BRuoxSBx9LzwVKF6++EYOhhtTepdiy6Ptb9Xiy/
Mi2VBlY/aWF6fVX7GAmYMAs+Z9zJj28KR2gOz8VYOaYelhGqWgzcOOT+Q569ks9u
306/38kU+Yx7C9L4nMpWSb6tDm8KHEudx/v0RORzY2meJb8rHmBsly3G7+ajTLHF
1JNan0kUJ6VJ76C2MOGiKrONQMW904MdKcVEQgt+bTc7ksKiY7nqb4euRePf9lIQ
th5vuP5mfPR9pQrYTDvyzDeIQYIUXSGu9IkuPE81JVKfBeewC3Mwf05giBz52QM8
QHFQG4S6C7kZcBpfL7zTkQJqZlBb6sgxhJHW4u7kDIETho+AYpx4Bd2HlB4jJoyx
gnaC0c5DNjn04QvFh/9LminZVanXv5XXHhjHSNyFb+xWTG6IB+CFpHLHTx90c0Qf
kbHZ9WXrzgTNbCC9rM1p6A8SbAl4PgIdCLSYJma09gitxJ6T1yx/36vpBiHuhjrq
5CKTLcXsH+OJn3yZ83B1/TAPkWdZdI5ZGN1RA5vWCIJaqAaCYjGhwo06nblmBCpF
I4J5hMAaaQHc6LY6qg7sM5HbvlRK3e0WGMY+sN+/UAIcqTy6LqsMJ8p+BXn+MWJL
jmXFH+NrbPK6PtkjeerTnjnks0iuQmyHbF9MIauaciHrmR7FXMPaKXhGFe5yFFXE
ultOMnOVrJ+iYc6vrftPpsTgUgG0YmFUMaHdMNLupbUUSEEEDnAKaopr+Izh7q/T
nvYCawtGFegiDTpSPbrNivU9jNqrLnzjOORn4vsauHMmQWGiV7tn4PSQxGs/RPWf
Bw3MJtYKgiewkU09a1PxeGh58sHXlfpfz7nuyX5rx/buZcyJGmg8MWQU4nE0JQFn
3Vt08CKr9wT7uPpAm9Pd+pNKLEi+BZoI+Qv0B99R8f/TSENIUi/2LjCsa8Cer3Af
tiwrqynAz9oOSfsu7v3S2EywoQ29SkFX+7X8iualESl7bqUte/F2rtxEh2Fmm+D5
3tv7Q5RsxkuBXmwm2CHf0Cy9hqSCTyRDGCk29bq1AcZYDqhhw/NKmSLSBpSgxZMG
nX2xpfRahaqSFwi45BPw+AFcNfaSN1KTcN62sMCcIZuEFfYOKgotjXe/i+RkMmG2
7XdWhc6hAGKl0CmPLvvBYETz4WW5gAnP3s9UQqFjnHT1w/rZ6QLX0Zad1jbV6Fel
eROditwDKJP4c8/qC3ijl+ESCNABiytHF5weC41M7lmfz5O+RyvBsRw2BBzpCGrn
9SQ5ItTn+FTrait1Db8D+rP3EDWPa/Uq8UXsI7STFg6i33tZcEkamdSGIefzTmJi
5+/J/zFbaf5PzfSvgkRenRn1fpqSwgyNJfKemYjNiQYs73LJVPcdPXhjB0SwSV+X
sF/oBvPGNp1HeaiXfqH4ZtkeGZcC99QJUvS/ihJHoaPZJYX91iMpj4T8b5XZS6/u
e53Bu+Itidpqhkd3RG71ImIcDYmHD+xX82rgfJF4ZvjgUOuMrZsC7l/OqyY0XiXv
Zr6GWz1IHWm5pV2RLDk3sZNmhwKnkrdYFE/levlazXASCtMNG5Nku4U8enxMRjrN
W3boX2zcGimSEuvZ9rZLZT3wm3G1YJTrqOb0v1lZQZsZiyGFIapFvb/T8lO8HGhm
uVBJWg1drTSLX1wdab82Fk1uQTJC5GHrJbBcG2OI90bY4w1BPnZ+HwdzREG3BOtZ
0KToZNcJaSjJ4uWjsDdz64ak+oZZm1tV4dICBGdwXAGg+Hv4T/OWPFlT2fccwAyJ
kZ8PxUaGvnL/FRgXSG6ek7khSoyIfXV2rJXA0MtCGC54jFT6Z1uUKRhXUPxnM28E
0lf5++Bgzvk31f8ju64kZVTDN1QCUaGUQpUycT7mSATSBzOpyoXnhdYbxAdGLK+A
AFzwz9EW+ilnK0hVmgkJRBkZtz7CH9VQEIOEjuvAiwYzXJ2wMlUyVNaurT/Pmvsh
CtJRQUXoGmkhctPl5EFmdXP15X8TQ69isGUzW8EZwbqLgvgUikKCj658F9tDgqOr
1lrDS8YLOqYhv2JHR7cKf7jdUifrUuyKKzRY+FwaqWzgsFjGcZRzknUgCrDUOY5O
W8R8f2xQ4aMPDCnWGwdLOziSCiZKOU46oMH7rZqchGyv7WL+/lKJqPYsCAjxYTp1
/oqgXHJt99aTZHKq1pS6WsOUDN7bM1YU+eFfgmgFps1FETLRLA9qT3ZGIsYpc1xl
GWJ5eV2/877dhwwWKJ3Mqiwwf2b2l/KLeXTKJWGb7Q91yzRZgKSgMOVRmUvyqcd6
nGFnfrq/wuyStKpFXov5/WHHw7DnSEcR55YZtcvEkPYH763SqOR18YIsDhTHqWDz
md+bme/iFhsXMH+0qokAIxn0Jn3d2HF6NzUWy+py25LgdJYvV+vxmZvEoETvZ3YX
/v0QJkt4WQ/2brgjB3Vw0kek0VLmrYZtVWrwDH9f41ldMQ9mFn50KJk1izIBsaRo
snLkBqI61ryox2E+oyaA/KddXMDBaXBvO/P95nLdCEg2JrUOLknRQJFkA7Okiu26
bBPbHziUwYVagSLFE3Ac0AXvDK+eTPa3gultoG2SCX31hhFmNKU9+ZtxBKEsjz9T
HcoDNoghO+g/O9V2WVvtahfwiUT1v5j0EZrxAXJpjcFtbm34l9E/YfUpL7X0brsN
azx4ba1zhP7YVbCBBOFG4oYjuGrZH6YESoqS9b1fo/k6AXf1LJTTB1jbNupTDyCL
eP1JLJm2A1Lu3fGWjiWj9+2+wLzpiHrQtFkL7tIgiQMb0Rm9A5KfV6IbiDOFx9EV
OpDwEXiyFjlhSuVt1zj10IB9Aiory4LAt8Qbo9Wo0efrqf3baprynasKCjTO7sUO
N96mLMidXN//nXN/1WkNDQeBqovAjxjsHEJkBb9kQnh9i0p3n2PGtwANo+8R78rb
tmGvsFXwrKvgt4Ed194kxl/Z83SfQ2PqEoa9eIvM5avBUSSbGk3vdhEpvQ+c7DJH
85HwairOiJIImkJqMRdFGWVMkNLPfHrxiAHPQNL6Wy6X1MowRkquXtFW2zo+h/Bp
MMZ6YZNSRWuq5liSWAMco0oQ++sCcA+MBQ8cccPP4Eh73wPIdyOAmsxdIR8P3o5S
RwEddK+RraS0z4hMCy3K6Bx+jzJkT8i70EDryKi/v8G/FSYl7tXstCW1v0+gORWe
e/X0dntxbS3PUni/4nojGw715+erKfp5CK2YbMsPzPDO+tsYr8zE44291PCMy3g6
g1wVgeqg5EKFObK5hblSM2CXCSh0lKhq8CO7RlaKYiom9XM449z18A/EHnuvKooH
7bVL8l+/gBFStKJ61nYiTBat0jxyF53J+kQ8BZB/AHPyBHOFGxXVVz/Wb8d0JcZz
CCRDvKnndMuYYAq3pZrUVrlbOGPj5hbj70WYmvo9BtcBCKI4vQWBKlCPNTW+sUtt
yXQ+TZI2XiEUpqmAM4X26rsTzej2sgLCsZWmq/2ke46NMIuagfi/4/bumGGTtgPg
FVOfH0OUdhEELUu1VOmCvxNlKC9znTMtCfxyrlrAPc4GrkTc2w9jkCHIe8PL9e6t
4UcHU2M4iKbi2SKPTuLZUGoo188pv60FVnJ0s1bNrSLVNDg5pvf6BQbtltUMVUuu
Bb4yB8tKtPvXkd2tTY11tSPy3daFEgRZVKmRkKSCBYs3AhL8Z+ynSKzO4T8h8Avs
XTtAmBXrPqzR1RPk2t0LQC582y/N8Dy0xrw9v885RIBZzAfaLDoH24HJ+DX0MNhL
D+f//ncSbV68mRhP7lUhJn3Bf0RGblOz9EiH/dNtOT4j3H6uebyKirBqyGrkkfbn
zZf/joPsrKSFp3H8lTP+VXP3PSsQe9XqnWqNo9P9iUkH/ADSym9sc/bJbqCS5dbq
0W6Dn5EEmDPNYYyJmV8Wc5a0yU4r9ODvmNP/NtiyAlK/0Z9CgQzNOmQkkFHk04gn
978805Nn1RISUgquq1geG36LFz61dwqbZGh9znWH2mAcIuJcSrvF9tUIHcEvb8h/
fiH+SxcY59SZELW68mC3pthvA/i5AiHKjiBGXjk9ns+H5tSxgN+/TxauTiNlmY5E
yooHTRO884p2Gc2JMAXFw0qnmya9XgDN4lNAqONFHTNAwIICOl0oYQDDPU6TlVcg
Rj8iBwNKdzArf83+EQGpzpscuHdna51JQPJqr2tAJAnc1h8X6hWkN8YDV49HK6Mq
dasQxwGWz6u675OkfH1/De8dxeJaz+/C6kSh0x0LBeNyYOfdkAyo0bvg2WwnGUpW
yfUpsomlzjwvfcvGqD0yw0HiROk/bAyWbv9LH5F4L69PZxlrQf4KWewvidEolff8
ZkXix9gtlZHucRrExW94KbSeM4BHk1uqR50Pu5aVIdRmF8es0slCo516F2qlAcES
1OwhAUeVJRaA0niKeipLm4sQpbHvVcWaGeDi+QfjvxdtqI7fFLdbLhYbZ9HKr+SQ
45Uyz3qUjADiIgJGMSYcgRyFwcb/4d2PB0NjPf8FtktJ8Jdlj38q60pcWC2FksU1
SsOg4ElR5jXpoqv1phB3J1+BBmgapnd1qolDTliDtG05NpR4hFdu6wPE+1lefplm
7/Iv1Vc96YmKqEg5WFEHhWsEgEpT1ODu2MyUzDky55T8J7tFs1+RxbLyQFrqkipL
ETdr3Tc7xvT1TJ6FY50pRKRjKHkCH4Co32uhGkh5eUVQuZ3SuH4Cdgq1OUcq9Ikn
4xX+y1CKyQNjBgLvSZSeVcSZxCxnyCrp0WcIPMmxPXxVR+BAE+WeO8Yt54Z4l377
s3j7qLJN2p1dzgPUqwPF6f7A4OHN0AIgmT0iSkXBOWJa/45lI9nALMrvuuf/nEQr
ynVfPWvzwRbmz3+ufQzUaiANu86TOBxS4WdqSmNyWhiO6+KZ7+zpiaWgifLHiVUI
GuWEQRH0bCjQeD6byoF4K1ORSF8JXSuE7XUGo6kcdOv+zVmq8iqY1M+1Ebt24UPj
GhHZtbbvYQyJyfOXx2uUvooz1Aw6ZbZ/SIqq9h9gb1IYo5IfNWPYIh8QTHbFO+Mb
WnYXyy1qtcB8BCBsbhFWfstu06TYP/MhK7D4Dv6zPSWUPUmSDZS3zubJl18YtlFQ
Y9F36sE/LhYAL/pkZXfsgGzY9BZ695BwHZSAHLEJNUYA8hEKmCla5wHiHciNtow+
O2kLsSbRm9yxcs7lLhFMa6NVSbD1ix/gSR5cIKbmQmiYrxHIZtSRnmNZOivn3g8l
GNMoUIbQgNoVt1FC2ALyjUNohyHLUvYWrdYgupQ9TFyRKCkqL0KJv79EViZgUxXZ
s2TTYQzjsm2FR7KlwoTouNnxzcQJ7GrP4NtWKQ2ceTiFfXmvtELD3bZ5lmcLQPo8
T/kfKR67uAjsiQpD2l+5uiHezzlc1/C1ui2ND1+4NeHAP00OTnN/EkAAIPyodM1i
zjGshpjt2YvlOTGmqaVi5ufD5KiWS2AO37ErxrAuSOjf3er2IfCXoG/7RSHiD7zI
wAy4ChhAu7G6jwX0bRA0sczB4HaKSCzGIa5XBzkfWuPEuCNKR502LQ4srXFYy25u
nSV523lg3pF6qKFXFURIjj7lhzW28rLZA3DaeTrm/jPD2YZyrfsbIiJ70s1KPNG8
jsLJJ3G56j/q4YUzZwwr/qR5qjJeoETYkOkpgqpIlxb0HtICmN8A1HepjFYiCjyN
2uLwLZtnguopoTQBPh8yaGAYLU3NJO/MUQc38/gjrTuYpM+Nk4rFQ+d2j+8eGnUG
Aqc6udod3XSLL9f4xlc73VbC607W1IWe16U9i2GnarxWGytF+mPeh74fHYkACuTM
iUzPKeg4tv4+E3BLaSUOXugR0PuWxJm58aDM62/w27Y5s1C/Wwq+kHb60VoqaXfj
sOTxLp+zbNwIuIqd2wZKFKrSQTJ8JBBEhMA1WBU0j4vKK067VMSMkQe4i9J6lFAk
4+2rXGtO5NZnsAkfq95+NlfFVe3wjMpbbor5Mc2ta3ZWjPey9HqGwYoJGBcCpas/
HeGrvjIEV3y4do2CeucgdXuavjCpK8cfqnI+BwkHBo/CZA/Yf9pL6qbd1FMMaMNZ
p418x1h6fsOJpvaAvqghA/VoTME774KGud/Ny0bnWyo/Vjz6g/OkUyRzhzixhrKI
9g4yNIbn/cBNLAZF38zK6tk+0cAy9oUDkAqNrbnJx34b2N8BVgoTUWvdDMOQMIdj
9P6wESh+SgMrjof5cvXd8RpP/JZYWueXu5MZkFuh/MdtTpyNoB5UkPXUZN/oHugk
uI9QacIQOKzutotl7KbgZzHp1cJKFGlTeFp6AVeZuL5p2G31kk8YCTg1MJK31YfT
Mh7I8f+KgboGeU3vU5B4XwNnoCBFUfDMvoYiT0BN4VQ5VatQepQqiStoIhOo+XPY
J/wZgoGOgteVln8jbz2jCuP+xPpTQk9NxM9P1C4i483x4NnbUnqOcGpGc+MSFWpT
xglNF8yKqTlWMF5Sw+xkZPSMTSzObzTMsQceQGuuoNTJ63hpYg3O+XXSuc6Z1KLX
rcqFc07LUL7p6Suhwb8EwionarBZ1CtdIUt+HT3obdu3OrR/dPyn9AzZJ34I6nB4
jhv8t3hAXqOkShRRai4wsPiyGstlz3RVPooH3NWGXrz3BJRmI2axmRE+1qT6d3Hv
KVoitOPvKo4SOfnYb9u/nAF4eXuxhIfS69Q21BzJJsD/gMa8fEVPcH6jchnuaZqh
YBkwhYDhFfUzFE/Gqcx6+q4jilqcaDqi9uLtOxTTdqI4quzAHVezKQ3UYKsrU0RG
5YvHo54Tiu3mEiRt28+Al7IYR4eXzgPP9cEyZSVkEwg93v40MVNfC/WSn39eOVjG
pp6T+N4l+BTgv4v7JHyxRunCWCP0gGdUTBu4afSSRQIoNGa1O1wDIP5Qa05DAjTx
ffd12bOAXKGEPowhEFkYGvgUa43jXDsp8Pg2fNSwSjRUS4K8Sipp/A/KngiahUkc
gmUeflSN2nC+W+p/GpFU13P1d4WvqHsRHmP3iljln5T5jzG404suNBrQdi0DTd/w
+jzkgvytIZoHcjphXBm962CH48fmyMSIcMNnowCyPkvRH10DxvICu/H+lw8izCiN
RSGSNLaxsV8i+JrFgqFTynlA0KyieqKeKICf5PIYVQ8HELvLZ6qXjxf26R548P7r
WLj0lwyTIi27NwhpOMxLv3kW2l+r5pffM+AOVtVZSwwb9ECBdPDJOT+6KQLgfMzb
gLbzyI/QadAtxP1QeHvQzS0uGUZXO3qoIXJleVLbBNjb3yBeysDBzXN3x+q7+Szl
wtAc4srf576tAmbVtvOND9G2XwEY9gI65bj1jxQmlIcnBsuSw2ssx1LfsKshqIFL
Gsq0VPcnMsGjYZZX9z0QNmjzWu3wP5mCUaG5kQX57eBRxKgjyUtvGQvMpEnatuSa
GZWo2Mr0AuaDB/iiYvzQif1wWxEWmA+LwPrw8YEHJ6CVt4Fkgfd2uNW7HIwjlZst
yoW5TYdRFhth3VpPYswAw++fB7XyVW4ViiAe10RDk2425XauaUcNDKrxzSZH49Nb
g2xVAEYcp6EayzHXYiWst3QlSqaqctI+DmuKMQ0HxFXl5uh2Hkw2yIQkPrXg3Kbv
2y3+IqOmJhemFe92MUP2IQ1QgJsfKPEdG6TfjK1qM7cS9UKSAXnrN6z04TGy0nI4
lJ0H2REz8MbST6V/jhlz7SDwvXJDXFXpJSXr11MeOQJ2hogneLxha1O2G7TE/yrQ
D7/+ah5sjh7s88MfRQ21D+m9N5ls71lLMiAXQ/wHITT/XLw6OROe+JsVXLuS1FZW
0QSKTQ9M8HGKFqLN3UNquA9uVve7eBXzhgk7cPa7eRj6pYy2/Wki15h2G4W68IEl
V9tiGTiJFtQOJ2vkN8FtCxcQ7Zv94CbvbWEp9/Y/5Wm8wr+irOTB93aOwiRt+w5s
eJN5L2G1f0EwW5Z3YYzuSgFHN5gZaiuHvvryySp3qafqi1MJRC/ehY+1XdLmKjDC
CAyZiPNGgqp6MvlyOzMIh2u8uIvyDo7MwH4xyQ2MNWJ1FCi9h4RiZfLEUyp4Y573
p82OW7AR06nG1L2UJRqenTa7OMJYm5payr79+sTb5gdK0ddXVc+Gw762rFka/lAK
SXFhzofKUg0NOT7ejJGv4KzuAi0QNUHw01nhSMaXEUkZahNbthfwjp0nNQlVisES
sowRlW0DBZepKmroMemolnBBaMxf+sBZtQJLtA9E47XEfkS50VJMnpRlPg8VJxaF
op+Ep2b4uTlWURIJs0xPHsNhIbhk5maszWZRZXx4LT6OHFkDbvGsd3VDy7u0Vf5t
w8l11SCQoTHuwe2QpdffYHUCE+cSAsfHVPt1gPwdHiSI86prdlNj3s05RA7qJi0T
3ulcNByDuRZm7B4ceuP9KRKPi3YDQMvw5r0Ko1jIFgC4Z3ToXFt9vYr565ndEnYM
bzyoG6qWXm7UH8/hkyHeV3wOjieclP/CTMyZuP1ZeW9dsgYt800rZqZAjaDhPkyO
Kfx0TdrAewJhUo2Ycdvcjg0CY4VxZVFwoGQCZzSXSy7fPZlZpGtFt6y9XFLVlUwl
i29H2R1GAQV8WuEXZrjk/GTbtr2OZOv8SODLUZKddnyRQj7NUn43Hmm/etHjbnyR
hpj1IuVLdW249EM7QF6WTU47NGkRyI3uI6CisNn6U37HJjyi3ASe3QLTdgbaFzfI
Jb/vi49wOYcL8+uNz4IVEPh2GjWpSGQES8deszAMUwHuMF+yuE9QattoJ9A97pZ7
xtjghFia7afRRjl8mxnq+n+UvU7OxQOcYcR2GYykcGW2M8NOZxp42bDx+H7JzxOK
Hp34eYAqEhtY9Trjrq/F1+VUUQVK2XyWWRLIp95zn7aZBcy4uwq05P0S8TxtHs55
CJPzWJAp39i2xcVwsQBk5Me3o6q0D8uilZF2aJ/dH5DkXBEgZxR4bVWrFYNu/XXL
IkKCsVWIxTOMLF5+cxr3wHtkjqCcrpxQeHNfsFtvWhPGTiuihC/JSj2hK5A9QpdU
KTaALYUc+Qbkd7MW/sV/bgbweUdSQCdQTCdgLAdIkbNMBFGDWYkv3bGMkyspURy0
y4ImjNVieDHChUiPjxDwEVInMoZW8PzCz3BS7BmJp1j35rGwIuf7/aciH9idxzx5
/p43GH3rnr/v9lfDLEeLM79KliTqg/t6sTuMb4HNrx/CjFP2ba+c1aqwW+XBAEVp
eMNF4W8xbp/H48dUM+WvDvUVQvkno+azBi94WbRslgOPUWFGf3yvIAlO5u6/l/WI
7MdwrCk+VwL3htD86yw39YyNSWUl1s62Tnh/7Fh2zcpG5uNzku2J3sS/BkMXfoOn
WOXqwa6RDrbtqb5vrQi87C5SuYAyT5xUoH7zJJKcH+X5JdNeyTX7FvBSm8gogxNF
zZD8mOl3FrQQmqhxYWYGB0MvnZ1B5JV4BFWPm+sxrLbgiuLUrQAnAuDh6bGiCG0o
GHzwFTC/ezKeY48/iJjynQ2087GnLpfjeP3A0Jtl1Vp0V5fhsDTxvesUfsiZLmZN
Akhf/AffezqvbbL9wHFNFbQ3CPocT8Svipxy5euPkyM2zbH6HrquAzc0II/BOwsj
qVX0s6wCcgSc0Sii9WFqCzpKH3L/Hu5/FApbz1JAOdlYzsYYq+h81oIrKHx+6J8H
p6XHDz6L4SBxHm7E2saHuTS0U3wHWdxLn+HCjaH+7GJ+RN8sHm2Hyf9Xe7nbLxuz
2W/DqlS6hyCDxESZhOJglBR22GKLwvx19WrxlbtRrRliRFHKxsuRsqz4+1NZuZCx
7bvg5/yyba/w6ktu5ukloS6q+cLyDAfef0RjF0y2Y6Um/eQ9xNg/QA66RK2Y7dyH
yIvaUc7ZFgoveAtb4XfW+1Scsw64GgvVZcv2VKvZkI1A6CnTgNu+uqmZ4TwjvjOB
vk7RpF0S/1V2opxlVZahobFXtmHZPBkueTmM9mU69JAQDI87yZLQqwnJblEp9BDX
f3MJj5nF09A7s24w4qaNKOlFE/vS1vzo3H5sVEyTjgPnvYBO1wVt1jHV/z3ACh6P
vBiEzuPFVNQrL+oARjzSOqeerqYNFR55iaN4xJBP38EcDwhOYXU7DriyG2KR7QNL
Po4EX35emsjBcDxzuVYW0INS/d6Y6wGQDbK2Qt8HM3FdXwYNXg8cvuZES+ABHah2
gcqoO0GMHXqi+i9qHBBga3C18dMzd9RSq/ta08omhEBcMm0Aw4aPnmeKETkJnPeM
cBsyCEvxjvEYO1RMBVVn6TNQE9NTesxicjAs5vsHejXad+pZGYr3548gHYPRdRPL
MkpoGQ/xzdEr9Q9/MwTRJk/Q1rP0218M5t86ItY6og1mrYA15K9onjJjjFiAfxim
MzcvrpcyBaD1jkVZ0NFaBh60WTDmcDPPJMUI+bm9wwNE1F2cU15CBW+hGJMZzE/m
owHTBkc8sCnO/U5gGP8sVoQAZX94Cqeopz1sEpsJrL/RE9KNX7OgZTbxBUAcchxx
3EGgYe+8IKsZr++BmPbzy2r6swoFnnm16VrMuuWz5NyFyDDSnEawz8zZ8v+dfZVn
tDnafVYS3urDpt7b6wMrdrbZSQYsEGv6hCUG46sj+MYQ11Qp/s/1mFuon+obMFkd
QNhCyqhU9Xpy/nOoE9+LiSZHmGysLoLF8LHClGyUBXM7/HyEZiqnGaAExpeDi2Gg
ld18nCfvxWGO5coQ2MW+yhamLD/FrMVmacJOpovBx3cH19t8sokcUCn8X1sz3vyS
JuOFW7slXlLMJyakXoTfKGrf4CoJKRZlccLGH0cSVwsbgkHWMGy4RaM579zlNn7a
Uo6vyR7CtDkeKBWsS/YPTb6AH76iYCjKjXub7tsiP7DvOo3SA3DyYBO4PrWzBVIY
7Y1+PYaPSqzJh9Zu2BJibo9PspHQCAWvVOoZNiNGwzijCS7xGu070QTeBO6SU9bK
1MlVjUpmEsKlAmU1gOW4L4P5iyuLrHSZLDMGv3eimAHuiynladDbpYDClJBXlsU7
w988O++bdDFq6zfTt3LWupHM4SgfWMRsB4tMix4bb4ud/pVR7THVetfShlkTtfWs
/1UMdBb34K9sHwV1Ee2EuE2thKVsyl3grd0rZrJ4LgOJ3yqqjf5iJ0W3xmCzX3HP
NZ2uXv0RMrNu7X/ny3HfVxsvwhVUBTxWdIQQ/po17yWxZ3BfPYuhAkQ+/+8zVKf/
sJuzc+fzSZ5YhBj+IAdOtan09AVfejNp/rc9k1KavrPSKIBGVPAvUA6HL2sUKU8q
p2z906e2/7gQS9Ee0vNp8dtMx/udxtvNIAC51RRdJuFW8o92bmaUdKAbL9YfqsUW
oE0c3UsYBTdBH8OhIBqlQ/4Heux5idBBe35jGSo8IE+otsxdCO/xaDPgiD55XK+O
3wjcSqIJDzrMLv99e2KLrBA12lbPbIu5PrLsU/4LtF82CFmmNNLS3ax86ZrWOvCc
eRd9DnDPgwF6qKz1Uwk0GJIa0+DTYmudZpIDZr1Jab21YAZ1XiyklDlGiGOoyS+0
q0q4SKo3wZXaIsV0tFUYORaSCaWV+Kg2DmFQi24+obZcBFNH32CA4GKYn6FRWk6k
sNWJ4YL+RwiL80EerFRtHj+z771Z5dSU2CuR4nP7uYuFyMSUeW/S61uY19NCYkkg
3B5EkHQFzyvbEU+4Iwl8YCxgQ12ZuDAgMqSrhQRrU8sX1g/xllrUu59JfVFvHb3D
7Yiz3EN/Nhj0umKqwaPKyqUKaa2KjcaZ2P6p7qQPUbNjaS+5rxbcZ2YjKTJsXEtB
FYkRSW9LzImzdyAXeOQ8M/qaqCftPWCtrVvni9tPkJkZVi4nzl3cKMwdqyzJQ6qd
MNJv7sJxyZmGOEEelKPbnOXNUGxw1cv/HiDTnPQmxKa4xK4McIenkD+xQK899GZg
2tVtlNvyu63q/gC1cpR89x8/6zKPLAYfK33D5tFSMnUVui5hv15XeL/xyYPc68rK
RzHSyUVfm/ztzp2LZD7KFIn0atR3+kdSY+RcsFOTlpkXzdQr4EclXik9N9qnC2iX
4Ht9d8tJP1IKb9JWLypZ5xJqvM6WY6hAc1oqh0i5axXjTmRtiPlpfQEhNBy+nTH0
XUgGNZjCKbKn3ESugolgltTilOzBL50BwIlZbyngFxznvcGsk0PUAB/lXg4kzboK
6WCNyrQlRCBlKg7Vzp9YaYexNxJ98Z4tNp7v+27LblIZoCBFWWi8cChsymGVsmX3
+hJiyQR0j0OjDARoOmTJ7OXOWctOr1HbTTsc07vog+mDqIVICjbJesLHu/kuypek
oOEI9WG1UiyrA0KLew9y9fmCaY9PQW8i5ECmykrMhudhbPQVe8XGhja8WfLMvN7F
NLx5X1nmFtk1EAGqbSIPtGHQKeGgJhwp1NvVctLdmJnmB5AupE8pNHYEjmK32eLo
JuZ1p9JQl2f8XfOd6IgGMyFFR/S5BXq3IZgNuTL9de8breHnjbx+FHQ/deu8SBWp
/8KaTBBShe+XXRPMRFYV2AHyf7YcsPVIBGUm3awr+ZuhrGxPjhRPzEA2RLCqQDfs
gJrsz1CxkOhYgjYJV/7oyDiohEYmd/cPeFztVUTu59327c/54nwmqimbhyRU5ucO
s5uNwI4gP5VKdVoziESiWHGqod1l4wdESwtXxgXn7MWiTRPJOMMlOgWw71jCICFN
6vxlL+Xv/Lby5P+uDGU6sQaK8H8Ku1HiIH4g2IW3vNwYL9dkw2ZagvpeL4jbcT7E
oYhI55FTuadXVY6+DKzbKgFDgJ4Nn2E9yS33v1WxSGhacIz4zJmOrUIH5CES44Ja
Inqz81041oJOjKdLPTGqCX40BtYXQr81+eHA93JxCoMrTEcYXHoHeYzJ4RD/lvC0
1WtkADJMeUZKTAhqKI8A+pCt/nJ5tXRqCQRDebhObr7rcoOdv2hn35xIJfTK770B
BIw1lhht6twdnRX1n1AC1MyiUNAS1KO8D9Nw+63AbGz1GxX+O3URnhaD/c8HjEWa
43S9rJJ7gjVKjTdRku3ldBdRuFZBdIUpkBd2tmAFK3XhpEG2ve/uVTnBAvVUPXpw
BWGr1JMb1v1n+fsUH1EtAiOzzk88k2ahnDr4QU6bqpaNlxgr/4m4iy4P1DQ8yFZo
F+LuAs0DVhq4EVxW1okWAp+KmOrWjQAYwL8SQRe42BG/KfMGUQ7LXoUZ2plk7IVQ
oe+mImJFmsbKavPc+IELoAuGlDDhG2KsiljZImwamUctEdq+hZDC75S1mYKOHvUa
K+1H8PKXaC0Fy+AesgVGEx6QN9q9QRhqjyj8IRCcKR79Iu1REYnfh1b+ZiR1eZ8L
zErIidHN6gFW0Nza62nFjR+QGPSBE826qBuujK3GNZIxyhby+C+dsQ3gJf4DXT33
q53XTE0Wa3i6JeYBb5+wLPbWxIgwpxT98SHwU+EjVg+qubV0P9wIvZ5+VhIFZR4q
yr8WQAgPfcRsY1V9v7IsW/a+Y7PmslBzY/MU91DaOweNahELgPzRlNOGfgonSu1X
0jtvssEObgjPb/RmvfKzVMixsRoRdFMkUZBFnQbyDnIPN29DAuIuIrzHQXXVGwvI
ZsGWbVHKkHUBC5ipSF9V5YsKIIsC6xQE2wo29YhFynIyNi9iWlTKwdNXEF0kcBUM
u/sONsqG6HgL5baGM/4+HwNhl+2pqkKYj01/KAQMBIylLmi/+CmqH95NoZM1d0mO
O/cSfqaJ1NctRzzKY9UujkagRStlNFEjo4EQBPkNHra3sjYpjcAZ0HwpK+eAgDtg
llfmw6K1YxrDqC+J6nFrZ+/4lOnkuhtDE8Iv01ZKmVkGA4Hod1+L5kK+vrAshNWZ
Q7CRnhoWXsyYg4G36XOAGKCiJGoC5oxvBWoJczZPzI5vZw2anibT7fLTsRPChiKa
Ryq8PnxtqockxMWd43LDr+03nC5yKRee732RfNjmWw0CV22jDn7M6nVhVgvwm+v1
bmKqp1J6fYorrTma4Jhk82bqM5AXRpj5CW1VFupbkylVrbY4aVOAYoyaD8H/n1PI
NDLlvVN4HcJfkhs5OwklKUD3uYkGn/b7nuXexWJ1NQWGLRRUhRgzJBhaurTE8Xmi
0AhLkzXWFwRLdxCZJTOaySgO/K/5SFqSjuh+M6otKOWuGX9bENBk4lO0AK3Dvavq
gw4Pm0eK5aQxlm82ZsB7+KcEoMUgSGiRZrCv+sCuyodaFagFuQ+1HFzMJWDeU6Ln
W8LmTb0bsuWiD5jbu0nyVqqwXZ2uu0kQfx4Q6UPbErSSYT7CCzd9gKz+UOqUVyz+
l5sdI4G5nGRmdSu3le7wcaLiYB7eMaUpYGWmEvvGgz/sf/6oytPL4YJcqdfL8WoA
bLcSzaxjadRzmeFnWrfC5PjbQ4qwkrq0bRRJceqmCTXwfGwwDdIaZS9f5njN+hY/
7reAKgXVzPde1Acb//cJdPdLoe0woA9HtuCwtQHFrg/NY/RtBOMJy++3Xi91+PCi
9sdJwFy3Mqa1rb1ky70jIc/r1zVXsQFVzFr+BXHHUAlROf2zB0fvuhQ4Hw+V5N4T
bjQKWWG76vVnODSu0zBbJtilgoGo1O22Rw280TczXzATLaKgAzoYYAzFhCtGSdAZ
45r3Fyvn7Q4l33/++uni6dNhLC8H0i/oMAkMJgtbi7DsJRc7hgGdnH7lTxp2rtw9
efF6zulUiwfyQvuWqLUp/Xqg+p7o+dGlmVCCeYTjEhXlkvAZvqIlV5yOKaEm1fsp
khJhVr0jh9RjiI2CiK08yfcz2CCja+vEd3k4Yp/s/FFU7OHe+hKm6pooE0JQ7sjJ
3KJnkGoX4zQayalNiyhYxRlSXkjPtBUqfTU/l1VAJH5cmT48okJJsNTdC1Xnk0py
9ZdpjVl4nbwlUQmbCUDO0kGW9pkdXsgZvz+TjiU/jMB1X6cpADqhIZouBzc/gorR
sSostbxIHip7dMMlM+gdEbEeozmRZXPAmdv+wHmEibq1bVdfDBgMAL+Ss3SP8LSF
5qzRpK4aV3sQI8v64LIi/u0EPow2jLAOcY19E676tPVDS8xKdgZQASwl7Kzxhbpy
Rfa7Imc2D4X7nL03zfwc3pMkF3xVeoKi83i/bV+E0lA2ub8FjCpq0A90XM2uQIVh
CdGcj3yFbyAe1cH89OpSZsZi7aoIEYbeQmfBSk8an8Rc1qY/H9yghCNxxAJMJ9Yh
v/KmOpN0QJF2cT42hlD/61fzdJfagB+9Ta2aM30Z4T61FQBaw/gDfLifjSwZgygx
V+XHnOVl1QU7AHZrA2l80VeRuOgxvaLJmn+0ohT/wvqki4vf0N40MODAoTiTARbm
cJexmtpKT51DUXD7ERAkZvByw5zkSjPlCpe9IGJRa83wLlEq62SmzmYEawemx6WC
93grMF256Uqc1MPJd1EqClxFeRQMBqql/Kze02d25LpEHfT39Sz4LqfeM0Qfz494
wjuxVehp22V8NKM5LwnWBXDgQNBvGHqOLTRtWkzcBgCedVI1CYNG/kgzh9bJm5gs
sPM00VNNTpBUQKbs66q4AqicnMd0cj/s20zrmvMxj8QKI6GWJXymjvXlUFrKuB9u
YySKzARL3Hn+nXh6jnFJbelrYZ4QUBmMZwrHXYLjekpbbVj+ouJnxKCSz0+b0sZn
1uwBcviHuqQQprfu/ihsYEYo/mw/QVh9iKSE0WSZLNa05lXfYYLn/NRnzsxGzyjZ
0FQdRnnZKUapGU/TAx4LxT4Oz+6hEvziXWHZn+dhBtSkQ9msTQM3rolG0GkcJjDU
HMzPZlgb/LKwtyI17269nhjZawxFQzMz2Pdf9XEh4qJvn1/bAkzo7WbAMru4fcXU
wpq2CkxMCJCrAv5PSjCtkyYCiIJOwva0CS/gHiVdYd1slBQwD8WZieeB9Rnjlkpg
uTRqKZun3+6DzQp03hD+wgm41VV0vlQJYWR0q37tGAFcE0VMSA9s/y0HurHGljtF
4rUMNM+Hv9Cb/7Jb9p6FAogdJ6B3JeSCdft5MI3koqhDjrUE/pfRY9Fhrv67jNj4
i3sw16kbY8GcaqtKQyVs7OD9jlG5BwG56yWgW3miEp6IbWp5DwgmEn+1fH/908WR
DYY8QK+YRXyD3F55mOHZBoQnfajqlvBOS23Q0/NeeLIANi1Xla+UDucGnC571Moe
960BywH7InV6lPLPky1z51aJie5E+Nwyj0x7tagBI9ao5LAd1S9M4P6u36jJf5Qq
nLZ2McROtSuSfxhZjUtMEWzFaJwpYqoIAj/6UHrb178hskuatjvMqdz2Kn5X3vy8
KnWFLmAy85mWZ5Y8UCTSPWjptgQ6K11h25bJbiiksENwa1hTlHD8xTNY2c4kIu8E
eR3A1mn7kY4uV+SPNbp2Ub0cNobh4SVtfCRVBT2Ya2P6wb9hwZsH9m9BEG0bzbox
Re5bC5L7HM3g0+UQRMOVNgV2dTQ/20PdHyas+EGc0pBipE/9ulYyaNz++9KBYxOD
T/rXAl15MBOuOKojBhpMpKjAErlEtXEPrb3F/x2twJUoCWbwYENvPtaNh9d+chFR
9QvKUpSynKKxCASLbSdVdcZaHTVV94uBCrBXyMkkcMQHKGrZjvL1NLeVQy2qu1pj
2ILT10f78fdwhfzp1oal621UKGRs5Z1ux1u/89AUBthYeZLWQZ9ak6rTYpbNYF6T
MhW8dp7YeNz9CFSmrIWFFn86BXJhK7rty/QPhvHY+wSsG7RBukV7Y2hk1oqDcb0y
gneNGsxG4GVOTI1Xb/G848u8kiJiyjoA52XiT+wE6X2JGCRrECbvZA+lZT+ZeGqQ
ngwwKp70ENcucsE/k6SyA3TcJPCLwNt79Ii360uysKrQcrnQ4pHH8mAYG0u6FZLa
IeApSH4x1pdymOBIfjpixDtXo3SnWFQmNCzBHPdADvNMpTBiqlcrRgL8Ds8p1eaH
4rDLSBwRx7qnyVA33jcuPVILSW1b8SpSdJuViKZmGUe9q34HSuafCuhzO31I2/45
KDNmhwSn36jgb/gqfR2xSWmWF4hfBdlTCIveNPIDFBv9MQuSXw9k8bmcEQOK5jTV
QsQfh7AHztznesCvCE+3cTC868ulkeR4uEHY32sjy+3h7rszqTBBN7EbWHU/EOM+
0ojdgqDFXMt04AOEcXUCYtDQunNssiJT5wAmMztCqxyh2mHIjvMMMc+nIhZj0R5p
xQ24bk7h8FJ8oyJXtSfUhKNlrK90YEvPsG8tCioyFASByX4Tajnyn6jlZDBFSyK9
PHWbf1es/qUAi7OrVI86q1/SanUcyoQEpBCWCRQUtpfmzuhjD2wvuOKY3VzVIc7Y
e6svbtBMhbjokO40g/j02CiRhT+heDYvBKmiPirIOe7d/9CiSViF1NFtLnp2oxvV
VA65L/bFNeyaWgENqp+cGlvTNkBigQm2YjVEWrUDShAg2YCpkYo6B24GFiwu08Xd
pAQtbSRuQvQLlVHAEidTZInH8nsedq3/8GE217HprFxj+asycGoJgIGKLPrfn9Ar
Bj6eq9nSKfz/m4rRUEuPo8mSeyX6O6UhbyJjRnIARt4WPHPYfISXL/+uzDIWwYyg
4zQjU9vcNh0O5aX5Fub0v/W3mqX1gfYfOahIjWlRwgz0zFConAeVWyvh8hUln1cj
55Fb5sZIQA8bLaRC6L/AqrCHgNuP2cZmCovMaVw2D04lNGEmyLLBK2pIkiB3lEzG
F90mEpKOb2jF7JCFmq68tEuKiAa3ZSc+RuvTDCEC0yjE06dz/enCpSM/9EommWVB
KlYO9wAdOeMbu0N0w/upkXHlRazCqyl1Y+k/Z+7FqzJOqzOLaH0dHEyhFltoRsTD
4AWDI+OHIk+41mh2S2bf/Ipx6k3CiP43BYx2RWVYwJdWuXe8eoLk5dvsEA9Tk/+O
9kCinJuWdMfNBivUKyXo0X9Rwut90eQYy1okLMqGhKto249pKkR/IqgtmjDPruHq
ScP4BF1XAZnPIE/ooZ0JmDTBP9v5Eil6qOpw/S32w2TdG0T76c1GdwHCn7TvjEYd
h/ZXQnwO1E9HQTCu+QwvS3QkNeFiXQp204Kasm3rAkn91jadkl0gEWr9LpuVVLUa
ehR100Ja9SnOGjWaPKuRQgOTwBx8MII5YVIhRNb3YDqYAi7Vs/lOLOTAxnmapN/l
ZIRXFF66qNd6Va7pKARMd9F60YsuIn2nFGTKSLRH3KupXnwAMJGYcpsrd4Alk+x0
6QGoD1eklPparQf8hsHwBEwyAPWgdGvs9K+fXry8h0FPTa+wUT37C1azj4OdEqnH
3YkJWBoI1SU7ZNv/cS1kPV1Ij4xYbOy/VbzyyoBgqPXPpimD7SSkucw745dnryJ+
lDmswUTGq5f7r6P1gWQqJeMuM8h60kZQoX9vBToXIYQ+6tmnLe1KJXun3oTwinLp
/5GOrDJu4w0UXqpi5OG7aZuaeBI2jaDMei0hw0heNMMhgGbNTdUxAXOTroNvIuj5
MYmCmE9HVbrt30YGZDGATMy0DF9IU5AwBkvjZyM4Kl4w/D+43YLK+d/uQ9aQrDCH
w9dX874Y6PVe7TBQEmQxTLTJmVbsD6V8FmsD39Sspgg6o3+W7OU7er0O4Q6uEi8c
mB3sWwi9ibY8XqYibpgcWdUGbHOF51p+GdwIBtlH+uGrEVU2LwrAsgI/OqjeMxLO
rUxiOpZLcxiGTC7P8OaX4fyyrUpGrhIYugPI249xKXuG+z1uT+3H0QM4gLOODxh1
fwUAjsr6sVvhuGZFleNKvcFIYlTgbQDiN4qKwDrO2x92mVjjYfRhANQrs3ho+2T5
ybhOYV92JErVGvZsnDJgaZTOW5umoXAb/oZJC8GhDci1z2vsedDZYFyU2yTTHlM8
G4ncD5LuvCthg2r0pmUTipCBx+uHyRTcMqfc9WOOQpUFzZBKZN1CEiaAiCF/0YX9
Qqpet62QXxGVAIduFz4Gn/t3jbScrBqQIbLEJIWgS3FchYhQJz2Y3OTUCSpfKLpE
IFNuGhVd3q1lf+Ez9pe6vkMaLNKRyZsY8Wmpvgi6CS+sQ645eI0UPJ7ACAMs4ZP8
6UkBQ+6K8mbUDZJAj3V0PzXKKT5VPyAIkWqTF/BzK1HKQEVbVGhk04ja1BqJ2B3f
2JHi9DEXaK+JIEe5Pb3cCalekp/2RE+ddxxpBjo1NTyNSSKcjvUHPuFarWUd5y+3
Fn1IT4O6kmLyjePiYixhnW7eW0wgPlTRm4j1v8vtbJZanvghgbpY0lXCp/Dcr/5s
v6BJ6udEtuGEaY4iU0MZ7X9nz7v/IYYXllmSNN6ocdcl5dneng5NONhqzLSkhnKx
g1X/M716ZV/ZjeDD9zsjKiYYFqlDbTDyb1nQBscAgK3fxJdjbxNKOEQTysHyGnMd
jpXGyDD+D9lfjQz5kOHCREx+mw6PA7ONN3G2vjMcffgI7sVl52CHHy/X8mJZndin
B/9eCAEyRB2B9XYiBZFEUETLiJuz3YQW6NAKaYJocbHWXlunGaPLnxnETvzP46i4
U/r1UgHcg+B8I2wj5ArZ+F9NOhbZG9uDLo43/b5SWvXm7WPiJR2+djdztvv9ZkaH
60EY6kAHSxhKCRModRXYGzpDML29qM4NOtmRUn60wEbabjD+yyXlx/8WOzku20V8
gSirP1A5rygtAjcSMikfLyPaJLHGNrqBZW1fU6iNHYO1a5SZVQ3uxGklbIwv6u0h
8arQRW7JQ2alaHRYuk39nbLzSIdHW/afioT7ZRWPJvwQ9WJnWrdXc19qzI3BHcpa
aLeE3oqiPlXI+aAJAn4gW8XzsQDEuaXNF2nRQwp//gFackHo7wXJ5uDLBIYc7OeL
ZVjKJTLzR//6R2reocpw6PP3wXAIuOojr/khqpIjyqmWBCXetV+tFPsxMRUHrKQO
toKx1RA/SMIUMQIqGIDHVyvWRO4W241+4FOYWgvgndWe4MCK8sp+ad5U+koGkf44
K/Qlk11Rz7KukqIU45XSclN5QVYgC4Y4MHsUqG2NdBBOwPDbPaXkaWBVrUcTgmmy
hRN7h0tYGbtPOj685U/IBMk2rrOUoKdJ167hrluDoxYHB3DFTz8cFk3OelAu56tC
dsX3bt3GDuQ+VfnXV4sWcPzPw1oMkuwlxgoOcI0/WzM43fJlKt+EBNDY+krdzK6U
pWLacLU8Q5hjbyzeTdjtXH/xX4FYu8V3rtXWlBrr3FmwhOOGjQo7+i6kU9s3tqXO
bQwre/bR5NqBn4G59dW3aW85KvgBJCvdJijWe/r5cDkjWkyI3VXSYIIyrdOiNN9b
XTh3Mk1odSBdaY2af7Qr9U6riJ+oa0Jqq0nXqH2dGnJX/vfW1mFQTJ8gjBkTDDLL
Yd0galXx6ejQbvarZfwKGyAuVSKISNHgk+Zo1GisvVvSWC2Bsv5QxLk484067X47
u0M1qkI7v77lW/DOeL9ze0n37c79flwa+OlBMOkvEHkG/zh4ngzQAkK2M5zXV0RY
B9sjTirdHgkowQ/Zet/QxW4A+WZL+vbVrF5Z61S0+dA1W1kltsYEKDPhClMzDnAe
LQqd0EVXx+cjT+IkdHJafSEOGES3OUzqn1MNIgS9l/4fc1t5y2qLtd6+3HpU15lx
QXkdHVMVQvb2g1IA1FiHpkXe4lMoRw5ZSkUi6AW8Bodj63BV95pF/K66f6you2FA
5VwFu2iGtqtqM/j40UEC47t99Mn4yjSnHeCZK74QReT4IHlWVYv/2gfhujQITJa0
5pnd3kR5EHhoNwhucP650WFX7TCiZ7Gh/JsD4S8BsVrMxlYjEXf8EnbUtxxDJNHT
NJRMpBIT+qWgGnhSOSeZy5nSN/xeY2IlHkYbaL9jeHUDvy7H1glRLdEta6ana8eR
b6izboa+zQt++bkaub/8sXPG3szVWcjzS1tNGyXTV/5qGB0Q3bGGxiIqWbT7htYd
ibx04IKFFeG6iSPUd9HpLyiaVE1JgN+IcO4w7ws2kpyHa2xFr6ChAO5InyC1lB5s
glBGcnGGs5De12fs+bq4188jx7r4iZPH2azYzeLiQAkhcDEWBz5HwNyBPefD+PM5
GZ80+IY3fRv9Lerxf9y5QbmLq02nbUNOFHFtnDv8VGA/zNdpLYNaBHoxWQswrx2e
vScGS0HuU8Ky2dQ1/sXQgDdg+kJY6gqTkA4a3DrT+Q4i85rehbnHZSdpGrSZIILy
Z04BRz3bJ/IScskF7ZjrDacu3c0tJm+DwDE2QnZunTUgluq4ENZGqpV4S4JUCZ/e
76UnPaPgsnNdh6OIjq7WSRZJ52xGWXZGRGuZmXYqDWe7rXXDWJF4vSt8pw/16adW
MPsszlWltWAhd/Qx3FT7VBeGj4DZZewlUeOMVxBCotdGC3ojydDfx+0dMBrG+hAV
o8Hms9b4OC7qAZlNNqodtTmIEmqz9UmnhXvgFjpielG8vnrJl/i1lNR56EPeAH72
XCA/wOxXkO21Xyt+dd1pW553azNruGC+9El0ocSjXjZBxGv/vI9HjbX1zNRYZyoD
opuEUS+WogQe3Xbmc7oCeBpfKzf7QLOB7cSeFXd1aWHZm3DmbrRXqe/XJqWy9OJa
WGYMSnppDbiHNojZwV/9xvOuvtvhm49T5BYa4GNKrvSXJ5XrKeB2ylWK5Ib+snaV
LJW7UrNDAPkshXBisdHAwZRk7Yn9GKsqOiphJticTMqGL61ueNRJLYHyaRxgpa5r
qT1e1u3+wkxmN1sicD2vd7KurW1p+lasxHW3e3xJmsIACpb3sbeRdOorwbIQ8Mmv
gAoBqs3+JQePoyg0qrZyUpaq4a3aeTlQ9alb/53+DjadcfUKktl7zWcQ/HE2cB+g
FhiFZsJWmN/0/26onb5hH6k207uFfOLQ+nAeSdbWc4z9kfToWE67efPI54Wz83mC
+BW4UEeMuioZIVp5EHC8j5P10ZpC/O7iQLb/trpB04CU/kAWGmS3Z8j82cmvBR04
e3w5Wt7g6MPp/c2bGnD4DiiCzbYW3xdxyw32M8/8R/ErOGm10r/95jlPZPsn45To
A5bjts90eaXiQFrG6i7BtFK3tTBjnhROg6fBBVkqf/fp4uSpMW9tl9kpK83U4xjC
ooM4BryPQCYbRPxjKXO93UYyo3abTH2HdYbq//KmWCCkoSlynwXqr+PRQuIUmKyG
M9eAxJmEAvoOrBz1aRo9HUVIEkNpjcGp19uun1F1GbfKMYLeqIVG9yqjN92Hs6rx
UXB0Uz/E4dRDeFQBmfawUNQIOz5e42mggLzCAM4E+Te3Ij5UH3okzmmvujzmPhZs
V7q1mjyFtS3yVxBlss3aaGxtNzpRrEedFvyOxcrEYWlOtqmAJ1pDRuDOUtEgKZHn
tBghk9ZR5k17Aq3FVs79eGAgwgFKeBuK5Ec//lacc8pWOKdgI9x0QEzWSs9vlFWx
P/vsi3OkMhQgT0aKrN/KbMd+qGQjlZ3TuU9TXuQwyw7iyg0Ba7/TfsmkxKV/NXir
R41R0kLxt7Cb1WG46yfkuNUWGcmcQ2Q1dek7GPiCwLMtSXnDyinzExDde3I5jdbI
W+Qk2LBVpcdnagQigw4D7HlaZrlkMx86bi03nwlBYFLQGZmyZtAP+c6PV3yZPNCI
ogKowGdxz7LgkgdhH0psB5opzaqF/C9D+tf1xM49nLg0zoqJvurNryC90EcZRY+q
9byCwS32vfWZgGxqFAr81pf0b497HCbjOTQSg3wAHznta+OnVCNYHCfLjamMhu06
P+Zp1L4XYG71HsgLJ2Qx131pJ34u7ABjGxlw9icprXFQxHkjbXxslEU/FQHBd35S
8ii5C2hSp1oVJNTFGwZy5+38zeXM7dNeR5ZyNYf8nymYGO9vl5X11cEOyPsq7PgG
/8CF6Gwu5KRCQxk/11CzwDxYz2Dw0AofizMXymprFbhbBPyFFSieRS59dQ/3xom1
B3nL9ByLosvJE9qSMXsNK9HdEVEyN5weBL9LzXA1mZsjCm3CY39xRb44vcviRjDs
17m1wfZX/BMcis4fkqCWqKaBcpO7aV5tOpfxvxYifK2zes9vBUK8JsnnK8shPzut
y/NgcU8UA9Qz1xVuwIMXbpX1I2F07UvXJJq+RNR7zKmjQ1Hv0wUqNcJrodfiTHnT
Z+/4Kv+KXARhv+wTXLg66bQHh5+2s0nT/9wmrC6CZDmfPm+hw27Hbq7wxg0mEEEb
qOWqKtNOf/u+diRGP+GnINe9v1VHlPY7q2vS4E9E5IxamgrkFspQP057SOJSuiYh
4qAmtvtvAeRkBS+A/4Sh0+RQN0gxqzCRgOp4FKJqB+qjas5z6Tfu4TMIj4zIsdWR
G7+9n5Wbxer87XO4d8f/E2PYKetNvFWn8cMbnFNms81+aajqpDgV8qhvcabPOQUO
JrOmXXZYId0FP3yYASe6BWuw8DZxQ+H3Hxo+471PI0BJ18AfsFhE06jAMZ7uy+8F
G/43Gc+71P0LzS9oe8JsE6hBElRuqp4d9Cp0T8x/fnqo8oK3D2ByBV0MyzEbRIrU
4ZTAD9775jL9Dhc6x1ise/qG3d/Z7jkX6FhOpSVruG1r7wLznEPLDpRPBuNAmn4O
rZcnDUhZTkREaDEt7wFitcr3+jmhGmHgNW9bQfN6p13itgTlqBUj+4DgFKgLLVLM
ZOsvk0qEc05ZtctHn6rd08Hpai2FzCJDzmpYZA6pqJrB1tIX/xLDeO3DufSBVRvR
evNGaRmaGT2cZx5vGot5QQ/ZlawdmpwVBB+xqQ4/TgS5MXOUwgd12nT/eGRBVZxP
XvOC/kHE+9JM4V5j0BvInp6pZ/FIUrF/LUUrPfy82VStWBpFKku7360IVnzNDkVB
SUOxYbbnQ4F+6zyxLXa5rXJXySEQr3goPKt6lWhesDUdYGCrChgtx5bZW3PX+PtM
IuB/hYfw6TVZ8xbYoiJn8n7316lQoT2Vve99OQbFZY0yI8d4Q78Iaxl/G3dzfTob
TJ6n5E3sKVJOYyXJk4eGegWy+2ESs02evqr8uinE6mZ0/xaEFOnXoVjNE+40aiJM
S1DsG0Lrb3E+c2g+vOxbx4g+X8VdqN4Lx4z5GWZsp0qYvTm6+9VxkFOzHOqlVBjH
leJKiEeX7SREg2KIKKu1DqQIrFiDgYt9062QIrD1AO9zVjjLLKHKi+UBF+hsRcKO
QJgvH1sJfEaN0iD46f3F42qZMJjsH5X4dgTJQZC1vQmxjobGAo91rtcYqzp6NYWt
wy7A9Tiw45kpt9ortGjWMAXYixKJSKgGa82U67Gim1/ga7ryc4UekO9BO9z230iQ
r+LeBfLdTQvqeX+Z+rApR+qsxld5T/ThLgH97EfOjDMvecZeq/j5MT7aqgKghbtx
Qr06JA7LJ6FVygmuA7MBHVLNMa/vtbe12sPsjBIstEycCiXHBLWg2LRerJazttXj
baIVhYf/TyxteQh5gRVjq9KY2K76Kys0cHPNkDp0NS1t9X/wlbEGLHK/vXJ7anAg
PkI06NM8ev9GeDUtHn65/RCvD2OxTIyPObxntPqBb/8k8pI2g5ps573yCZyOc8EZ
MFHiEB5lzso+xbOdOko4oshaeF4jouRZ1haNoCH3bOp8aE9Eg8h3PPSQHaMxNjO9
ixiF/j4l8eVa02dbPyt8Y4wKkvYfIBtgbjYKtbGxtW+Fo/DoJ89U/mJGwXmtKMEP
aKgOTR01sw2irycp/6/U4ya7s5pJA8XlXhpD0rAC+ARjXLv2AGvzJu/lT1MKqyIH
yzzeoTs2GKidRVpPoqu2wk6v+PQwZpE1jhvbNISTKD8FhiQtaaMUZWZtKMhjbeRR
SEv0dfXVmjmU2+rinTQuQpL30aaIL6fz/2yRA27S523xCz/NcwMnIiDnrtBGKXEw
2PLsii9ohiSL3E5zzvxnzLGRm3KXNs8+HRLnylyjbEzOv3PiTr6mUCH1xVWmRfU5
Z1ZLLuIxbyDl6xAg8uj5X9zS5/05NnA4Q9cATqMHJ9ktMzAcL3YFuhXSVKz4heF+
cnm09t0MYUq/Yj8udEkn13hpjIgUcRgcnMg3V7lVEpVRzO77YZ1fuJw1yp/brYGN
PNlFz7QEoXP+pe7pPW0aEcGmVbacmB93nfzEJRZNn4fvOHOkeddAUgARQIUulHci
wK/rOW+HPANoJ80z1XVaZ3Y+BGjAxljfCKxdaEXuuf6aDakjCagjkKeCI9x2pdyG
4o7njTRS8GQ4nFpVZwS0P/fv9sPcydNU4+WovZXtDICMwgeFpUZIV9OrCb86jjZf
ypWYi5oXVHt/l52+os6WZ63LMYqen6Lv9ye09EQpbzOwEGIb++iNifF/Jt7nHALI
9eAAirbBqtG6DrqPMATQTY9ZV+htFOYjODvdTeQGJBScpGQTYg0bZKKKRnUqEj2P
ZMo+PL062bIxiH4bGZgn8dIAijfabf78pP4JaXcxBPtxc5nwkxVKyoSqJibTB4zE
CpMDzrle3pVDQ0S2jCJRublgV5uwBGFkhVX2mxye7Fj+rkZDFSVE2VxuKc8cx58W
/C5lejQMbkWPgXB5gAVtLyApd7peURjS+lkVK1fG1Mo10xu2yOln5l2yKmamti+X
sM3FMCD3Pzg1Tm9vQzu8osNr6HSAUrnC8VzAs1V16Re8fVIe82f+3UJNcfVED15h
YN83KYZXBVau1STYdikt9t+DAFm/f9Sf0n8NlI+7gy0ewmVlDYAtTujDYHZIchfw
EBD38pA8aVFqzu2LtRW6iyAPjQTRvCXdqMWVVeuA+MixrpZ7e47uhN7DwyrsM6eU
Vrnrm7+ElVyGCF5FLOptRVJpa9EU13CxPK9r1qokWWLiqe3DnjOiXUeTXFYgOa3H
D5kGKlSK4GShjeT3rG95yuS2N9Duaa5a372ApPCrOEfxwDb2d23rAov+MLff+a5g
LVLMBTE5WnU1EBS6c9/0d8nUTzuC7Nu5J7TGw+mrJCF8hEAmTdUqyRTizW6yxtsW
kGlllmz+eXAuwMpHxMMkiV3SP7N0vLxwsiTG24OAWhRvDb5WxfK+Ck39LJW2s2ve
RYN+wexRacAU5imHYcw4V2eipC25sTQNaz/BFyOdZKIDJFd5gd2UQHMNKSHvO+Zw
Ptxt999K6doNva84GVk5d8d7XpbZx7S8Mg5fThcsNWuPB12e/S+n/dWk9MCs+KgU
0pRFoGi7FeqD5eCWUX7PNuBF8zUJM7+588ynsprtwzuyZAhtGmaGsq5b8kh7YcjG
D4pO7fFMJhEvwegSWEctUcr7StGooExYXXaG4/3B4kCVpzBDg5ycH5Gaeyph3J8k
GNoQJX4FpMt9dsL2JG5h0xeRglFhqpdcC57qyIRC/YX/EQ4/NZhPpC/YThQi+wuT
G9uMVe48lqAD3mdkiTIkNQGc7TQ+WO+byKlABAgr0eCp6iWLGwNGp9Gcqk/B4Xhu
1H0mpk+M3NqUd//ijItpMTBzpiEpoxmMpIzZWA6xaYckHDg5SksjJ7UVInelXE+G
qjOqe5X35QdDRr+R/cDkYHMfFYIRnvxXBteN8PRrCVhhiwwMx6UXoWNtYMj1I3AL
4hX3NdDG7lHb7jsNjMUf6Y68aG1JrXwPACIpAsTwUjwG6yQ4XC4y7+BmbA4fZ4Co
ytVX/JgOY+6L6klP9qxJtVwcO6J5h+9jK7yxzEMgefc6kE89BAxbKZlvZ3Y4XF+f
qYYJf4j/qSko8KcH7CFz9GgVB0bpm9XZfbZ1II0jDvCE48X05Covq49yicX1GZ8B
qk80K/tXwVuwVkw5XzRe3xexlahCWmj+VDChs8CVeQjcq5dJRnEXiDPmyZ1cg5bW
+l/D5EaD++chI1gTV8woOSIRO4oEeUGkYvee9jIQhqDSaQAcHx2tMULz1M6vyVGe
N4y0fVhyzdae/KtnnjWV2YbCQKsjr3qS1ZozzSg0Ma/spE5u8uMXNkRsc9ifjRrs
AFO9C7wInEDvtv5v3nPZu4LKRzR4StTyy5c0iVU52v4Kl1nMPdenNzlAGEQ3wmaC
XqFBABAFZQZYrG5B/3epvt3a87GvDU5sfbPkZviIjYMWZMlmBfPT6wrSTZKx/N/A
KpouiEysq6VGYr2/s0+Lz6vndscesqa1aeQa9HxuSZE9k21EkAjl5xnogPfFZR8K
/BmoqjJDR1AbZBzGONjBA1dxE95Ts2s0zqHQPVqnnGOCx2jlbtkFxilnVT+l+u2k
y220THds+S9efsfFY3OLNNWDD2SG2CzuZTYmGhY+u01ZHXmdOMzGIrLXlEYrrWhI
Sqv35bZFZpfSMFV7Rr2bOA0EyVWim6C8lNUPdNZAkgfCAjIYoMhKvV1J/a57BZMK
OirQcM2B3EjDsCqpuxADLAEpB+6NiH6KnMRIUga0GosTMwP+x5DdiQpxRO4ApNpX
+sg4EXVNR1AHSakgX1q4uFgfSKr5U125iatnBQRlxN9GA5zmBEN+8WSgpvj+sI7u
L3tcOZxwAGD/JiaZBJgt0x/xQa+6drUq7vx89rQVqmTmy5J5O/WOTaGpMEeQz4jh
yGcWJh6EFewPA03dPgiMNu5a4qfIdrGkEDbP/m/4d0S4UPj6p37EHkAyZvTxlg0Y
ugtV5tVhTNBAEIGVR16yPAMAMng3RXBO2bmZiHvIAyHVQa5sgpMypbRaHjTjQyOc
47v8+RUNwK1YvjUMg2UO53rfs2AUfsPagj4q9Jz48vzhq0zjpU892S8KgQhOqE7q
CnFto8awohMNzgeCDEOX5oYvaJRG9TmNMdjK4PG0ilFq0sXizCmhb1NjZKwbb/oa
N2UY0qQWRWVQQBl2AgHPsDpETNfIpfv2MLqdRyy+dczEa8xUSHcQTrtsB7CYx0Js
QUjRpZxvqwVym43TPwOPBufSC9r1fy0cqAf3usnsdvPtsB2jm4iVLUC5UwUVcloQ
1FXw85YYJp0Ms0TyctFjeJ/oIXSczJK2Em3PYbhD+vN98RgioJXlkgdGlrJafXBI
Wwh1d8C0EDY3hO+rLdR5YwGc9e2wHRJDiDEndZ/JQEOK6Cawh6n9uGFlNL7mmTvD
lXf7XW9Y5MYxhDcrUKKVXELHq0HqJ8EdPd2Ka/yIhTG7vZZI6zN21YTrOuNIH+V9
K00snxlaZgcn/2vUFg849p3l0DC0b/V5R4ammItUoS9JaZmksay01Hfn+dy7Enuk
cVNZTxxJ3RsFwzGDU1vgSZIpLF8Pqn1RqXC78jyT2dstii//ISrmligb3wmGEybh
Zn8se6kdPd4olKFq5RT1kxTuC4paMpzuGZ8/ybWvMw7YspCOobVR5kRyRhvH0xv8
vLxVBDDdF44uAHD+axwBnBKQwZvJUs1r5e6pTfkwOpBCT4XgosMOPMVJs/HNHGRV
dE5eP59jSMjg0gLFbm3+M3qyUpf48rBopttJlbgig8bhyLNzxOvlN+fST9+KcCQ6
JNPQPeAzncn+YAkypc7oFu7rxLorMQDfzPDRqOeD3/JMKxaqbOOl43biTU9RbqWs
G3s3SPHSvXyI21zcXNSS0HGdZz0cMXUu8FNSi9wHub+MYLLaUfYKvUcHkimiBI8X
ViPvHsGmlNIJ2aZS6qSn1ICo2oNlIDs/+GDkAl3Oki/YJ0nI41CEHQgpJnfh9mwA
p4ktqTrgCRhlSdc43Z0sgwDTdkv4Hno2PuXUqrTz/ZfBRAIf4eXFERw2hQxpCuWc
ChcldVOTWSZdQLb0zxW1ztJNUfxPyfTHEBbEORKwLk2EhDG8sJ2HLHYpA3mB0RfH
ERmpIvpT8Pt3kKxtdXKC5uRH7ZVllzbaw7YjMzAdWM9p1WmTG7egDnIanfq69Gt5
kjCNn0EBRxQQJ9knHuj0S53OD4rzGbR3iPI5VqPVxM9ZN6u0Ntmti49hgbJzeTiY
qVp/MudloLYAv/MPEABV8Tp9OaMQlyjKm9f6c1rVVvbVuIPHsSyfC5c0z0kxAKE6
7+bSjDQnZO+PenbqzvWFv2vouoSp4UcrCbPsAGlhwy0JuuT9aTKNyCM3m80c4dBz
mzL2jQXs/S5vAC3E0txIuM2/wjQBEW3mvSgsqO583/ML1xoqmrd/sJyhfsZLWEc4
OfWuK6Bn6v+aJliu8ZRJLbkGKNnnGSR4AaSDGqaA3H3/cAaAgHVg4b3ipx8soJQ0
veqqh/6rO1cH5+9V6XzBvvPCxxmKOtrpqn+vuVt1mYhUU4fEAwzYyX/h0Gt9RA+x
vNXmA5EnYuaQVODOT5kVgXiVn8TgFZzZ1aD5YR4ZIjY5trf36TsiDMQkbgJoWAaM
CGMtAGeG/bIhIxGq9Bg4xpS/JagMalnVvyCKTDbVOzHXPyvMYV1YFO4NY2GyEYss
LzHfKkcR45WrektcRlmVBbmVxog6EM81bcQGGwZ18OwZQ4QqL7LGcWKGOgWyBuRu
DCqqVqoqYQbWA1Nf1T9yfeG24XLXqwl5/17GnH4gt+6buUh/vz/m4zGJ4c44I+Uy
brSTqYqBq/Qd9fPZeFNwAHfUXSXc9udfjOVRWQguXxd909tlPHfLcC29GUV+RbuB
Y8Nn+NV26wnRwLv5CwMlhXBwVGr02Rzv4PnZ/VgQu1yrerlDTpRBE1qU1/KQiWbR
y5zueLWE7GHI5jC0mS1km151AHRSzWUptYKQ+hmMdXNRQztzSNP7y2CsmSYGD2Ie
iRY2e3tTn2KUc/r1fzVMVACPf8hZZA+BGSYi6wVf6RtRTCg9JymvBHxYoKnnTtP0
NWaHhgXHfbQ1vynk97zR1KFSWeqcvDVGWIwfJALKJwux8LxwNyLh703E5Rz2L5YJ
5fKQQ8n/Q3ANqDn3IJAmOa/axCl5DRJcFzNkAAyIVKZo7i0DWEvI0+nLNSTMWv7j
GwjBKyForQx3dQ2qrahDjy8yspQpCR29WCHJFkn+VsbAopo1cLh6KVkUwpESa0Es
QgkJ0kq9BqfBmL2DtyFjn9THMbb4ZVihg4rcXyev5BdzxJymR+Zkxs67QtNStu3p
lbDHR7pZazh8jU/qTZfwHPIZMYBbUxCfjI1y0TWbVxVVv23BzPkWpqeldrpjmsP5
TiNsOYcHsxBPDMwnOMkaNs9CkUYQJW3qhzg0p2CCMl55qcNaIbRTk9W+OdRH3S8d
eZ8E3sOIGimC/o6RHAJR4PVMqMMOc69Vyhhv3wuQ4bHhe61frxGPMGMSjQBSqbe9
iL/5I9m91nNfPMX1SPewQb5LSx5QWAU6uBKbBSsi/bR90Z6O6k7oI9KvZ7dDjufT
NU4T7vBt0ECKfg+NB1jzoR/CG7NqNFRkFhHvTE9Om89/8N3fRcGT8Uct5f5HgQX2
+7GHnE4gm8rlgHvDRL812dfwrZe+y0Djx348Gw5PXjQV7ueahoqutrlB5g76CXQF
aeFbNZL6HzeyVcHeLDPCkQtjmHcOhpZxtqLG9kWmZ/SeCjFLnHqoi/pwVkOJ+r1l
pMuFo5hiDtoPsDE+TunCIEQR+D8C0kFaLVbYaA2W6g4hduUNIJzfXKJaByGkuW4F
9qQoL1gmnqciC0RqjQ3BqseJlo5y/FK+f6QW0bxWkBiv7YIUZdNtnYuGoDFlnQhX
4dATpWKf3PBTiq6g+qCYMDjoJABBckPEmHKYbNafLuY5tWRNRK7fAjFxuO7UKVoO
YAgbQYMBZf3JuH4aLkQN1JQcTYoxU1Pd9ELusWywiby/yfjlpBH/L+Q7tGQbK5GR
Uqjcvh2/sbKpU1J2DPoZbZRh1V3lTtPPilKVyoBabhlaAwGp0wImPWNVCGkYT8nI
1BdnwoHp/4PjzGaO4JbkxmOPdEE0sVlIhb3VGbrjGXnkA27Ym4LFlRFzIcLcsbLO
UEcqzSQuYWTYBl99b/jW5l6Nk7Dwge6TZl4aLD+jOpNH6U4ZFLuQkgFzocDJk/4c
5H66wg8jVfwza9fFnL0AvDxBfLZy0rh03TgUpOlBLkw1Vjx0rh0SjnNCrg5IsJPm
KYsFyNsSfH5oe3I025snoxDE9Vl0NrFnHxan/a1ZLPnf4Sv5ybOeJDGTmntgTq4L
QYAqKzgKXLUpIWCqmFDv6luasL/UphqqbkPUd7u/sR7yd35MuX5it6Mctop41X55
y5nq7INpofkKE7/ZNsPL7z2OOyk8QI6+xvimFH43ig/i8Dwx6UmQl6J7bq5gMOQs
VlE+wPEQfNfqljN4WjOfys0cHlLkeocSFBMOhdQMEbkuJwPIdrimIE2WMA7bkUH5
MzM2ZGm56bLUECoJgsF5KoaI7gDF+cogDHxSJa5OE+Pk6CMTD/lt5IpWjkLPYb2+
YdjmWVwHo/d90/M+1P0O29dNdDNuch3eThEVWITeJ52VvW8uvzmPilrNcPKU4A7y
vZ0aTmjxLYriIUBzN6c/mSBd5AhdnNRO5cCsrVvsZF4seEck0BGJlooHc6RGNO23
n6loiuPm4UBTRdXcISC+Ojm+PiDtcjqvsdFkQyTlyv3RCQV4Jz7+DewY6d/UbODo
cBsyaL8yzlKrtLbqKEQc7mwyj9GJwEyHK+6Jvh0x5IHos9pH7s5gq8RcxdqPH80u
l80/+6KzghWEXkXocRX6HWr+dLucg+hJDCgjJCK9eLXBMSujPov2g5YAgooYj43V
inWuaqtnEC/IaERGPwS4buO9DC4GZF9HRx3a2eBHTP08+H+1KdOqjSmtzmhlKFbg
/KZqEe+5Wo4pjrzPR2Zzor3ATnjOADJeE0PiIneopn/2mKFvreb5cZit3hsY9gB5
3ttJ/is1Cxmb59RV1M/iizJ+9k/hGNpd6jqCcGqiyJYe5x/03IxniCuM14Xg12qh
deAHMhV4f+JBZZ/WAWGlJMjRJT+MZ4+JuhQGzsiA5bfbbLL7+J/6ssRKkh9cPYsb
cDZtLYRULJ8U3Cx2K5l9ogDLP198twd6LZINJUA0i+fUubW0KqY8Cf/ryO7oWdcY
DU5bfEBM67iiaDV2VIqe0O1FCc+A2WmAoY2g2yCElu07y51B51MKrlcYG5M8OmfJ
aIQlx1MCqbUvH2fFliSz2HHLHw7cfqwCA3NdfIYj6DBpnLmks2aNa3I/B2nuBZk+
SQ2KdJBQ1M3bwGa2mmbSK7NKYUAnVN9lIViRMPpFN5sFBozredLRR+yJ+LLMTfOD
3hOAJdEUto+nmVXhRP0EIbzh5RCF00D130H1/2AmIFFevpx74d3m+f6GHJStK7tS
DENaZetgGhcAX6EjckEGl6NDDXDkz+nXjQXdz0fRDq0DwWkUPvKbVUglVeKQfpR8
/avGFoHsSx9ArgfqQ5bLB7RqiCS+3+YDYynio6Hj4R7TTVXTugAsyMFR/y/e0yPZ
kweNwLrmBJS8PUTjCPvpFQYXK+xGAIQW6JWZj4fvlEdwkM/t5NX1QLTnoz4jWysd
uWgntslxC4Z/fOtWP5t3hTjCq095Zm5k6LDZwSF+/ma18stnygoCdLAjzlii0ONq
MnvkqfBc8cKvFu0bwyscyGLLH8Q2ydytYTLkZQP/s3ehUJfDmcyqN9nwj+gsz/u8
3YXLc5TQL9AbYQb2+tTSkwZF6BY7ToZmdH1EFgcGr0qTe0OPaTtvfwJY/HP94FQd
+us4MlTCr8xd3oj65ECW+Lw3UlsC0qBW4cg4AXy0EfPAmoq5bd6mt/TJX1bGKHcM
Ynwv6yqvLfyDhqdXREPDDwMrblNPl7SuneNdGvFScgXaCyke9TDdAj+O+cM9kxiM
quYQ1WkgRXrg+QPmgHa4sNThrxTl7PA6G8tkcKNYKp11jPvwjMbAYazHcTKPTNPZ
5/BLCzOShg9sOrjDhpeDexxlDE2FfwNb22PT01qP/wktPZx/xgcNygmsytRBEkjk
U2puPmeP/bHu4dhclYEsVWnhJJZrnc19hRMU5ulnxCasUXoXXw7EWbshBuGeU/Ma
R5Zg8XJ7q7gJHnGkncnRBJwkc8mRMcWFma7GlB9zSaC4lSxz3kEJhEHXV1lOfMRj
kR2Vhl+h3RR2bxxFBIPzfhoJfCr4uVbuHzVOX0zRVv7ij9bSNboVISL8jGUavLDF
n1+IwhTwPa50iUMSn8jNZnIAnRxv4tA+2jSYNEnltNhjG9RwfRHcwc9yGnNDJEB7
ewHakt5Wvgd/H5lWiZzgmKeJHmdHfaI5HAXtZfwDhuKX87rmFyxF1lmmIi7lhnOY
esh8GurzFJIcZ8RP1wS3K/kRW0I1lCHggLa/cRL4oCv/lS24+l04PZnn/2PRdNrP
3cK9RVUpnuPEYKpMCJKJaKAlpfq4uv5krAEMT9bOF5nhFACr2cmaAfBIarmrD5dL
kTWNqXCqMoV49t/2sfbaKOBLr6bN86H8ZNSIG5ZMeVn6s/uhlc7xVJ3YVEGcc7QR
bkAahOe8ST4k1TjPkIqEXbJS2okyK/jNlmDJrv9FRIuGwARR6iTXuV0mhZZCtfcU
8uCORhktwOdFBCN/NptD6L1XTtgkKDHXwUC8CWG6atPxrUqIGTqxZZ+thNc+VgOZ
7XT4I3eCjhyirXBbtfS/fcn4q91ATYIMuNKN6uEeyXdKembtnlJErpF1XQ9TIYJ/
Jvly1XwjpEAWtputRpvO3zDBsTFLGLlYmpJV6PeuNb9wSU9O6H7aNtpkHDzo8wNY
7SlwSfk+S7j4597U2iar5pbYZoSVYXxEXdN4XRYYu5FUdpIDGXZPQ6KJsdShbSaw
m9zsk8Qh14eOoSYaS91VwHessUKjsZpqxB8fQriGXZYIkBdgu5DlboHoTBfDKxUg
EWFjCXVYUKVQ0cnn2q1bJLN2JabFWL5E7VF8VA2qD7qNwJ4QMoUkufytpafeb440
9jZ5xyGnJqlKZfunuF0nzdx5hqq+3BV5ZYvbDWAuyQ0OBalFsUKV8CV91vHGWjKa
MiAHS+fZfGPLlJy6M0+A36hZs+Q5xL9kDQ/Z/8Dne0xv6cr7PCHffOA9RCdP6Bm8
m2ft5HSTT6HAfoun+lluhtDz29+VXSgeV/GKc72TQc/Ogv6qTwpsBkJorB37xidH
S03G2Uh3gIouItbug48rl8EBgR7jypUoKZaHls7pFAGhReUd32S4/7PxYNw3s/55
hAjt5jaItrXOpGol/KMD8TWWgSIQD5KJNXOBCnxuAHe8wLGPtvnstoepLueaZTJC
NXcuZ6MF+GE/LuS6Uqf7Hw4q4KtrKsAhIaH9Fi0yieAjMBSk5MHnFQBAvVqv7LsF
gX3y0QpoAS0oBEBZv5Og0LCAhtKMcNcqCqjpt3c78yBIK4sI8UPinH/47EAYOmBl
dvxlXK9oJFD8C8zWLTAw+ETv3HmToHRRsT1ujND4QrBrMjWlgF5YC/d0K4nVT9D8
nM8hweTziJwasYdrk9j0hKKtmc35gDKk3p+zg2DTqWI++YO6jwiD1QSHCiZQu4tk
bT/DpcIbFkMalsRvalRBt9AFGz0ZQ/JZG7TMSK9R6JHESRHKO4MFTpS0HSgq5MbD
YHKpohvepAmFITfz+9UPaBPkCYPzs3gLxctg9+sLU0LKjUwONP2gKss2cRbCKLdR
OvsuJnmzwaPvYRQ+nxus7gpTD18dudywLoOMl4gbUqC6xYLG+2eWHc5RDGcY4wwh
hBmg5Mrtj3A7ziaeX44K4zXqpEL72ZXIL33CoJop+wIj9jahTUoIH91hZz6pEvKD
kpfPJmtmA9P9EWzgxFsY6v0L6IGHcZmDSYePgtC7ssxpoW1BF1N3ib4AsEh3pqNI
iNmwVx+WIdhNMKLW3f+B7Vk1jdYRHxfbGN4JsPwOa1VH9HyMHr2V6AT3d15DCa12
2wDb8psF2tWPVYa8hlUVFN7bur4hz66P6hegBnF0ZiESCwSolVPZhpNAMWsqwLkc
jSVE3/M8O53G0y5YFqsusCwG7XbtbxmwhRzrXC6cd9B81lx2m87mOrsSPFABVkHy
FMYfaKN4/1839FLyaKTTu0Y//l6cTXGEUBY8vZI28H961KC5PblyqxLTcauYA+EE
djQUUdc+ibSpuXOCK3OXMUdIjOOJSfa7Xe1YyeraqJkVH1PIoQMo9TTATEEwKyKX
/+NjcQ/ybSclIQVrFHvvVXELXClfU3royyJJYS81Zb/9a6kRwD9YVAXguiggbard
z1saR0tzlq/fGNs61eVlhnGkWsVFkxF5jLiZoqw2ikxkX0hIVM/mD3koUARcPkU8
H2mchOVfxoL24Qb+k+dJ3jblmJbDvFozUWRUbsteXeR3IKP2Kt9RGC01pV+YO3li
FfZ6FKFvZrzcLWLzY01Sg0GMF+mQ4878OeNpDVeoED/ht4ZKG0BWuCQV9L9250mQ
zNfDNpw+EOlaCNN2Y6F/t1FKUh5p1xvXMUGZNzvX5Od6PNaZNYyNIEr/SguCfYIw
TSiZd6WMURUcnuW5ERtZ4dp2fdymuFz92AXVrLLGcxIdsE0ZsWJrb/+tIFKLucJm
IIo98G1zyqT3dnvkn2AaaIhO9d+uA+TolhB9iEOwU79i3nMXTiWP68GTrlxRKTb5
U4feNmcXu7f1j27fb98TnI9Y75eIQ/6RX2BtW8IBU4T8UOjBewGYXuzVTK5E/lvf
EoEbKHbZr66VJd/BvFTM8Pee9+U4qX7nbDS6rvMcHlXqwAwrF03B3wa0y7/oVVaE
aqLPKAO1jfrSU98Yb41dHWZbPZq2CDuMnDBSgqH1Xqd1Qd7xwCdfNRod6+vAfNyT
pfW4zm4TmuV5L1asB7kWSQI6igyguwTOz+mTcwTu99+RV7wKnPZeb52y1lI1mxex
YMbGo4zVy5ATkyry0wqu8nt+Ei6fQ3jAjm9XwxTVSJlJPxK3DkQRTS3Op+65ueEH
cU1p30P5gN5KyvJdEYwbJMXdmgE91gAXawUwVy6pUsiaRy0bmQRv0XS5KBHfa2od
N55nuFZBIrEwB6ZDcbbbm7C4MyD+ZHrxmVQegyeaa0CjzozBIhVGqK3hi5BF5gaw
zrFfqZQhmDkuEygEUQhhxuhHXitXEhpGRVjNPGOlHME5baqfn+BL3MelKYbydW/n
A75ktF/Xg/RJh9LHqa3d0fQPtxxgupCV5aV4oVpCPG3jjplyLmRuGihd1+X/Bju+
pDmosuhzFFwMNj8mjT0vchtMPpwPo2+qRvMAdXhOEcWy3nKyjcCU+8zqkpL2T6FB
+dAvfF8sDUDPmwo4IJ5Xvn/mBqt+r/B5Nv6RXYh4V9BcLG6AG85VKah8iRElcqx8
vkdZJC5zE9dune4fS9gSlPmlgLLOUbwJgjs07DKf5qrqanjMlMZ/GZMVKg+fS6Mu
Qu7PL0C6rfSBeukFk5+mfLz2+BK9J5seh1NG1lM9BKORlTXW0p+U+IpGzvQ0GxU7
ILxMaZ903qPsAYk8GF0gHU4ny2JfZI8ETgEDjCl3Q92Qfq8OQwvy1FPy+VbJG02C
iCuYAaaOBP26VvFBDbDheS5zkUJIKGCgefd7DGeaTX1usckQdfKRhBg8MV8xCU85
BRZgj/DqH7wYRJD7VZbiFnL9sA/PJ6Sy6vVPf447i8nILWO7TkkJkZ2VZY14bEUn
D42X+bDd17H3xlG+uIQQRa0oio5iyXBhVHwD3E2IcjoS3evh5m4aZ9iW//PpTlxU
UdgOIYnpbvj37CMmu6wNwYBeHw8OSoru9shMPPwpXUFSUiLNxMv9NDnnNSTAMQGn
odTvIanCk1LqAddUkYQGysRiGJCJeuVB1lQiLNqn1tUV8JC9Sbl+R+9KjQ/R4qeB
7MxY1vGiygGzdZX/WUgeIVq3Ls3AkbI6efBQU2xZdY0fXtB+GzJGhMBSXIk3oyqp
ETQ+3qpH9LzmvhM9FSWM2t3JkDyvFB9St5Sb1t2xnGEkNx8yrllffUIm/SYpnvD3
03w4gY5J+5oEOo8VlI1lpiRkchI02PPzAqEw1gO/PWe0QijUsrHnY8SdVm0Jy6Wn
XBRorVcxiO6iu1dbDFkFt+DajEwR0Bommk37lgqgKEzOQETAapxRgRRZ7bDgbdHV
i7tmx+jA9zUfz+B65oCUSZBMddKqxoHVTlImO1wGpr5shmCD8GnLmc9FMrJhjLI7
yH+eJp2jBCJ03NwvXOjvdCSwWf0R7RGrz1o6r8j+QSXeh0F9HYbD7zgJY0fquRXA
yqHkHLKMltse4i881F0quBmuYOOOkloT/FG01iX6xlTJzsz94yHcCPP/rR8QMHwo
2NE7LbM/jm2h5lRmcw+tKl8NpipAXpQoeYFqFMmkzQDZz4rt0OzgGPeGWyu3jxi2
7Ury99Be9LLIJC4k9cLa98W2xFjzUUbNHRFlCJZxONIP0MCyni45ZlHQlb2pVMh/
BMVpxyu9q5PZUZqtrue595lfhsR52ZEoKO/7/ym2PCrVaeIXAQ8zJUNjPT6mj+DD
RedSes1CD6Ytsg0KqjJaVZ5lmXwmzbbHp5nU++DKdJ0H1rajFBp913yBrk1rea/X
6Z9qJhve3I+KKD8t9CxG0LT1wLFqWytCZCohEciRME+dG2sj2kk/PrsD8LZUoOr+
agoF33b+veNqHTqMpZJRKsGRj1MjpM8hZzp4HH/C2AW7hKtUIgAJoEZnM+tTshJv
bYYljayViVHxnNgvcp/+g5B6LEz7F41dWgE6YhdLEYLrCBRC4o0cSDb3NiHn67Yg
THOWZhbMBvtK26HdbXYsNyhmL/YeP4HhI3H8qNa/Afu7vhLSAqYYtpw31vC1Sjkd
G91AzG9jsnxtO9ZJEba8oYs9NDgXr+X3Ln0dkjOKkGnFIneJgR5z7K0bgkuF3Gsg
HVOqzkhpOi1YexHvilsIyYUGAXrSxZt0mVv+JbXC52o2u8HTSq8B9WXaf0gkXXpt
vSlFV+bblFOi2bV1uULOkyS8mrz91mk9yEPYtDpALjkPUWAndvoqBPsqps1QVXSy
TFmOqqpHT3YkGHRR7TWvH0Bj13pGonnRyjVWoJ+dq79T/BzoJdYP4RWztYRqM4k0
1GXAS6Su7NDLjDAkowpPUHJuobZH//TfmxpUv0NHGbg04jXX1RxjykJFtplZa51c
IUQOCA4Wqm6FMtRVd/QvPLQcLfQLBRITWD5lNBnTKsy/LjwdOhOktRqgTPLTVZnQ
szLeHkhuJVTEstYdpllxTemJ8vDe5YLGjgysXqc0naA7T3HOWRcSx7ThwPn9yP1W
ls+cThHUu+xaRlxLegEFtWxhHcHS33ci0/RnuQUTts2kxdjG/qGkIfoqsP+qPVq2
EeF+4jfIxuCVoT8xAAyXSC3miuGNSZGuGvVwFV676AChARZRN3aU76rf4XL7hS35
vS3PPcUXTlVfncx02JP415EdtXaqQKJc0KnnRrlguoXNibGyNlkgIT3S8feLVCr1
/VFRoaryE4fqTU4WQ28YgzFYJNDvJdzRC+68OE6PGzQNFcwdqDmprTYbx3htqxcw
rhR9Jb4zcwwohseBzZmoALe/LY9UUKJ3ywZTkGKIE+Oj4c27W55CzScDT6klgUG6
a9mFDZlT++kHkDbGXvWP8jAUM4Spnb9xsKDKX4rliohZERJc9tHt1UCn5gHZInZE
HeXJCGmv9uCK8Ri+SzlUqVGq52e4jXFZ/h2jt9CgAF0Ey83iTBIh3hez2VAiXN0o
Pfi091O1O4c14oV2LCOtzY65lm1GdPPNlceOqKVsF+CFxca1jph8BrNE2WOt8ZcC
fG3G7/q3+9VwrV4SzAnV+22/6JXQ6KRBrIAaFfKFvkSa5Eo8N9K2QRH3P+5YjPQE
QfYrHsItYYBFQBdorXZK64w0ntvNEZPW0ljfkx5KZ0/PnIIOQW+zbihsxZ6l+moR
yYvcEaVEJl3BuS6d5QtRzOBd3cxZ9OtcZKanUm11hwDF51k6BE6QNY1Ssg8/QWEz
/C8Ia7To1P5PJEge8HAdHYxojcj+jbCRRBps41cXycylEILic0oCQUpdRf1W75nN
Ea4IljCnK+V3HGhjEdwoZAu1J1TzmFvnNYUxfRXI0MvtCha/DvZWB1/8eX9e5cd2
IkSNzMa6VwLgFzV0RyYqzDsWGekqoBMMUoYymiOS301NkGjTo2cmVYwIPeS35w9O
hF+/6HYL+i70lDDNWyDIgSAr1iEAUQuTI6I6VEFLgBDJG2l+/wZr+rktIic3K6uN
Awlp4RFTB92GbSlc0ZtVz9itqb4YAP5dcHWxaHbOeaL3JSgl6FFj1hyDfAHdY7f1
/p+IS5+7ZQrZYhY/teRS4IdvKabIzo7wPkkrj/GLdXHU24AROignQMSaYqr9YDrV
7K2jrW1jC0sIehdqOOmyIlHmpeSzzFTd/GukXxVaV/64KQ1HJOgpRtBODLE737xW
HGaqoKvTxhDNoqT1zwFvByVDg14zfqzUX5DP8UP2HrgSY3Jl4qauNx9IMHUiY02/
TuGdYXKkTmA/6xtPTX5U1bZqR+jG8YWv9q0epr1e5xqtTY1XV4rQ94/tpS1KIn3t
p/aRhU747zydk/D9NFPVL59ERfWfvh5ur9aCMgVItuZ8Vd/leDaVCOsW7J7pojBg
WTtCaxJ7sILiCwtX+8McJ5fk+z/WDpSd6Y+MA2a6C0dfiLIPX0AhKDgVPlJjQDf4
EpWTz6ArcLhShb1VdqAqt65PaM3Y0CMFXKkrcHLq95Vyp2/gVgfL++Mmqy1q+PpS
DpGt6YBZqfZd2UP8aVUihXqfn7bVb/fxnJmKgCmVaWxSrpPGMXzpnS1DeTSR0TmI
3sSgjK3HLH9/B0GdkxBpNTrtc61Jz0wfJ/2/1whs4h6e7XhLD6PP0b2dupc/Dx6a
C1/2UnBghoRNPP8V/nvqhNKxHxOF5ZolTGNsl3gOgKQFEXEwpdaxxOjS1MjCZ+qL
3FigNZXukjmLc2hG9pMwj2nxZcveXxTb1cjyHat1CA7Yt7txT2y0qt4VXOH4U05v
S6tj9SzFEJ/+uct7NwNYvWzLHz6467OcDxCeUutkD3g9qkM94QRuFP1od8Da6Pvf
XLiLGS0sBNsfDZcw7iaOcT5d2Y1u4jyNvXFBsFgOoWew28XRIMA+gdUJHcsZvKno
Dl5Trp5t0x7pvkRotBgbd326vIeEVn4C45qklmZY1ULTAVdBHgTMCX0WB8Pio8Az
qQwSRnZmHyUll+EOTtJ98h1IOSMyBMo1e6aaysLXoxvtzzff5xDbDtOfs6D95Wad
g+f/N0u6yditCsobvlK/hRcSSscHFJBvz2MAxEi0ZTUN/ZfMIUtJeEllrvc7tldt
KWZKUpS5F+LAqxIqoB69ttis7fC/pNI7qHN0DjyYj+WKh1reFr6GEFNIl1gqDnD2
k/z9h4qAFhQ5CbXZlOIvkx/AGDqtqDUL1CfqpnS4mlvu75cGZVNrK/XjC1+c4b2v
m8fTUtUe+Z5lROmKEC2ETi1ExnNWDxHvRxG8ZnRU01Aj8fm26K0ZJG+H2luzmR2p
O5QGSuCNmjgJJbsMYObdcUQ92rNaWZJ+9hhxxMzMb02MtKz2Jaqqxz7YNRtHE79e
q4TlgwxSiSFiOra9DQUaHH+XgjHSa+EVgCDd2VLT7E/UE19dXNf2FgRVOyzSRUI5
ZmV351Ji3Go/zov0tl4blAgBZyenm8ugoMouoh/2b6l0j40pq645MxO/T1BPEEF+
qzZ6z8pN/9pdttgAQD+0sFDNUX5YetJhftjKq4V2Wf8Q8iBwcDyy9TNdFxTgP2Sz
ZzGc/C+Q3tgaYCxw4pzP578EKeotYMK3DrKXtARpjeyNTnRthsCD8Qkdiz7kVsia
/RPyunxfHvSuoxcgODNW/nt5nFQDTUTYtcSuiN9bBiLlF0/gQw1rMxnDZyg04dl6
WbduRJ3HZpP8uI51eQ8+JkYbbBfaryU2E8IYTzQGojPPbZ6+cAQ1p0biSDdIFK53
sFpoKgJGPXTCtqRIsztcBsV7Mivl+r7m0aUGUbQR9apjgw4LpgUtb+tSxF9+Rdkf
0wjL0RDcSV1NXAZeDInB6sI5ke8V8TLNLMglZ+iOG0AJU3jebXCeoJup+IS7iW1r
01NvviYkqk5//41nTEeDFQ8Dv5kp2PJ8kq1ohPOHLW/OJUisYqCvFqXW5FLE+v8r
40ZwYGdQpWPBv+zr/vHBEGDThogund6wSbXZPLyd0PNZCHRMBC07IzUojgpk/qU2
9KC29/j2jMzS2MiIcg48ojSo/xpJZKWy4yuyMRLo7jSqMbE/H9jPAGa1p2uRc/bw
/pAyZFZzPaGzunikXcDvIQwX0ytF2ZwjYqioOODbDEQz/AHm13FaCLucc9GK6eoL
9K4Fg+rhLfFIN4C9KZiH70M8vgHAdGiFcNz7v4y67kdm+iKgdOVXbDgPxmabg9gh
KFHmQa1+0Tmb2bqx3kD2P22pwd0wz/jUJeBOuDOMRXbj74cJIdlunhcXQlD47oa1
61y+/FGow5arGQLkl4DWrBmJ39qNFzszsSLj13taIE4Q8JZMCIFTxgCa66LhVY9C
2RkVZLITdCX/eY9b+pdVb01fugokwlst3owlrZ2BSV5yfYySFYu/itGzKaTZ11BK
7wRx9dZLyErQlmEryul6imPc3xWtdT36rvFIDx/43j8Gg9XYy/WI5alE/oCgCco1
q7jjY7/+D5tkxoVcO6x0M6bMLEkmdhleupSSQcyPTdMXW68s43oXG0Awa5h1j31v
Lls3yVkzqnlQ06nKsH3RVDJ2NqbgNjYHh2loJcmQB7jeySCZhquRT5vEXMwBmUFU
zfr+KMj3v+RHncE07Ye1hG4h6ILKH6ddKa9gl2OmaF4nP/MomXhwmP24NhOUpJTj
1FBCTxe7D1JONyTlSvS13IvzxD1JxyN0QuLJRpL+LPTtxt5CBaRtejsat95M0QY/
CrzHWWRbUbI1HnNObBO4uhB4RIR4NnRhYpe35yBk8h3JyInV0QHNTx4Dyrc8XecF
hpGFYayW4jovt8u5AvfeWDvZce5hVu5Tg2fQgzikHXA6AxYTyN524lsu3O/PM7h0
i2fE4sBuy5FjJE1OqjFIfinrMIHfREbfA+IYQsHSlqN7eAA0KJTxj9yNAQXuvkaO
Bo0VWtsWiOAGzmAKVbq9v8UcGRSNPdzO51IHUBV05cZ07dyLIUcdVI7JuwM4aXns
U/7n7QgXwLmkVCIcUT6r+r6Sf5OtvLfKfA/OUIPL0SpOzwk29qxGi8clta+5wd+t
4Q29FbQsXiLmh0RURctJ/DpwabEW9on2ZtHlHzzNng5Z7xvHb879J0kBL2NJEVEL
4gTGoxHONR6oT0Sy8gnwNP4qgCEMXJaL0w4H+Ft8+HYADU037A13HVOttFyOBymA
TqDoeHjBXov5DR9AZ6HYHy3C1Lk/eJc9dAiIg8ln/UX8xttVL98bp2D8neXqZemE
TTYsSifcWih0HMqZlpPS0irMP9mVxy9z28NvlC8U82av7f1Y5e7h7dZmsrEiIwNI
Uiw1G+PeWGM4yK+Xhb3CKHJXm5i63Ze9LxJjQ1COPEZkaqXy6b4Lfrm6QHPCeJZW
O+5K7fS+kGT/gBuxvZoGNId1md27mTp0USxmgOD4MjqLrhOfBschgMj8Dt8r2wG5
kelCYjgt/5XZgVr9+CTYA7Aue6kfBN7vPUjugAaS1Da8NFtQLaz+m2jQ2DhI5FaP
zq1anzmnNp3dkGyJmH1xuzn2wZWxGVeKQ+zJHILjrdEzyffsGtfV85CDzawvVN+v
dFKk6vXqDyhPuCxao4dBhvUJ3TxSGdB9rxWyYCmjCtdAvI0BjWTpIOoXa7g6fgay
5JsT8n17IViPOutKOLm0syDmncvhoHbt/yNe9ad2f5XMb09ITSQ2cExOUrA2rf9j
EyOJOX/WeE8UMP4oFfKj8UKErQOMGd/HXv7oF8/he5/GHnLlPISuH0dguofHXLdL
QyLKdW9NaEGYVBpHL1su+/WoxBZhkRc9Mn6OW9BEFgMMVZ+OAiB+/0frgNFB/Ikp
mc762PaZwUt9AU3uJ7g3K/z/Y8U2Chy0DaMG3pk4dbD6R9HwCWmir7bUY1aFNo0r
BXJIy7++crrK/nJ+y8O8Mm/F5Fi36A+M9+7qKxZTUqA/NiQmdE3DR6w49vaVBzuo
G/65gSuAwA0QUFCtgK/K2pG7GfKCtPrdKLpVwm0chaITpKyfU++cryJ6CWoA3wYR
0vkugJJUxb8/IwdnFMM2Zz0Xg8RNJxqfBFKUfW6XI6t84af6BR91XjM/AjQ9dUu1
veHQdY8GMhD0fejkoQYiA5YlmgT4szBvmuBPdVvfJ/1Q9v7iNkfnV0s93nJixR2g
gAHH515XhtN0s672+TWtMmyvSfSFP/IAkmIc86pomLdI5Wq12CnCuTBf5JRdkfo0
BYoRGK+P+oQqPl9rdLd4ODgth/i2CevOYZwzh2y0/mem+V8viw2PjhF4d00QEeYX
gcYsSaa5F12iE1EZsBqItlK0tz9K1OVIqi54j4tMbj03zDW3n0bb2U/t8pc0QoPy
FQv84io4FyKdHdN51l7HwvMGswp0PmFdgl/rT1z04bRknPJt804t6rpHO6RkEkT0
A3nc2ukD3YlPdOGUL5Lfblkp4/RhhXY+/eVciSyJvsJWBp3yDtaIgC5HD2fvYYJN
lf8PCK5iAHvZMNgGwUaB6akWZRSgPOlVVy0YvdZQoNuh0+ku7JbGTeuisqJ6YM9L
wWmrPEqEkMSFnR+ouJYH8O6cPifOQjiXd/wRhUJBQ1DmFlAzny6r7xLBL8mrGjW5
anDC6itcRPyuQDnVvgatNlO3XQGtkMt/a0YsAMiFtcLo1EPH8Z1xm+aoEZVZkO5+
2zJKWP9munhXotSXmAj6Q4LqdEa97Qn3v/mauiDoQcGrJJr2Pb8LolIQ2mZsMlRk
e9pkwbrpKMxQLcD1g2ztiLWH2AZc647paTowuNtKTOBQrP6/kiVV1onkcYQal4x1
NQU9H0kI9J/DYuyHgjBDVoDKidTpl+OOu14O+3xvKo0zfg9cqMwxmAQVSoQIPGrs
n3MP5UmCMvx4OMZ5hugJ00/YIS7zAWLslv+y6/jw2ZElgOol0f4x9VYyufVylL2X
enQiKk9ufUdL3Pcv+X4p7yBA7oZD7fk6uurZ6baIt5RHczAE/6LL6cFSkzUoJROv
vzVd3KLlwLgOXK5zUuOkGP7u5YcE7mxpTUf2RbQubgbxutEJdyiz95wsESYTQWZo
PNR7TA7U+ou2wZ71JmDvJnQE/EKZmP8wrEFTdO34LA7mhVwtxYR1119TBSFPxZz2
2h0UmVfc09R4PLBAYMPTvZPxVLP3DpQ1z1IHx5K9oTv2p0McqANk2ON1K6b2Ue45
tiSVSTZQP2O/GSzlhviDGiobGLCNXcFyHZJ18yNgx7pP3Jqn7PG8CsvMso7blQDR
Dl3426D/MQIROjOEIjIHTUx9MSnf2bPe77gtbmhkCPVyWj+4/cvAGJq7TTf7YqnV
kDR+HPXhKihTh/ZgCbRsl1qsMAT3MYy6TwpR20WUQx8vApFt5LXRNvGqoonNXegc
D+cJ2jzposF2EZxLGtYb+ByHDdEXQSl1EjuUzfwQ+U2UjXOwDq+0Kbc1LIqYD6D5
kFo5Awtz4Qmp8ZHWeW1XsRrxhELRB+17SnH2dc6ouBAr1bMa2pEnst0LdKurB/70
XXy/wEECvo1G5kllz6BG700eX1boULvPN4J/Crw6S8Ac7n7/dGjaYpTr9CJpI74F
70yvVxraJHYd+v08Uq7VRzGObAD+UdOL+wvqmOu4/JToT69eZKy/7+WrA/dDr1sC
9qWdWNYW6r1rsCeCWWu0nJyyH7dDsqP94u+5nAtXpI9usmvVuKyKnNLeIM86H4RV
xKJkOjjp8LfhMJY6AcHsoEkaJcn6c+lR83mZW05ur0i+aPTT0yPClCcK2Rt4WqSR
ZEast944qDjd1qu73Ph5j2h5T/9NBwKLaHtBeFXX+gCRe3RWWDQoKsHGtNnfCPFq
aAJmNvWDp2HOtNbv0HNhU2HfScs1fSnvnfUbmdhruH/KoEtp4czZzG3Rb+ndxE9u
bhCUVg/XKqI53tfmNnG2QOrMSe6j6nO8j5eRuOsjiFVkM/Dt3dZh7PcvlMq8ros3
Chmhym+f01xwz9fl49TH74zyYxAyf2UgC1InBRcTkd/0m/nb0AtKiCApBLUZTat2
g2n0x1k3gCImPhP6s6EzmVOY3hhClANAzfGOh0Dtf49ex3iUrcooER6DSEo4aCCi
EpfHPfqPqcBLgOm+3mVc0b3a461JcsrR1TrnyUKpWzWzXP7s4P0A47GoeA3fVN2b
VOnsqKiGrsCQsmP+a58ymFgZqGbqUXK3uqdOKU95UhtK6hU9c/KokLkgy8SKwQLw
yNOsYUkucSFz7eNUcdRvSexEo8KiNYfKP3E///aLtcSbCqQHNiLYym5+HM5J0Zaa
QH05uIX1jFKboH+wxtTKP4PZbzDzYSDtYK7Nuz4asqCtGWQ1rCKdpmalrkEvn/+f
4kXcdgCQ2yy/2JIENPMhIsxEWpxrER8uWhGPBYW61IyldONMoMaFiSFKvtl4Z7xz
hHfcnkIMinvv7RKZRxQ//Ja2sqSHUDQU4KcNQbjTbvAPBf96/ifgBy1WJsins30G
vNlQszKFYRGo7Zdx/djswrzwW2kGvg3yRdLKBioYr1xvP41M9NYSdX0kl0QNbsZA
m+rC/Xq64nE2Rm7uNLeMD8RsIwUidA1N+G3Fk7xWU8fZQS4tWx/wWzazpjECKmH+
khtscIf3JsKv4K6UPx0kFDtNdmizsEuz+lLkMg2ibtUYhMi7KSA2ooLGV13au6Dr
D9Ywh54gdzojKPr2M4LwGhpXY4Otw8L3zgN0ODp9xLUOHNpFIGSebz9wZqJNh6Ok
y2l+xVksSEOcCdm+zTY0kzqQHz46lUJ+VDHk8njLPxohQI39WHulG+Ag8upcJM6h
h/9b0xxn3+hFnmi2saTMsUGVfuzN1qYvAMcGHQt8VZ3POkoeZ4f3OH7cM/2ABM4m
mswKDvUiUuBBMIe81XYBGa/nl8ML77G5VoKSZH4jOawAi9gFtonw9Qf+pFdnzObH
xHGRCaJhmUEM3E0iTzq7NVRR17hsE54LS5veNMZzzF4WBdA2ukLsHZSFsJk8PHoj
Lk7tjZRM4gI18fITqP+v7Pfuz8+YDheRlxEJS/MSURo/bY4pQES5nF5bRkSqVG++
Y8VnNwqgeSzcHKrTUhZZoiprKmf1gOi3QR2qLKgTWy5gtclmta07UZ4qSaVHfE+w
2umAVFpLRL6O2rtJmTzLahLrjskrfWDOTJfwlsG7FBI8bk/fcEWNfHXVgIOumY49
Xd93foYKCfYeeqm9R87mQKpmKu056hOinHoSNumenHEAGw57SD+f3/eOmX8/Lk4e
Bftrw58ooWt4ZGZITqF4kLpUcTIBIhEks5O786Y9oFqhpRB5XS22xSzXac58tgsK
L1XoD6BkA3En6ubSJ741SBaXa87ttqdVYzsZogA6kDOJC+ZlWU/+fxw7DYq4jJq5
3kOvqiPvmchsQDq4kHizEscuuJpXatxYE1iWMsYkO5sgX66lNukag6lA4DuEcSEp
d2RGdLIjt3PYE3SsztSnxJC5TMxr8V2PgvNSKSP58Nxx00lzKlr/4D8JfNEnsRA5
5+CpdZ2+r6RoRy7O8vmHXx+U1y0q6gUCJwtfkvexf30xw80sFeVyCRkjivjEVi+m
fE0niZ/oAjdZx/bU5RL5ySS56UyTZy30cImvO2jktUAO0sbZ1PWHgWJx+BUNIw8J
3afuQnl0WVcvIARIP1ab97xgnq8EyUkRRsbywbpfwjc0sqCcwno9IPzCm2fuiwcG
5bUHbi6RToJ4spIsWFPn0G2I6WV+um9q9G6/FbQiWo/rF10+aSZ+8dcKwATsuGH9
emvJ7j1jSywZA7lvHF6OuRRnmQq5Q1hLWEqFBNPVFWOFBNrAttU6RHMPTzzZzhhw
iRjYak3XveGgj3eEKhwygGHUrjv9HJdQT9S86wTTuszh2pGezkpbtdfMMEokjfdI
s4DrRCQvYS2Kq51OrSVusEFdqIi8wLUzSesoI/2QleMkZifF14ZRa2p1FUo90bS+
C/ozazJR8U0ZoTAd8EDj1F/JdlVsS6CRyy5Rz/hNnE7Yc/OptAPlU80mE03MJeRU
V43sbx6S6chlAfaUeGDquMs/kAU2C7ebSBvzNb4vqcBOEQ/uonAn7vDaDVRmJQks
WAItFJXOxJlhbJw17gP84X7yQLrWPgyOK95SCKeRFKOShl0eKZSGQD9b+YvemFZ1
qVa+1sIbDFN3EMk3OV61PlxBRCkV6whKjB3NqiYKTjO2WazkNI3z02hfEHDbOzsm
tqQmI158SqBsA5c8aJO5Ep9IcxlB3khv2V9hcSwqhSN8CQOZ2XlGO73k0tecXNEp
jC9jwSvIp0d3+/PQmrzRLzER8DyQvogqToUyN+EWAJZcL/kca/BiDBWDoT+Zj+t3
QkpdnavCFabqhVJ3mZgXARARBn0Y259CnmWsNcxcxFhIQBrZ802hqnsheEIq9ZjH
6czVruZpE0qdzYMjFGmB4v+5G0N9Xp9C1l+XXeBgWn3X6XYQlHOXg/ZYUsuz2Pe5
zPV176ILUwuBlT9FvWSxl+aMSCcKPHKmfzoZ5QnhUsAAYCmdxTsjLLxY5cmaTDIe
cvaxg2wxeDG60n407T3tfMLxnUVUxNtHCt9STDAB9O0RBJXiCbt6mWaqwluo8Ktj
qjBzpAtgTRSAk8QeTgt9nhaYQQKB1jcA3uV34En3fMXTusgV0No6WpYHsflXa/jr
BWheplw75N8UJkF16VERPpPD3ukHITNCGZz1giNBwFcn4VOOD28LWShLM57mKfCw
wGYY5Ku8qsGYWzN+bJBsl+ynFnhqNtlzS9HQmxjwzNyuUt88HLN1yfurbO7Kzqw7
yuyZm98ADjVTsvcw51e4lRcgQNj6DSChyj5pyaYrIl0itmwvfm1CD0q4lHd5hC37
h510GmlnCbRASCf28hzt64uIWw1lgA+CaPUtNXfXHucCajXNjsfEF9EwqcDDSKPy
nnH3+Q98fGV5iuALSAQwnTEqB6QgYR3Syhymc0vQ3C/5k4SllcFlMUoDR35KpnYL
cWsp5H9LGlrsUZoJRpbj1ztOfPKFtI9OczGLomQ+K2Zou65birhBLl1ZOAyxhZZp
KdqbdqdSbEg8/bYQaV64YIt2PRFGhfdgCwNJlbsYyHxPCTMyLQCcmI2VFADUSJSJ
rZN7YwsVC77jd7aE/9ARCMKjL4K9cKGPIugVJ+uGZuVo0UOc5mq/ESKKmDYOZRru
IN09thQLMrMeee1EGRNSTp23kWWYtd9OpnCAxRWqXdWL9g3VditoM4acGRUPOw6j
wxQGJshM+IdU22kyr2Qo3gWpv+Rl3WyTlmajemD6iqOkcXoVoqQYsK5Ph98rKn33
Q0G5XQZ+FYln0CHMthr14jbemGxlrJqWay/HarkeO1tMK9vSHq8YXx3qEZix37al
psOI+uwo399D+XCMmSrXhjqImzdqiqa+m8YWVrSQ/3n6azaze8SogZW0DTt3L0SU
3TLqCPgCLnJO92D75h2/zJo7kd5X2fsQWbbW1CZ0xY+vXwYfCW2nLc1xZYI0YU/i
1ownGazKNRz7UOJCcimhLrvCEmBxEVAC1GmyBEK1IFDb/iUlUkgAjZwtjQ2mWZ2M
D9y+5BferZiVfJXdbyrwC8rIcI+gToI4UaK1UMW1uw4Z2AiDp5BiT3xt/uGIMaHF
M4aJg+posK/RGlZbbL0pFAZWciYb++pPXCqliW7N8/k4H345UnYViG4OcyVK5bVT
pNpL/LWNEtYC6XtSRBOF3Ka87Ye4vaCkISUhtWD6fF9hKmOCBAGwKP7uAEMi4nAL
t/nL9lFSJzoqgR7lJiBse3U6ynEqUMK9x1IgF8CNU6XLkCYVP9rRdE+YJ2TcUnCR
xtEko4I3O06jpziZLZlm01xNAk8aVwv3beyIgq+GH9fR9cjSuWKX4pvLMsJdbais
jg7Ns3bTM83MA6Ka5lOSMeSmCGmDXuC0hQdyathGpD+BwrfKg5iZn49/2xnkc6MP
tycj2i0IM/CkL/TrkRrvHHD+C++IPkSqo2+QEFylxPzL4XTLpmpBgN4MSwgol3He
MFqXNbSVGhlFDcihhEoF5T3PbO9Vqhl31gHiLIe1TCKAS8qAB6XD6rAvipic7euH
YFqNBa0pfuNcIB6LjQBxZuAyJB7ds0hNLj6ibkLStTPqdclToj+VpqQGjQ+GTaGs
5r5VQvE52k4njOGLuoHg2m1ZLk1mgH1k0zW32+aEhLo8TmjcmQXh6580EG9ObfyJ
D0fJ0MGGn33KhGA4qBC7kMJPzWL9aXDK0vRC+gpNsYMrPLUYIIeWZ/+2xISogC0Z
P5U6ToKu4OpF9ZdgTplXry+VSDu3nsoOZf6p027eRSxpZn0W+KXSvKmuMhvfxGdY
17iqWvHfn9L0J5dw4PK2EhDHozoEKBHF1jnL8NbU5DkE8kNYlJVTmWFmH2DtSm/R
QQtgZMOZPmrr+1ulrcD2jGHwoKJh0DaaaoxmV3XKtaDemg/9zxAsnozHCnntBO4N
SMAK9NEGfGuqgIBTbmW3/jL8REmgxnhK9ET2ZyaE4MdbHKXEktiAJBzH0F59aSIS
mBJLz/6LmiOrBpBZYl8gAjC2rvWIj0EYvwsFrcaSMSSWNCP43R+heRN0jbMcW9nh
IZB421X/qrKygQQmpBkrRlDmwxDX1mqq12NiQXOfylwHm7pdeO9AIPMD2CCKez7/
Y8LZSvukICvlxWCfuRSy7YNpgE1ZejTew+QaVrpcXJRCSOZRigZ3oPf15ijvHaD9
8zzVeSVX558oRKMAmqNIRPrwnJkmK8B6G0eJj1P06cGwKx3kH5MxGkBANdryyM3E
d2tqKfkvL2R1quesgHC/H4xpwc0MXnMuveprTNkYk6EC7Au3Vh9KpG7TJGIqL+Fv
beiIOjMdepqoleiOjmaVoALjBtC/mTiKTLjicecVxqjmId7OHgStTpJ+KXWSC2Cf
QbJOxOHqCZK6EXmVpdWBb3SL4wTUPLowIHYYCvynugE9i2IF1CjRp9rP4yCOcSUb
0dLNX2KjFitG3Jln1jl70y0+oiJwEj6iGqc08tGn0Y8DVBCp9Ty+Wb/SutA1bawR
nRAczYrzbXbDG/U/z4n2G+fb0+G+nJv1nCTnW0d0ZKUMT6d4H8NUPrppAUB9ONoo
L1A1sRwde3U2Zh2+mWHAz8qtbsEKUeQ/wvkR9QHYnTIlcIr9l7DCOeS5O7V9Sq3D
UQgQy0Lz6m4aS7sR/3dAT/t7rh//9TBvK6+F4vGhvTCGmEfYnpQJjxMXKCkvsbxe
shUXIfE+xQs25csB4XZ1Lj6k9f+1SyUYCwdhe0OHuwPXONf/aYkB1jl+exPt+9FP
R+f/GWtwIvNqc67KzOSZCexPgIOODetcG2UjugViAGsN2gv01T9tKz8O3OjTKau5
NZeh5q7ckH2FfTCBINdHC+F4zWpLrRIwxtPeM5JxUp5U1tnQjFX+zsW4kZr9yaxm
JYt+PGXJZDR90vLNwWZPfei6iGIMeO6x9XaqFIa94KQWTeQQO/OlZmBqNQk3PB0J
tEWpSBbZPHk5AiopdqkE1oGU75BfDom/ZGKSsW09enZJFW/DLkW0FP1OKEt3vOgJ
XePa03ndQ5BU05mnLYoudr0CXFtd3nGs7gfJjj4qQIrhX/a4Enso0epqFk684lk3
IEE9I0+ljL2Gifx5GLzXCGO0sWPpK6tSS2y6hgZXhqm+wtYJ+qDADZadhvmH6LUr
u093TJXysIyAa0JS1tTddo7r0tAufaUfucGrKISJ4UOxRbMaiaBxi2TvYet2JtUk
zDvGcsroYKmMcDkhOIe7YvS/57n3dj1J9oUv7cXIq2V7A5hzfzrCHXfYQRuFyjuM
A4tl/vdQYb0MdWL+YwIvr2HxW8hEU0gdu5o+LSU4elxcFlQLCOz7BtR7b1nGKdo7
sikZbw2KJM6eAsTinmhbr7zDitR3WJv3WOo0B2ahJSJNUCrWiUd3/cnxsZeP4E9z
qblN6TnpXJgxjZ64FLZ66leGadQvHENXB4wK6UUxyZfA5vzE8lvViyNW+wdZi+FG
R7zRyx+8zUynXwaNGesm8xPQ0GB1NKympqQOfrScNmDbsUUlZidkFjNjqQDWhu8q
5y0ByOQjoQrdegYFYb/SQpcvyJPwWMN3mIOGefZhp8aq7vknfpWYzRlw98tsk7Ou
RJLlV0Kg+26ofoH3ZbinrfCYU3SVbeuPklUVndAJ5H+nqwiQcPxllpy46is507Ft
jc2L87exxHLcjosIelbtwIR/wUTAqw0g64GvoAlNi6fEZTeUXhQ5VKdbLj1CWUdC
LwxZK44ikI/NDdeBO+7XtcrMzt1kP3ltPaD13lJEW3ohi2OGocG7tVEHiAIidKzK
Iu9Xiv5h369hGftJUa4ofuEoXUY/D4A6IWwq3JJ5G9qqNGbmkZsi3gaePXfjT+3X
rct7a1POl+2OaAoxhpF22tTzGuO8tyxYhczc+fq4Ifm8A/WgPOTe1epeDeF+kp5I
lVf/AOL0I8ibpQ+0kWkQt2+xjwsUKRonTo+cbthMBb3PfODNu0OwRQ8u19JZnnq/
rDocMbzCKYfMap6wO4aR0CiU3QrYZgiyng6aKEmhMasM6BHWU9SdWOCIM8RonEpk
W5zPEVbgDs82FnAEH29g3d0OwacD+80TJQOY3qGIQBFv/PgE6VZBdfOJ08wI6yD1
tVtYWzDOpr9arp7pPAOX9H4/pbSvl0J6GcCY7TSHBBBUz1aDUt0tLeXgkmJ4LWg2
OTFM5qt81D4eRW9hKD7g1rxDFrcU1m1fFlMVIfrSwpdRC4GtZFF++KKWWYrd6gVA
wy5uvTV8F5zsHSikLGcTU+hdHsIhkmwdpkgGxFpVQ15kp/HEDX38Q5sdLt3RNZJH
ksRQg/r0KIHMXnAwgSS6gry5auMrbIiD6U08KesZBqio0mijZ25/NtKr2x78g7Tn
t6FTcf/zYmUM3xOdKrqgn7Yj5VPJys/ARM56N9bH4A7WLpL9qbQbHp9RmWGqBGVe
kM9k1C7bOF86P5ReY5mWFUHD6DN6JNgpe6L140mp39bRxnS51B1U7VnFokgNEJkv
nkBNuze/eA6rPe2BvKI1MfDsvGEINnaWjoWodcbk5E3/s283S44O/2Y53YJzJgel
WKz9Xw1UvcCKroxvo1jYmW7m3dA4lpAHXITEQoIOrNsWV8oYG1ruI4D2GtSClFBx
43r0cfhwQh32mQWdltGv9Mxtw86a2j8hlRIT6toT/AtjgKsun4/7+ANSWs89mfTj
pbMsS4f859u9VNcD9iBdtdXNgEU8plBvuu6uE2nRm/5yF1per3B+6we5bQa461dj
0HOSUldhjILJwKokTbdokoff0Xt80Gfs7MKpJTjQK+tgkny2+O6NYprFmoraxci6
DXppICd54kXoLtw7u/UssLjKn9oWagMbUiITiO4AhLSGJdp+T1n8piWhuAiRmic2
irehF4hgTnreEVn9B1+pFOiLH10YsgmruCXnphIQvlN7WJ73jba/hj/bb6Mw83xS
dxPMLWxQdJyk32jr7EqwW0gnUPM3BWdT7bUiJ/rJCBj7yHK3KrKihrIrlsk0hwQN
U9UkqXKhLqtRFi2K61tCThuNOtltCLu7EkySDwjxlX454JYUFsHAciEU2KgSSfS7
euXDPwTtb9JOlaLwwnbTP3ztKooYfUHay9tgapeZz8lcqPB+fgQa9119WLGw5Pbk
c0aMBsPzaWf7U98AMxdWnZUOSzhu4G4SjfS3wr1xDhUFumL8WdF9R5kNoGLMa+uA
8CYggTnCdK3j65DRk2srmIudq/Qj6RXwwGv8Bh9XEC3W6NTXNWiLRoQjQSY7dKVr
wGu8tzI7JBC9JDWE1jKBVvUl46tkP2nuwiHi9jhTfH2FjxxTBS8irK+W+NycahS2
ej29hIri7lkSfZUUPMEKSUfTN8dZ0y9fjdPQzMSa/5h++ozLtVRjMWMcGtgF95g7
71GoMnbYxwHxyUgyI62dtJvYLWO5HsMaq6IT3I4XIXt05Dfr3BOg+HF39749oY5q
6VgT/NuM9Vqnu0L1kn6gn+oHSQPkeNbL2AZet+ZBf+p4WR9g0fehUNR1XZkTrpQf
l8wQgrX+GA8bYLFzqt0Y4DvTo6lVgqeLym7cEVFla51SxwbQGoviry/cGhBP121O
OCRMiBcHXA093bXo1dcWGPHDth3sZnE0dMCsOYNCB8hdSNKt7MYAiME3aJVrzlri
iUOtgFIO5NzLxHJvlqCrfgYzMraFvnzljj4yCmf2ORhMKJBG/UbcSGYikWYAZxYq
8PzduYTSFfT7wCNEUE1hT8qTcs1YQGgmTikkReV3M4C/6z4MYQviIFfuzjR9UcGY
RXUsDCXuVqk03asKBJhmac52fjWGaPZvC/VY5ut1DiS8ZckzMCARR9WgqZ5OeE7D
DaPUwa45864xwcI30NoJ2Zic/b1zuG0iGU/p6CXqr1IQjLt2/Gw6JSoNGXc6WloB
XTMg2uB7uE5JY7UV/0ED6Yeut5qNIS16zHxyCRIcylSEE+oAFcqKJvS/14axbnDU
oKoBv9KefVerbwdW/8TW/rE/SnYa7KJLhE97YoQkUmFI82nNLRp9iZSEQUJ5w3rI
VoavY0GRnx7O9ctgUi107rKVWnmfUsSrRj1llfn53Av9U87sfFh6jwqWwgxLyRcO
j2Phq6wDOfYO7UCnkICSU35sROzLUxTtUQa4p14/cC9ct4hHhnONoxLOkCFjWOPB
/drIhT+xCAH3EBJWfH00LayiaQfce1otpJP/1Klfq96t209fDZNg0uV+d6Z/+KN1
5FS4EB3kiqWHoxsVtc+ld1TzRSamlLAD0p7u0u2sV6ZtlrEwlBsNcp3DdQ9Ge4Rs
Z2diSt9Hpbbe4mb2BrI95I1Xjov5Rj4oKU69+IrbHEjZzaE8ALLGwG78AZACBA5A
zQP0ED/vukboXG5SdY0+ecr50l2tmpe4Xed301/gr3tumapvMubs2wgcPEbeEl0U
pY5g4X9nJVVlP0Plxlq1896jTElX/e4fqzzSdkN0EUCksW5F6KiluRgKGxXMqh07
94EUWhlrTgUXtgnWJHo+HRHtC7Z4fsUgCSmlGygwQWuMwnwWwbfmDDTaCD1ypf0G
YBSWEWc87FbukwJE2hlhixyvVTLTCgffk1UF/KPPnaZsHcoqGy1p/qzHr26BhRtj
QdqkNWVCeN3vYqmtOaH25Dl//f2vsBJzWZa5lBIZ1K2gf9S3xeM0a17W0OfsX7LI
vHigcEKYAbl5w6BrJ7liLsQlut+Sossbm5q+zZTdo+5I1nJXqk3ZYftihPj1Yeea
O9ZjuetfUe6k0AhsNR1FGrneUPVNB9Ygk9GnuE8p9f2B08lgBILnnJ+jnIHIx+w/
hrJ/qNI3eiXHN9YTw1flMlfTVnOR4q7eGsl2n1WOkT3s0P70uKwHqmNryXmtBWCv
nmLPreFxojEbLLsJUs/o50XuBYXGA7z3f0cghVpiIoHlgBO1IYIhQiTD8hUGBfGS
Sgx8c85NKu3cveVbTtHTnPm4ac3UfJtSBGEHJ2mKzkyMKFItvRs3GLkQzmHpIiRD
ENlz7kVs3MKGrjuc/wVxyCcDpS5y8nG4NWGd394s9AU0vq7JYwtMOfZO+HT98xPy
SxA0ecAWSG6S1yDg/a2x+FrGBCaRR6oFnb5P027Uf1Y+14IexQbuRjrOfWMFU9Xg
k4vnLwnGVDx5U4Cc8KUOk76WYZV55ycDyQj9HhesUitEUN+0lp62Ua06YFih7SIe
8hcXZKN4W8PnD2Qur/eP6z2zsGB/L08bRpGaekR4lOpISZiq/3eU5Y1t3UGCqPm9
0U2OfolIe6bTmqbKI2PnpP6swfwvlv8zaZ5n5AZSRxxtosPbAeG7iD9kgJ1zvPgw
hc+8VKIsfhDerUPwdLRhy2xtmcRwkW5E8KN+W5dcXBj8Koiw5aIV8otV8NBjvH/6
WmapWeCvTcM6EUZMosiyZDNdMY2ayQoM1dCKaDY34Wl4bU+l2btXAMwhRwCqpHnV
7OYXduAkKDMVw6Y3LJIpyRmOKHRlgGswAsh8N+BLNxUfhFNM4p3xXfQigLEyQh4y
Y4ovOuIJ4awAe2ZySQrSGYx3BUcWyxeagPyBFG+1kxiIV+8LaZ98QgCHBKOIJaeJ
ud8vSo1ayBT2omreBURTDiJnamVM+BEZzWr0iRZA79TsvglOQbdMhOjn95ZZe+u7
TjK5GXkgB1YZsjcNglrimrLo0gt9wPZGmiLMmp/u2MnEzjq1TDCHj/5eEB1/yI5l
AAKJ1FfAxJg+ig5nO/JRKVFvfv7GE59QKFzeLbW4pzHSoEQOcQaFmJDejFBqHuUm
trhrJW8YHSLHwuz1KAe9yXTh3zl3yYEmMK0JKC8kdWYm4PrbUaMji2ptZU6US6K6
KjnOgRSGc5+bfxHpEERmA2/kKe0okW7kZwT/kIjjxWPR6X/mNyeN8j5DPsOhB67E
zigyM4l4EgBTj4LQUvikz3fY9epOZvgxomC++fzKtyB2EusnKbXUN2FflHr56JDi
3KG3pEJYIb7sxWa3dlyprBwQRdPZeGevBMws4Q5z9oIysENweM3CS2lEByvGKBvA
Kgkq1Qloy+I6bdJo4VcwOOmlJZl3qYtLH+/9h5rOAlGMP527QaXjD5EjtcGJCYHo
VVuPr2GZBv8slwOD6FNlS8NSKKP/vmkYN7VPZtUK2ZG+0o6oOKINQWksS9buquGX
YTFxLZ1/qqAYTBW1kBgQbR4NqPOPJ3lDSXRs6N06YtnY61ETOhxMlADlIwKcp3kZ
47+n0Q+cqWekYmekwWjkVtyv5yRADIWxIcnhn7Miu9IpgwqNyEpxhoChzImsWU1S
RBhHEN+tROqPlHQZF1JepeHfOjB+9bDasgG4f0/TgRsJpr2WrYZkZHtJTst9BJJP
Ucn/XewHac8I3lduaydstM5Qh0eMiQ9Ewe2qICp6CviU+P4gj/SLlsa8Xbzl7Zkc
aRsWr8rT+vgH/1CIJuqhqJrx8vQDQa7Pzr52p8hxsK/RzAI7NTXbyhUC/8wjtnP4
RqBo9ODAtvD7Ew60ClsxeTafPDWrVSe5iqGzS5yREZaKu36/ncwmIIw31LFALkWk
2rndHWqaxfsXKae2LpA0CrVZiK7tTsaBihT+13B73T+3WUtkulzrqXSxMW3pM1oc
XBU+G3tAz4VWDf8VWxG3lzncnaJjk6QfewTnqHSaLHWqL462/I86pL1IYRZb8ZfF
7pBjnGo7D5zbgf9HTgPg1GWgKkiNQ27/eAaiG57lybxFOj+kY84kByzwQz8/QZxF
U4gc2REHzbV0lHU6Y5m0LfSXexZiN0faCe4ydoZ6EwJm/cn/Qt0l9wsYgl6PL7yi
OHP1Unf8hR6mVCVpPquxP+6oLcncKF2u2ouedzmGam5qknvvtbcxJjC6Y6RlVHUo
Zj9gGo2SQCE72TlLX9eTPw3E19SUjUr90SQo4UUHgBdo6yN15yPgJuHKiXvQD0up
sdsOkzmMjPvZ8N9yHk/54KPvr46zAeMEk8XdI/8eg75wn8CE8wcjotCjLIsCvL80
+IC/HGSCMEj0aoC5zGTON62foDBB5ZTyM96/73LhrR4Ug3suqGsV/T9ARSGpgIlI
BTO3oxABJmClSWtRNaZX6Doa/tPQ1pQJniVMQ7jcV7veLa0LfWz1KVaMRMMlwwPN
172PKXdqoHyI9pnK1CbN1KKId4H6qdjpaHKqWB9jdgzwa3gQmMBhmTD+6fHCC9lK
EJYlvzf4DdkJVVjZXV4v35VwH/NUpqG0ntGlFS7OBTNSt9+CrhJrrlRYZrFg+PcH
7SobuM1DaXLxC9+OW/IHNKFkZffi7SLymerqQapf+h+P0Qb0ffHGVkX92D11ZZqC
mnvuX1MCHov1flkEELsZcaX/iA76ALs5/GKa6mTijSuqgOxqyfo4pK0iciJOYh+b
M1prp5I6hc4NKWRdQB8jPRIEDkaViSSHTuvyYy1c65O0UZNl8xnQi24on7Jwucwk
up5DnNZNzEYi9FsSN7/jLR7gojmNiOyb+FQhL4d7mhKlabqIl3ZNCjvmIEe5x+Nx
qumubibs1WN4MjS4TLKVEj10jyd7uSCKFW7axrayWGgjHi4J3GyMBDTYDAb1+yrf
K9gLS+wp+G8hFJ7Ctnt7eHxKRec06k1K8dHMqm9jetsMzvndi0REEEmQsC4tmpbu
hXmyjW52qACgUM/fqHOkhqbbH6D2OouovwjRvjTOutg4CQ7Qcad1mVkF1VDa2C1S
0SrIqsRJst2Gr35fGQJTP2j1Ldla+EcK/J2mN3pCR3ja33aq9IUMb9sd0S0vTO4v
K+kVWW+bGcBmuYJcKTrt/0nA6KxMUpNVAeGMFf3GglePWm+CvvRjqoZr+Kfvr5r7
mvOXieijLW9ryT54iurWyF4psc42TjSxxg0v7Ihpy+Jcu1rtaeL9XOS7WakVMHCf
EykSP37fSGsZQhE8QwHofWSDd/GC7fFzeZMEIu92Ozw9URuCwRg2rBAsMD2nh1KU
Nu62tnxtb5mP9MBmsJfoQ5lEUlZF+Tn6EQvlq1gNOfgZmn3e0SqndFW73SO7TcDh
X9Jdw8BxxnlTeW9RuYLVUVy5GoFzw9Hg410QeYcbDhRmZ7qAbpDpA/obFSDFsYYM
aGSJtJftc+GwjmYJX+ziGc3IlAsrOcX3fwc7nvACnk9TQfX7LzH2G9JjVWVecDMZ
DBMYyBhuNM9QA9bvOin9d7tl1LvmeKFMKjAyfYdoiypV+0SPpDtH1ox2fF93LcAt
UBkVQ6MoCPw09xu5U+O8khm90j0uS7H79pM0ITqm+nvOIQR0AvSr1zSRJ3Ags84p
2g3JRfjyXz7R0QqmWVEUSb/VU8iugbDfpM9a4uwoBwOWB/pUp3pydmeTzya1mPVU
wpkNWrScdR4KBw4Up5t323vmpTxP4oiFSak9C86uB/TYuzPaeFh1lhK1+W2zjSui
hHqDAENEypmh7u87VwC+lCaG++OcknVPSoOm6oCp0RnHvaX8IxXpvXiKNAj8ovxV
ZMQq1W98ihXcuw+HU5MhkuencoT7ToZiz8NGf7GMtUa1l+7ijLymeY1AjIBqGI7p
eC0TNA19dGjOqXeAi6KK40H4qeAY/ySOwEQQNDe5Yhwd9MnzFCC27aSzoBzqya3C
3DhqY7LdSe1jNrYJg1IdzDVLUi44vodtVZpld3P7fyFIGlVnuWCQCG7/QlbsuTeI
fWumh3itldC7F3hvMBhCa67Z/S+qEZHukBfOVqvADgUU+NKY3PBNT++482aUXE1y
1ffKwn2+Zb8UappQ67bUzWUo8egwkFK7FhFmbratJ9WA9jVM4FwV5Mxzoazxw2vX
e4aexMgIiG69kpGMkGme8ujA2Acfrdla5AujD5jPuI34cgKr3pD9pIIUmrOJwcb6
r5jVpRkiEGE6mp6wisms/J0/2nxdLVUejCkC7XK2gp/1HXgaY2HEI2zdAmPlQIxt
aV3f3WUeoTsVBkZKYfV6WIL1rmkG42bOk4+bS8W6jDQruBZp6S3hkJxz01WZFjRk
RbKcGQhZkhVljMXaA4FJop5Prdp3TDiHk9YXchUQyKtb6tpzjAP0GFcgfqDlC6a4
ykiTdnEb3Iush96PeNqSdpBt19TCAT9nFtA+h5q3l5xVNwDd+tiMHRnkK9Jowhhu
HbIqpj7/PP47EPKXEEpx7F1gVEU5oUc62ks4TRv5bm3ndytcj7FEZj/am5/btPCS
epOk+T9TmWRZxmLpC8bWzuHE2u4piQk5vPF1oQKadQAZl0xqFbWvGCeD428hLPHR
m3igvpSBbRBbkEJ8bLGlG2n2M6XZzvVf0yCzud9TlxcyUA61+30U9t/g9D2FMcZ+
5TFcLxEb/sax8AGoCbK3nBC8w98TTZ4WJLOoi+MMviKOeXFJlEgEh99zntUVv+Mb
MnsVjaFmg9Y+OGgm6TSx5KeFRfbjR0xGtXvZJUDyss86i9rGk/WfmzmjVqB0guOo
IeBFPC6I2RvNii1iidXO3lmDW3zhlLEK6PFbkkIuAAHrJag67bacTWRrjKTyaGsl
Zufsanygv2YMDXsOkCDCfBeupZI4wJjLCjiih3liNB5oIrALfsg+4S3UvtH1OI+n
voDLWJx1JzQXJL4Vj2pjrSI1YxCT58VyHxTKf+jRK1H5EoPXlQD+hZkqCuYNwOPR
afXqVUQkemkaFUWSaubZqJ60VgpVxIJ9NbGN6rFmN5aJaZzMNF7Rpev80Hi7wGdc
8CIKr7TKelhtc1CHaj/0GOkaANMQsslP5pJwWxGJF0+xl098xsv0Qgn5FemoUCdv
HSDFLgP1fO8don4G2gpY5N1MDzbXlDdDlf804KYkir4=
`protect end_protected