<<<<<<< HEAD:flexrio_deps/PkgXReg.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
j8CKRAvULn7NFOL9h8Ek2jHLzoCpEgRSwRgxdOGQjWNkKl8Sj3Om4QOMwRjgOH7t
91sEuzZsuTb5kS3wajX0TVIHmakZ3lYqCRRAQXjKR2j9Yr548nbLu+ZGFvy0jBEa
op64wIb5lvjX1rxDr8knEyjkN6h9Wou8thApRbB4To8IqMvqCNaZGTKaz+jagwYd
Oak+ojn7doHqQ4gVuatHNjbAVmI3Bo6/05J+fIzi5EvN/fZyi/BVPQ+0Lyj3weKa
j2Xhy+qjQ0uOOC2EypM0Bo5sk6m06pYVN992q98YAZ2sdNaqbXAQMTaQETpppTYJ
wGW8a+W4mFa6a4az9Iy0U9ycQW3xHe3rzuSg+ooTyS/VGXJ5/TlR+P5ad88+wBzN
+AsFYWt/nxyBSXbzMvvJrPew6u6WwUtKM4myBqcWbtlVLtV0nGteoNqUE6Bu367/
QHQ6T0esCTKgBOyrzxtkOad2kfRS+MTJzRSRTT0hPT5oy2NbLpe87B4gup2gebJZ
qK5ICEcm07KZxq2NNqhtN0GDrFYr0a57q5idclkCw45zF4RpMkrpYi3+UOF3M6G2
90U/044O+U5SRUZAOhg+d5V3eVhPDsNSMnfFXqoI9SNd3WG0qUGw8KKNlWewqKXS
C7XM5A2PkJK1ryqYKssa+JYcD6Q6v1CFH6J55baQR0d9W3LBHd0pnvbwW1yhhhyL
AQt1eMPIMneym2ZyQ2GHeVN/XM7KvBUiETSFBTzmRstF4JVxqsPMqY4CoidsUVVE
YfAU1RXabeyb+N0qro95wIyYAWFjYX4luAFbYH68PWzy6Gi+ERRc3/eQXFi25TH0
BrCNbDWr+mjufDllJkYbK8W8ORnYkzI0UzZP332kh8zKiygu7cqQ0Gu2YCccFBzQ
QTF8rBdZBZgRDfOydrRYdq40aMB2MZzpu9XsgyL3QNDo67gDp74/GQvzCJUutVvz
xjQ2gszlgDur8csoDYvlZAW5poWccfEMTW0fMFvzS4louxtq94NJsQM4ALtOWota
Dv7FdI2x5aUxUK0jb4rz9QyOSDTqrmK4CaUyBWcCPMIsOWcjQlJlVpnIimqNE1DF
ugGjicAVIL1Wzo6fI4sj+ALqm/GFdqfxxRl6HCU/rbyYFeeH910fXE1sloLu3kaO
Y1TUkG4urORX+4Ypg8mj4gnG0Kn9gnNXGX+XFqamCzLxtf8neVvPaJN/aIcNmHaB
ZDQCwXGk7heKNVRueN0dyjaVgXcGvsAXKOxLifbcQBW8sYz5MWD1zvf3Jonu9D4U
pD/BZSG9lCQn2K9OSBWWHToYx54RB1urErIFFYr3ceHpv3lRnoJLtUJvTSqUJe5C
PC7AH8ZKJlvDw6lxX0jlaJ+/wdQNw/wIYaiUZ334fT2Y0RpgaM3YkIdAKEtJVpIs
VPI1LJ1BBtueRG6idQTRr70CyuxWiik+6y8mAsCv1aV9Vi/1wJ45GSlv9E/S3j66
SLsqmYdhUCWoghmyrJVp4zZfoZDHSw2crw+4HqlqMxUquMRj591GdUCjk+HTFLBQ
krDPlLdk9ozXRQs/7e5JxufDgBJnHeeM45J8VTyy0JUef0TQyVrG2YRC6MxFlHqd
jI86qUdQEvAxmLYs6bOyYhQU5qVbHjnx7H0co5i8rTqDKWJoOR6Xu6zxJxcSaEMK
oI2etotkz/wRKsjzAGaV50DPoKfb4jG6/nhYbTdHdPKiRrrcVD1yhZWYba3e3weh
CZXDRAhlztFxu6TUejs8uJKGFxiYs+9Nkns4vmhQ08KquNEGKg867x7qhDMopovX
BvxxH10YqEItWBLzp9Yaii60bEfOvqHLY5WHx7aNf0DQig3qUVkWkBuzUKSSHowt
vLalRnmvm3yEkS6e2XskwmDCFoC8yjND8/tqhnNQu7DgdDoU+92jwGSjH1tf3wyX
xGHvqy4448GYJ8nSzWBCh0hBQ0tCm1oY5Di4JiJTlX20YxLbJYNw7+SczkrR6eby
cIzTl2AilVcUsGTpkbWIpM4HdZM7UC0TBiEt4vtYcNPGls1KnE4rSloDKPmE49Nx
adwDdJdQ/n3s4rQhMcDYFH30DZYN2DdbLW3+aWuf6XWCqTwLtez9ykJGMWzOfwZA
7oee/40MR6kFc+T0/EZpnhq6LhVLe1bJYbvKNsf0RO128ZgIwbS9pPuvxic6lm9H
pcDi18kyHZBpY0iczLcMEVcQ7hDvRSQq9uMd9/bkCTZ4jszD3E+yUKvY8CeExVGM
HoMSZ9/p0BRSKSQPuTH1xrYTeRMOZX8oa8mEwAtJ9FcwFazM98EgGyhJkjqt+XIb
KiYsAbK2xxGYSmc1mBYoPvq+mq3NKR+hwQO8HgZK6BkLuHJXNYWlWFK0kF3P6nqj
bXN0eokfLoWlhxgcKzhh37LFOjv8k6oHFsPzcgrvUIa1/pJhfF44veRdI5C3k+Rw
nMi4QjcIiot/IyDqb+Leyxv0TGKgIfyVm9sXKYnzgfXoWmuADW4y005a9JzVkRo3
jD0NcF680PJ0+5H4c+SpNqMZ4IKA8yHPhlzyYlzrxY+WZwjF4DjrTW0YPk6sypQy
qpUXMe+k4qQf4Y/e35eW+7o5Ssw1DFzSIsj4Cl0f6TE+L1Fgnh2bD1D1O5nc/ALr
p0Z7tkD37ecHpD/hB3xw2M2v3mAJeQ+u2vi28FboQe4sBEcKWVDxDJh7KjpOaezI
cz3sU6ox6s5XlhvupnH+0uO059DXqN7lr+R+kY7yTHZyEojUIMXYSnVdb9driGHc
PonxFT3Lel5jV8/yFZLiPB5rCL5ic1Gc1okynW9HrlH9gJDkuRSzm+sDulqLpzrl
5JiQB+QU69IuFfasN8KNCzEazggY4b4DisghL4AUzYJKeMhy4YKYhnAWsvvIayD1
6kGtfr6Mlshg9/UkYfHEZZnFuTp8umKJnKgqIkGh2Ju13eUmm3wCT59ydAjfjBQH
dLzJd6NPCU58Joy3fOK+e0S2QjTMWE8SHOqaH1yU97fQaqHHjgMEKraInXocd7d3
RzgOHaF2PukMQsYofibSQlWyhK6xmJGHYNMFp92ku4zkUIXLyqwTNS2SD2+j0vJY
ZX/q1zaAVBqhWnXLV1fZ0zjIglmAVT22SybH0Idxocaztd3CAny9FKxZZESE0dK9
4FquYNz+2j/PjZ2f02Hs4jhxD1lcGDplENPNwTNGAXNhTUbzb473/SaGuUlM4SKg
zCGOT7VKpP07tAt0peWoT/XZlomgrpniHga8lwMcJ/i30yRjve0nxXwgqFGYNgNC
AiTFS0YAEFPSSSA9MXk6nl8V+hMiQ79Zm4IJeq+CZzrHqI3DJI8HHar8Lt02LkRk
x+I8yBX78cZK8bRM0qAPrsJhHkR/kdC39hxNssGYDrrPhKkyYM7WKeEp3Ar6p7Gi
BRk6C2asW3DAfIEs4uAfoc7HFApOs2VPiLO4GtwxXNERo+wzPKzZBjbRzHl86rXz
eaen7sec0uNpLpVla2ozm6Pp+L7CkCgjGQ6jytwcjt2o/8lFXYyG6leJw/52+p93
EIGWlg8JBNIGBdtsWQ66awPVtRD9lm1USDKe1ddg0Cn0WTTGkDk2ZepSZIMDrYc4
pIlCTWerDKiwLnuMcV3qTsReAAYHupaomgZa0celbPGULRtgRCk9zjhLC+oFXOsB
v3CgT/AuQoZOvJRhfQtw+9BKoGgeflt0DIhVuGpd8tD04S7P9f5uMmhR+2cOsVg+
3VJs4iWmyCqHzLy/U6DM7e3CMTOCegdM7N9xgagyfpe6kYSJZ3CX7Z2RAuYjp8gj
lI9EhMSDePKXwQS4jMOij28HbE1YnhaqkrcQv/qnC1YaYIJMp+Gi5/RKMT+g4fDa
ymusE+ZnMw28WwqkR+pJ8CVtj0RtET5xsxNvdLhi64o3IMnrZsRuJ0EVN9RGur4X
gpKLo8JhevHdbiunQ0XfBj6lT3g1Mm9GoPY2DCCNf3ASHweeSQRs582n2PEJoHUn
JOtBAn6hiytlUb2GKJ/YbqO9r5IJlYFZwAU0DR/1b7nHF+pTdzbCntCWE35jPt+o
CET9Ag6O+w9nGtb2kv959FcANfazWSsQvEkxpwKMcQyykjGf50DMNH1kiXuT01hU
AVl7NOTKrZQzZG0+z/uCNNIqGiG0vYeqI4YwdfwQGFjZUFnytUft7ilKmVNKaIVa
k7i8w3s0D38hevVqL4PE+Q03f1r7ii5gJXJGUY+oTMYuZ7+ZD5hs9aV5VYEPYinp
H9sVcarghkO/slPfQW697IgHbzC0lxKB6Xc3WUZw6voemQy/Dlpcil+X5QozZOMg
sZH2N591xKQCF6S/p8aLFrCBYdBpDvQ0Re0Sho57mqB75BoKW8ctbHniR0H1F0Z9
XNoxqpH1xD8g9tLCgWumt+LLz+Xqb7vXvdw5MnKSdtJl3H23NrwRA7GWLTCknhDd
yb+SeLdk8KJXenlX6n8otNGKJD7hu6m180dAgakZg8k0smxiLC52FwortY/fWUV7
o3arGcYuvTJ4UlPRLXT8xPhi/mvXx4HqdTYxvGyQf2Xudpt4PRLmMN+gnMqavsVR
15DwJINVSFjXqi1hNn0UiNTRudpZqxM+wqQeKTjU8X2tsU6h03QQLIHON+Yfz/lK
bD1f5F5j7UmborypgIVbM71sccI9d7L+Rb1oh1AQXq26QJchyln8RSuXuunHDd2W
Qu0V+1LczUYX+Y3jjiLI9t+aBkB7yBHPXxc0Cg20+LeLLsif0S7CkFkWoZ++0j/Q
32xlJ64twDqFGcm1TNX9emq6KiY1uK9OfXCEOOaTsyIgmk6FFAhoRjvJyTCTy8mE
r6C5Axb4ipq6nHHboCnkIcVm6IxG8ZWg6WFfEzD2rlY5DNj1LSagsupqThGLPM6z
KVzxLxYoBg5O0z+tif08UPj1U6T3HJqsoXax0eR1XkXXEJO85GjYkjLISEmN06cu
EGR584GiVfvk+3OF5Y2H51CN5RhMzeuUnh0IHkBlXkxCgKW7K87+yYYdVWCFUJim
y0EfjLVdPZ5+kIMgND+SKe9462tmDQbK5CXLta5Q3gzZWTocrZG6kodnPmeSr+nE
mUA+WrCmBvyb5laMKSnmVuRFU0trWaT7eUUGHsPcLC/ynRn3tGE+VcXpFtIbsnGs
YVxByGEyOY3qnuYMUNCQ1sPXOEO3OoUfFdEGPGZacWwbrjNCCCytKrxHhiAKHO5z
34JfxGmoDdja3R429H6Th35494V6Iio/bB3nqdmtIEkVSM9Ib9pr95eoJlD1i2AX
infhq9nPeAfWMQnTrfdvjVyXF7VwkIOsN+JwhDIcyDuuC3qXQ0b+Q3s8J90UZZEL
WUQ52FGZ5t4wYanIK5D9UgvZQVLq+Nu2ZpnvUhioJFGYVfZphAH7NA6fr1sAzZdp
8PJ2ywLNpXF1eejQg6tkBi3iAs1eJnbl/pEXEhQTQI5esh0oleLet9VVY56gIrlk
JNF1r3helEb49L8oGqCOHVnYNqUZrtXzVvlVFDEo1uQDrbDrLqetQ2dyNfC/FKHx
vuVXu7FwfJBzkO1eWXugxHxsMnH7l5Mbo392NPAhchKoi8UBr+JcAJlVaJLaPpgn
a/Ap1pUrfMRNArP+aPPIDO5Rxr/7Onw0Gkld9OQTHAkSNm5Lu8Y1SrOCPZl5PUTk
Tul0NT41zr3CuvCWpyto4xnV67+mg3PhhNUMuz34HI4t20t1/bdrXs5Z8G7U2IKu
xBemcUvmACFfuGBQl+v+gd7xwzjHvs7TtAF8TwqvGisuDDwJ8FRS6CiHa+QoFdW4
Yb+wKlktd4KpXXZOFcXRgiqLQt2L10wiGH+Uc0G7pSGOUWCbodS3bmZSvGnSizDv
afGF6BxV7x6zmc3WXWcTxxiiQw4sESlYJBhFHS5yzO0I3xi9afHi/FD2NF7VowC4
9TRWJocfJ06s98h1FJXz2HBr+DWXXeZyc310r9Wxmvo/i9T2kJBMG2wF3otPngHQ
IlTdpKzZi63lZzgl7oG6JUjj5TVwqlttiJOUGkmnq8OBZ761EBy7ZzB2HCmOvyfN
esPLgQbgtAevWrlT8iN0LPyJHonz6qpVDvHHdNSVIiA3dV8bu0ez6CvlBy2T9/SA
Ze/y+ECviLEBv1O/j4Lzid9ekpZduQo6VqjLFi4SOTXmKCtouqAGlD4000fMTBE6
YD2dvYR8CE00L/Ef/QJMcE61W2i9s1B1dpAsbS4q/GGmO9lyvg0xJPPR1ExYCaXi
lFW+56UIMzOu/cn8hec/q6nHxfC8BmOXkshUFxObkZxjktV7EeHCKA95DuRwB0t9
nlLnauSv/UdX9GU1GaZoAh0q/akWNd/pxlmqMceAD1H2AmAxtQxm1i+foaDn88hN
HeRMl5XleRZxRHMoiFNs2VmUSNLmcdaBeKxga3X5VnlwJUgACMzKE5WV5+FZaH7A
Ucm56YVYQIN+oSw6VhdNtvcD1haJaMW6ilUz7XZIg+/EzKzGYxxi/MugnGwGCNCv
1nDIFsxb9hmy7r5CQPDWLeZ8YBchjAmpLeoKADUMCIYWrErQ7E1Wc1ZniTyN6JGp
UVVoCUa0RZHpYSk1+2P/D7Ns0ptGLsz0Anqn9s85F4a7ueHeyL0jvTa/IdL/2Kbo
8lDhvi6exXzinuBN6FsSaHDWHp+VYguTpl8Ier3rguuZ72Cktage39bS08L+6H0E
HAUSU7So0QEOTb/bX7XmlKh1BUz20+KUpIu9m6kKEU/QGrN0w08RPpdEL9w2RfM9
6xs0nIxzkmNEYf4GBRFADeoqYsYzaacz6nkZcqZNoDHnS8ijoLuHRRwFkJ7gdqTw
RVkA/RAA2dxvO6E89u4GvutwdA6hmQPUFaTn3sWrqePGBxTbAN7HFZTPFKijXOcB
dwEF+DFSZ0DsaXiR1mmLoeL2Jr5UwDAsnD4KviNJbiHu6uKOYSe13Z89A1tauPGf
oXV29j4ISY/yrcyQ8/3VcLk87GxJQYJzmLY5bBXAUe9AlNMUT4WlgwvWnbjhENtd
Aonlkh5m5EuOoHHvuZfqjy3KZ3P2YbGaXhG0DM20s5DsGkhu5uvvxml3y/7LsTVw
t3DDRyz0tVOaCvfa/z0vBsWhTlDdXpWOGFLRJOUy0ov59+i24PU7zL/GOArJmUD/
wIHgucNd3wHvyOjAVlV/tiWfNKU4nEbivskqYBgHNzo4sDuwLmb5a4dbF7j92VSD
GHJZfNucNnfXucWKbuCclN4fpT7XcFGBnQjWVFKo6lc+EDYAznGwzvxXNqIHarw1
6zo9lQPg7gJe5tX9GJhVqQJnlQjL8vpkGA6jqZgP3ggDXs343gyNLaImkoXW1a04
cjR8L8aRYIw7UTqcBWtfkecFpkMhoBB7caW5krsBwHxFONQ4vD93fK8uOKJRRrBp
MZ8eDPcfis8sUq9rP20EqpnEKf8GmusV8wJOCIODMlKM8cKfhDZaXm3FdQmNfGDo
+5XORgr9yhxOaj+zTD0q/axBdQxm0xyFTKWVDaRUrjrwx2DvD1d3iSpnK5+3xZGA
JGsNbO/LrDcNfuxGGlS31xQevzCuk61bV4V2taGtIvApj3oZ8iC+fXPU07/0w6nM
XUU74gNQ/B1FfQAODkSD6DmBMmIt1QhAP2//Iu1zB3XC5AWdcIi4GDmHtoNa4uyB
ZNgefm3qg7o7CDx9UYhAlsmBcmx2QSY19kVkmky4dAkwGB26G2dbvBaPMPdvdJB7
U/Wq/8IY3EtB7OS2QVahs6me9HSRGxYTxF8JqG73SeNknNVE0bMxbw88w4/QjjGa
8QaRg8MdengJAtAOcdUDeCwi2EcQHStkK/VjRomYrydmvJ4YWJBSrBlIbNTP4e13
DoPn8tBcRXjtApWWA6WGQODxBKEodWVbikSAUIoOk+RlegaKZxcvm1RtHRqpqntG
vRKXJO8XNEa+verYisow1XjmB5KhxbQZ0NrIHn50oqA7wVk2oswbVH04bBYMSFQ7
Qi4hiVWDNoTV6OH2hki/yN8uTSyG7Y2pEQJgskpBBKpjCAB9ZGw3hCcedV0cnBsO
Or8hZDR53PMSk8ZUP3GDKC2Ld31fiwlJokDUCmGIJq9IqeP3Yeitrru4at3WO/wa
A+rcIZlbRbV9eCrNTQVzAeke/urbzriiiPAyg2RjhWDPiBnIiti8Ai6WFByg02vR
VGLogNDIt7HDedLnxXzMzwTQ8zW7mZ9HSwZHlwHbuu42ixnraAPxVVovCyLXrvXq
Lhfmg3+9q38SGU4KTgNL+jx+RjSDmRgXpd9DJj9D2/2pvmFD9CN3jmE6zC+s+4wf
E4ZjyUX5nLYcY9xJtCqnqvXxP7Z+vp7gUY/pttxxHqHDGebD+BJPV2gzkkMs48fy
BPFvCw6/xKq2jvWnBiFpxGzgAcOYNkmQrBaQkoY3siRPeBZW5bpof0PcKd9f5ObU
Lf6yYscEDysZ36270/E2ZYw9WuSf3djTNKC9s9NUhI+QWgGLopibZl2aRLvy2fWV
G8BBqrVLIFnqhZrYl5p1zO/mKXbXNceMXeFj/CyMJQUkorC8W0UWvrGstV8m3PYp
WY7ijTvQJd1L0WwtACWfk3w8gJa0XGRgLWwCzN158uXX0RUIGlDYY6ZGwtSKdFOG
k8Gdqsfd3rloMX+AhibrDErn/vFtPH0DRsCz9XSmoql5ee8q3mRTcxAI0BCjgN4e
ZeQPGB1qWFU7QWrZPT9luXiPpUmNMWCLnV2rcbxgjaDXMVYY7KB7OYMVXBuo7Q9i
kljnzUpDH15DEOWU6i3TMWAoRvEFD7KwS7JoIHuENxCBEEHq/gzifqkhjDbe+Skt
cq8/SOIrHCLifo8NnGdWNF+JbO/d0QOkc5W+UyDIDCqUs/l859B3cBPdXsE/TuXH
g/sZtUJl+kJmoGyIkiU8YZIPJMviTy4/Y9XEmS2A1GUGXBUbltUW0IDLPZFdnHlA
by/GbQUpjsZeVJhwH/JzogvvQfhxmxpv11sIB+rQ+Bsla8wbdX8PsXH9M7png4d6
h9Tg62zm93/kEwbT8imVwgSxbJnC3Aa4qAUYOGQbPp0YcKAUBPYJ6hTvevn4I1dt
qMoRrb01GW8Qy3OfSd/Hizs9xmFHzgvPZy2DZw07UD7RQpZ8xAlOBUXeB6b1AI/F
o6SkRiUkQ8LPqX/mwFDQH1/8QVy98lBujx2/VVNF/2W+oDIj3NaBqTVOFfNb0HAE
t7TH5slNR+RTWBxAtiQYkP2uKVTny+wfpyLDSePmQimrxzy31Dv0BTl8HaYIf4gD
T82vc3/hcV5gvLtzCI4jd2ITcvQaVkfYAsQiN3I20Sfcma0rqywWXnOv9MDAugps
7Ct9GSwjoxhkldq7CGbyYTwTSTqZ3ke9AV68XgdegLE2nTzp+3+KKpIPfAec6J4Q
13JaRCLWZeJZcsD9pCypxnyGcaZaiXCg2VpV30Y68Qf7HHJsgU4TGNyQKURt67jC
Y+jhJSgZVqKMgbLmYHG3c9m2yd2GAyPP4DWRTtx+RdQkPw0DXDygiZM1BylvP453
h6uN7kf9rwkt7wVrZRYrOuqnmLZbjpmLSLaakVPWZwCIOE14m8XAIiOBYD7DZSME
L+OeR2qY+Eh2Sp3Rcklgu1XiwZXMqmSuX/vOJq8/3PptKkrWgtMW0VOk63IptOgB
eqxgiBHCmbcASgYZrnx59CI8x/wJjfEg5IsFADF+uGHsf4/LtNIbKyxulRJ+as+T
MKym54VlrbFlJpnM3F+pzTD+4eS+ULmgUItzV0Le+fNDah/pD6ssWE85nIfHgLdp
YaUvpMBZMNJmfdEwBzvlftgN6IfoWZu1lSriJUitA08i+RcmVw2r87Oj2XsBL+S5
aeyvL0v787g9T0Tsu7XQJ6YnO+Zzehfk+I0FqTTzh/k//WKpOohDx7rxvla8TKm7
kYa7Epjszjisih+2UcTTv+DQEniKEwyZZFkhoqHF0nUZ+0CzRNdlgWE/rtRfLxCq
e5IfDxUKH/vpW2BxpevfTYC3nXaqgl7vIX2bPipC7Qw5ZV5mYtYSlsWn2qGGQavz
qRHdZY+wUS72BbnrqP6zoXReNKL7X/bdoGXlWPDw6o/1ADZtUH/uetIRR1ncAwiP
r0us7uATrwmcH79KBaW6wVwa2HUfWgWyg9JXqd/0qW4i7I4w283X7ZITi/9gydW6
FViA4/FuGXSrfPkuway8AnmWa1sTm/pos0NU6PQJO+Tx4QhHhtdL8/KLLidJ8oLU
u0bI2rMcBAHS6aJ2zpM9Ce/qyBuenjTOaNe+SQDx9ADXwcrLgeoo1A5H+pSk4OHN
Ec7JtXQh/u2A23sCnmRSBgEdnX+ymJCv5Mq/oQyxOmoPIJcaBZySCl1uTouIuO40
Sf2fdhZqBD3bgiPGIz6sl48tBFQWzIZ83DX7yjFn1sDr237a/sZbYEvWSPINUenr
uMpF3YlOPpAJAbrU7YFhx/xhzBLegxapgwdJWhHBSwQh6MjKnkWoXbuQxQDZorXb
evEs3OMt6akzbquZrsMh0GW3a+fLkW1DYykZqyPPoH3jt2ii0ODVetKFhIKaXu8W
q8XWX74MQIbVwrbLf/FBONMRQP0zhnGUt8+pATEVestPboFcbpxgExjjm22J03KU
8cCbVUltE3K/ijXlV2+r+K1DVzsBnTqbEOKo06LaLnEYXdIwHM2ynVaNgFVl+ClL
i7UR6IvroQDXAji12DLL26/7VihhTnnGdJohXVyKJuOrM/SEkRBAnCftM+ERD9AW
MATjY9qLpeZT87BTEyMWEcNcw27hBSBKbNkIt9L99cr7NLTUqByLsA1LbmOAwlHi
UKDnM1Yo0L79mqzCBvjStjLmKTlg97zHzBuigREmDygvlr9uOT4zAhFI+4X45zyK
QqzQ4BBQ0jD8QsaNTJMr4+flJ10jM2NXG6sy9ocSZpxvpvEP3setB9ijm8++UBs/
gY1lQlLBRs8rPxVRL3I/+TMfhsBNUm80DMhEx2qBShnfPhSV8WhQHlIgLuNSvf/k
chn4J80Dvf+gpGkTSDhl99/KIqoo1sPVXSG7Y0tjKZdRPkyUW4s0nnGfkLuvYrwr
c5w965WuqTBYKZlyMuSENTf/tor7x+QSRzlIae7gyqTgnZ6Hp6jP8RmiNnQvFrJW
fJDEENfKwVtuMfwdr6dD7sZdX9iKLw7Cgr4O7JHZ8kAyGjJUAbxSM4DgkjVsdsO6
meGGz5r7jQ4g/WSGfJaCauazkHvlks64bgGn+N/QHIKLhc/MRgujFUX/T4Wg/Iwt
JuBGYdZIwlI7bhrrgq8Re453osUOL/u2gwKwncebu7GVouqw5pA4vxZXz+hyZfUw
lDvmfY2cfsSUxWMczGBtPsavv3nqrsXlQIyk3pF1EuPS4shmfhiV5h7UwQEzhxt6
8Cm10hi68MzGD7BeDhFXfqu2tB3UHHal/bASjr7iDpP4CZSfclnZlRiqfOTxsM2j
SKdLGexEJK2x0d4z+AUN4GwN2n16sPU+kUdnmYHjcx+PNZrqsoIb9a4TcQo9Q9aV
eLjeudH8GtCpKwNHkbWWDeiAo3x/hsMZHfbEtvEz2gWWt7OqhkrxNtDU6xy+ckRK
SzquzgHsjwEmSF4ziUMvVJYM+6XZxwN4XjsBUaKyczxSplivqHg65phezkm/6NnI
6wGSIJ0OsGxSNODk8O2TjEtUBSKPPnjP3cH+X5CvuMySiApvG2HXM42zeODmGm64
nUZQpXUTzoqKFVDlfmVUldeiAcP6rEV35u040SXLvrDGAW48wnks37Lr66J7qlSZ
ZVa/hkBZXmlUqjiVJKlUZno35wVqLrQJ6sT1IxnGcjeRzcMN+9UPQt9TjAGV/nRk
N7BA6oJwjsnlHuatSrlndzsO9cNm+4IrjY9OFcFA8cnzXG7OeKiLdZXTNBGddCzm
b3DUfncVp89HIdcpQJ1MThourZkTu2R60fobmCCyiaLOLx/GFTum8RlnSTJG0Mi8
33v6+OmfmldsYB6WRAQbWqoQXBSVvjFu1FppjuOlASgTjqfPEEbzo9MWWyiSJvvR
+JYf7fVtQTXFaacOugSXfxqFXOn8ZoNnLBjqI9v/js3OomjF0m50EhG0/uVI9rSl
JtPu4UEtxlAPbppygBcbVRM7EIUD5lV1H6+9bI5FvNtfbNO1JSof9cjv3wPtl9/p
9PY1WZSgvikd8+hhaZyAmxpy/q5y7Oml9VY8TAHikyotS50dMSdGBhhFn2YpKb3x
De1t9oudvqNeowAnqlklkuo0KpVhMxs4ioyRjq/0JI91WTQXerY+DeCKyEWYcOSD
jnZBXDtUybrIXuhosk95uueYRDIe3iOxC2EoSxBKa5ZDqX9icj/iiWGQ9EsphhJA
PgJ3FZvbbX3gz06G+1KUic1olzVVG2jgxe4zDVBWXrftHGEmnq8h0pscguOOYks/
Exu+HjS+u6vMqVWY6CQLyfp3THtTp7++ZGI/NB/aMojWHDah+mOmMKkCuiLvrkOF
AdBAVbhasBmt85VhKpmb1O1MrIEpFG/S3N2rjz869iXkPvqlOT0zYXBhm/+43UW9
X4O4Obyl0lpQ77IqEVJm8ClNW9jLEnaMzXKz7Ds7sJBKXzoV9dicZE0Hq30VL18a
VgkKTHGJrLkaMCJHGrpGWHX4oMELIzWrAFGzVQq4rYYf6wDW+qq5PxyHc1VnuWA0
lv4jmU9uQVrbGsdDvhAdLmUGizV32zpuZ5WEvuaA3F2ZyHY3MlLgbdppmZEMlYw6
BB4ryrIHjTWAKVjHRwZc9QzosVIvrJVGEAM++E1qDz7yXy8VfwDrlTaiiQL1PT/6
s8tqg2JB2AIZFDabgy6aLhhfUuR5hEnXNcjlJ5aGSNXutHFyoMHtXf2meTgpQSxp
Uu0sMzUOIbIIvkDTCW5aG7IWvYkCG7zJV+/qqO+za0QeAn8u0U3NZFAHmhE0AApn
2AYfpxiY3xNO5vEfyLxLWtx6X2ROmyMymtZI1xFBU3MUYm8MUeYL4C5cn7KUHQKG
TiCcwcVMyyVovGXeSXYCWbceuWH6hbiSrsdLCDyANLIaks7qXX/WXrjKucn4L6vj
g6sGQG8g6r9ca1R0+8Qf4FKdX2H2lUufs6Y4O44pGeHFLrLMkpYmCWD02eSZH8nB
IqQl0xVxczXkZ8EzbtiNBdMzONYm61fQjUxVhXeii7YYRcksqHk64NvJuP0str11
Mv0vhJlAO/wu1kx4m1rjGExvEgo1wz6cwOvA7nAFgmUGPNxLoSxMLkUPIkL2ZB4M
MqG1muGNx6oGkqzGDSN2Ai1/+yGi8uyYf8O+CSG7XYAwqeEa1cmQBdz9j45ni4cM
mZDsQ6R6psTEgABISfZV9sozA5Z4WAhlJKWShPzwK41Cjg6SwPZwf2ck1sawRKYw
b//FbFXqouhaN0z4156K60h9E1T6p6q3Jy69Of3jHnUK17GFWAnzmYExjOx8P7QK
FEN8rVvYwTLVGGGYHYajAOYRtSykWsjJrvv4A6iMhy6lBgn+/Cw/vmlv1mMCbaZm
ZYrjBt9hTCN0S2g1lvOgHNYe5hU39BGPECiFxcE6CG1RnUdtis4QtjQr5zH7sgWb
aObCK1Wxuj4o5HOFF1k0gZBYp9f/OTygKhaVchtZFaQTklTzfjrUJNf5F4gzaVuA
6aPgwKhgvkBY5cd5e16oN9bZGEbx0Omda+7hFq7SapG8fhTujZrWgzdDiOc1Si97
5EOBYYVpnoCWaV+sMnbbCD6SKYO8peXV7oU8RwiZa3Z8XGkUcA3g4XQ2kWKSa6ni
2Ex8mRAnm0Hb9fUc6B5jsVOFodZRT/aVXkcC0dANIN7BjWfhf0BsZziqa/cBXMlO
SJB9WeLnK1oiPwAJ4hZFcHiTKy3i3Yd1dMq97Q8nubRFcvlPkq98SrfsmoGoTNYb
9ulUR/X0e1c/W864QekYjkSRuTsdljxKW/WnOtyupM9mNUAPx9ILq/YXJOeLT5ZL
/mPlWlV0VrtoR7NWAwXAeILXYP9qtaW8ik6hY6ZdSdow6dbhvD6ppsLRN5YpgOcr
oqsmZkL/tw3j6+wPGafCZPEoUV0ru6swTJYVfMKXUDDN85QD3XbMUoZ1IpmPp48J
6GorTHzy+WfxpK21WRTcAXwI1hO+8tYqeaG2Yoe6GtrvrRaf1wiUAchJe63zOLyJ
fhZWk2gT/s69KHCgx5ewSmf4wsg4ne0W9ncmWp+QaULjPHWs8ktJLpQXPkzSIzlf
6rIg2VM1UwyMerEWq5zzM/Ks1KhVMp7UmBLFHcWOZRGYDk4zj9+uq0NDLnS8u8uU
YTI0oSEdQXM4Hi+6R3P+xIbyuUOHK29OPbiEZW8M3Q1ZkyZy/nnao5RHm0iJshSE
bG16bE8RR/GO4Qqt8c1AIFpxPdUzhRwuRvoUXIdU4kZgKnbG+Ifm9RGSZ9H1tFyw
nMzZUgiuDbUUMmbavZAGrI6W47F8JVAW3X95jeAudiEiS/jKmas+ItyPdlJUKjHJ
BbLEyn+c+VxiuboN76U7/+zZCXeT5p5UdugUQlTFtY0SoPhCAwgAp70sTqfnMwLc
01Hwe+8WrB+DWwEG8xNxbJ4lXJ+b+pcMNRORxT1CbMblxfgkGK0BX9AT0s4AX4j2
crVhIhGTLeDYvzswm4rzBLFMZCnWK+8RvwwtQTAnr2KsgSLZ483Myyf5NNYSfVf/
V+MPpvtRcx56amNW6sYc8Y7z+oZtzXbiBUS1NWIxdTsTgufKQMRwR+C5sjHa89Bh
pVTeal4OEJsaJJJD3YwP4he55KrI9MIyaqOcUQCV2srPF8HV9v90XBesq+Cwkmyj
W8QQNjG7ZojDV/oH9G5PGCbOMFi1qv68+l74ot99npcfJbT4Zw4Ed7KGrH6fJP0S
FjTTs7IctIKAx7jiglErUwD/Bxr/7KkRgK4mT5XOxw54uqgOb3EmYlz9s/kG+/0Y
yUdcJEvnApKgpwuuR4iO1ZzRs+LB4CQoE3WtgEc5YnGanJvGMgGYbNH0RzhxiBgM
3vKXxUg1DWVuAXbCWg1ifCQbkl7Bfto40RD2sGeTBOY5HprcsJqTUgTRciVP76+J
P+9Wuh+HuUGzDnS9x2oBRI/Xc26U3qfPQCqR7ivDdYcGNSF6n+I0wWtWnJEEljFL
CjikgxVTnNK5JU+cukL2B65fFjP1iKO49oHGT0lXW9RjD9H3rCRWVUvjIae9+chw
FvymV80veuDzhUt03jIT5lVXY7//wL1X5xkUIgC9BnawLGTCXOCkZwFMvxTMqnMw
TWOs98AmzFphIgYYdVfguAGnJtn7zXCE4TFM34jsQIHHan8qAQlBhSlyLfJ9BXjr
GgRfgrb2O/cYTRMIFU2yDshzF4XvartvnnTGMpNWQVBl/Xy6MI8Mj4K6afFywqDJ
esWJFO4WCTA4ucj1RpjoWo/q4OoLbH6FCJ1bn3syz0KxDOtvkiksllsUC+1sy9rq
uke+/kUPyx95r+kgsBGgJiGCNgJhJtgW/dnsV/Mbi4Z6ucfY2fK2kiY7n8QEnPFL
DsPh0zQHRVnWYXdGx5VyJkNLklcNJuWNu4PFCDZ3Mm4GBjPqZUQtWmPq4ByfehkL
7m1IyWlKkE1iJgZ0CEgpoziAMHmKv9DRbvRkXHMXPPMT+blR+a8M5tsf4RR5fFgO
gSgfCUa5lSGKWPx61t4Sy8UZi8QBL+jLQGRkbWtop73TmTCmBby65Otj7bxngSOQ
YIdTQ8J/6xfgEXZyEIIzP2LVaob8Y4PCQoL70YOwbRdvswk/mF58pNwEVB2Yv/09
Lsq17KO+dI8fOwssyRc/PEqREDClEmLc+9MyqVJULksL6xyPG9vep5p8UXCmESfY
IXhFeokiydBifHbzGbY1tr1PaDMIRK4mJcaWRxtdWAZs3Myr5HN9HCLiVWNub7aD
v3Mz536KFnrq8hQJIPNE3V9MzwJMztmio+oonYswszMzWNkGK+VHA7d2+SkfUAtt
KbWQudnGb9/RQAYGh3TO7b8HUzU/indkKDUsi4ddrbd7xuCm71I7spj//QZOxpPI
F0SoCx8jiq+mXDROu69IHefHCG/KsU1vYLdp/3UwlMHpMAvCB2CM+m+I8khbZoHh
gyLM8AqaCxEXf/T42qzfsLKAcTF53OD4wLtAKxo4/xBULNc7Up2+1oUBgfSuZFpb
FMdLViiX8wBAmyfQ21LM/ruaJ0ZLNBXqKF32en8znv9cKE5s9sQWf/s+9Ihx3QaI
+v4MbDQ1rmWAQ2MCBU7jDeaFCkcnEdFkRVdW0T4L5rOzcmLGO1fBMk5f58yx1G7O
5JnsMDr3Jloh9N+71uYqNh/ibubnTvcmbTiHpUgBRupZKLSCfPTaabuMfSJDsJFW
RltqAXx9X5viSxvv6AsNej6AEQsBYOg+t5FkRhr0MnSVvRM92WREFXsd1vP9goGD
ji+nc5G9UBfNAFs/jsi+vXGArXtsQKDQfzDj+388KVouqvt56krD7hc/7BjtwsyV
MZKR5eS1s9sJkbLS2BgazFOQvix62KF0Ylud852qEru0g4LV7wpOZM8rH9l7svZo
clacv/YfuKNX/3udsDJl20cumHHLfEDDDUPZCsJ+vkvU6I0eRUsLGFGjzKarGxi5
h90cLqvfNQIdvBSpBcBGHqJg/SW4RDhmWdDs5SeDpJNYmcwfzJqdhSAyvi2n4mo9
yv7CKkHNWJfe+kvQ5EU86Fqjugnsr6qZz5tu/PDnGXyNGUr2unk5DNWAPorSuVMY
n0FlvsaS77jWieWocx5baUnr+8VP9Omd+yxh0ISKRtYiFmga8nfIeb4tVKGclDv5
dQSsaiPnf1UAzv22mWplidWXkB0pBtMb86H5ToO3MV/MZhQ447aMcg+oWQWLOgQo
0KzQl4tnzQ/W6vI38VlYfnkLL2MpxzLFBRqsTMJTqwq5zK7nuhns4QME65/rvr1C
KxygrokEa4ONeiQL7FWscz1sn2ZnVDH4+wzCgwAxyRTCHa6WxLIFrQM0X2f8tZHo
6QUpRh3RBX5b8aOWfurjXMbir+sSX2rZh7jWS0YOcDszxX62FZPay3OMFDNhyO2M
GgGKe7ILQRdFH8ilBFJbyxTYeXfxejCYQQVLu+1yW607JX5ATPFmOR+I6iEzYbr1
/1WSs5nrDnzpEbY0iXD4euh1eoDzwen6Ls5KwtqoIybBwg8JNl1GkTdC8AlO25y/
rY1CBeXLlWo5pNnfqzlr0MqzRYPvB6mWW7JYvsW2wUQz2FPuQ97/E6CQsaxRAqhb
ZM6TcY4xnOvNYb7cifVF/Xq445Ui9bdtdgwWGHrQ0PqVKIUd4CgzwO8ETwZtxh/q
KPdczqufi+S7UkCEOA5BdrCiyWBNilqvkwQof/OE53ay3DjSQ13dEGyOGZMSpIdA
Nx2AUWpbqcya8CO3pFRy9Zkr1TjFxd/QuwdcYxObXwwlm7MklZoj5xfBDELfWO/i
h2Dq5AT0VQA/3EdKcZaoHA7Z8dS9JQRnYE841JjoRcpnZiUs6buD36w2t4JehgIP
m42NsWDsJWMg06rSw4yalfcRwn4qj1QNcAw/dDE/QkktAWldpkGj/AG8Q1rC1D7D
0NIcDwGPAafVUM1SMoxnm88TcDie0cPjzC2ltzbVqhY9NBsqxlG1fiG19wbWUJfQ
OYEkhQsl1gync/qO1ofnBa7Hm+mbe1UGpwCvPH4N8F5b0KLjJb7mKMDZfpN/plLv
/bq8WL0VxNa83EZIpxAg3DexhTN7ZBK2o4sW5agjSByvvrm6JKtl70/lzCYNF2oP
dLTx3J6mvEgIQvxJHf9Xqjafru3g2YzpXzT6O3pkYKAE9/wOhlO7hdDP/qZt/hOA
vsIZI2hIqD9Av2KudqprpyNUCETW/4Fx7+BBor0nJ/A5A9Kq5ZoMoXyQAIKTF5MT
v2FSlMNu0yH/BdmuNxbuPpfnWgozPdMuphwZvGVudEnDPjx8z3TKNrEFw/bQIVaU
mZBZey4uUvXV23l+NOhN62L0SKAdFQ6OR0Jg+zefpVx58aK7DEnbtzkAudvPJ3Do
RgIEZVkIgwbqFXVquyLNEB9a2+rn4TjV2tJ77uGMv5v4JzvloJ2yXXCvZXqRLo1p
g8QG60dNtiAG4z/1rH6Pp/7HsMtD6P3boXVB4DV9oF4rok0g4lsfcp6+G32q4Sf0
AM8j2nwm4Pm6UEf7ZYGKVfBhA1oAWV0inCxmYTC96BtIchOuHnXFJVRv5NWX7vc7
f6J3Xkz/UI4sv2tee7D3V7ES+3hhYWkrqLZnscBKRqMo7CAWPrJMRSYkDpaZS8Fu
wsfHO7lsBCpuxfaxTOBYapslqISuzwuRQUfnS5asmIIsawhwwc/yedFXz6e1pIWa
MySf4arAmneKoRsyEVltTcwgcRTDVCW663uLB/Yu/fi38We2Qw04Okdq3FVuwhu/
FFE1XWaIdJgLaRBijsaHNvd+Orp1Yh5I7kJPTXmfYTyVLTvgGacxYn6fYNxtDcun
UODDVeb7D2qAS+IIi88SpsjlIiR58hnzJEVbruxcJcjkHpjl6XrQn1c2Sdk8kZXK
dnr0iobttL94KZS6ZqYHJOgmYiUC2d9XtkdVyilkPrO2E9JQaQHdIs46aLYsmenk
lihPn1U/RWxZ6orvhJztpwPEoj+tfD7SzCqM+CsGFOclqC7dR4CSf2QYZanPd7sf
rYMRTaSkvGYucUcdSazUptRqTB4wzix+mPEQL4c3yMn6w4m+9bgg7rNdzYqC8MB0
YKvUfqlN7ZK5aPU70M1NVAeAFnom7t/zzTdLlDQ8hEvvvpDlhQbodMkQnZSmfUCt
amXUyGQiIEp+A3IuuODCTgDTCzZ0DAr97eDvt42tJVn6gFm3cC+vyppt+3UfLF3u
PZ2MTzVTqfctoBryPwqaoR7WYb6ISiEBiEV0+4vl9l9lths+0kHine/XExc+L20s
fx17lOemIBpaiCfk4GRsq39Sv9sE7GUr6/dOfTV/qLsEten8uW7V4NPmvtiR1zar
9XE9NHvMWlkHqDxRkxRQE3fBDbknw3LZ0Jiuv8NQRi0fBW4qv+Jogg7DO5QOHp2n
4esKImxFEEjaK2wt0V/adBVmvr0dXDtEoOZn1jDhl6EwdQmeSiMYA3olMk40L61a
abKhLjAGuZZ4ynBMFUM63JBn9+KqTB+cH8Z8Va67YygpGPcdVDOe7hQh5wrNTmRs
w9eGvD2Jr8DS/4xcx4WciLV0PHNU/WOfaakzThPYth7HQAN7uw6+D6ROK5j3v0RD
qxdhQ4/Z8AzxRDplMBbYvRKsssxOm6VVeLQcZjtUNpjW8H8dIS9ywe2NYnGlYwX4
bUy8AfGGAapoT8gsHWc0spbfFjkBXqpKnVAztMdc8fMhk1AriACwbLiq5JLWr5SJ
tkOW21z/ezlQctscBdRnMVFe21QV0jIwotshfHtIyeU3hsCQVD4jmJjPFONYDQi8
Uh5QC+54qIrItt/HcVoNcOQFMzzGcLBLQokkgYqfpgDDPA0WyQOJFhZ8fpwckXUh
BMOvWrePKe980HZpljmpe3O5hVCG0FO3ikHCsTugtE4k2551piPtje/Hl3rWzfwh
IGn6UYeOSE12njS7yAIGS6HCCQTICBXX2svpl/9onYolnVR/SxlM2ZXDJL0Eeand
KE1mas54oS73IOtFFYE8kpITePCfjGLsjkKpWVxtZs5lBHYMmaQQzHRVJ1UO5KsT
89HqmNH9/GbQJV+J8ZQMuGrX+rdHThk6lvrNs8gH1GyKLFsnotjN7OeGKD3t1Ffo
ud5QJMlGR2gSvFsTE/N3vt4F7iGyPTNSEpBt0x/d6xvdpXr8r2135XdhiP1u2A1x
ek4NIcRNQwV+yRdruXaZo11UOktS3EmnYjjbF0laTnah7/Ndw+7jHCWUyMlfcHqm
2V8cC0MrY43WNerykhHG0E6JxGIiMmOPjh3xlN6rftTnxI8trzA3v+94MaPTHi3y
bk0pyU9kNrH/mywApd+7fS7wj3dmRweY2sK3QyhGkxfuCwZHT/6RGkZHlEZcT9m9
YqDsufcEtew/hfl+JEoMTwoXg6et8Jhyvw2bnXuzXZjS66ssYrnwoQ5t+R7hXT+z
haCRB3mZRLI/XZ8SPBeBqWRPNxVabwGU2S/JaLdorB3umcoI0Wx8EEaSZVEMfYNJ
O9W/cZDcqNdwfqYEUc5FMdmJ1Kytt9+BlZF1KNmJgce/NYOe1Ejq0aoOhsNgPtZf
xHlXWQ7BnceLZNS4mCQCx7HDytYnoPnLeroTVODRqBIAXL73J3v1fQrHJO7eIbbT
vVwT+2fOlemi5pyHYvl5B6DOWuQK7uqvfzzoNFpeoQi5PA5sFhVdutw7UDAD7enX
rtu5S0l8rMbaVIsd1AtAGBoIzmHWnuR8gjZoXzg6VQsZZD6iexysf44DIYpqqyHB
xnB2Yte1ibgzFcXeqnR5NN/uybJoIq4mQbbImK8x+aP8xDxUGy3AbdK7i0bCLm0l
M+c20C7FDDF1KXRsbhRSPNGNXBr4Gvp14ZcDyrcFsdjXaHDKSp31XLi+W+GhrLob
f94qzu8ccO2j/ZIM7gvdzpDjJN3UsXtzvlOBXwFOwvz4KnKJQLXakHkXbmrtWtVU
tBiVx/4gWc3CiggJs5DKKsIRuNwS5RTaiiWkifnwvSsdLLbTcqqcDq/I75L/X/vc
FA+CY80r+9WVZc08eoMtJfFARqW0a5el/h2j8+RKbJ8LCs7YkiptFoSFJaf4Q2VO
GqbCncF8DsA0GMnV3Rlaxn0xpRouksCEzhyAu1ew/UXS5WkF/YubdENO8olalHKz
WFfCva8yrpJGwon4BPvaStBjoKzkaYvtO4Eap89qx8tZedgNecSh74sG58r4St+/
YUvmP71aO7ramrg+GA7zfLNXsauMtgVNTkwx/XC7vgkqWpHbgpwGTTkK9A+wvsyG
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
JZ50aiuLYkZvTmrSJsFdbnWgIgUxCjz5t0DT7dCvZxHvDALJgmGlaP/w9W4RrKUv
CPyZNn6L7oQA0WTiT8kcKKiSrUOaImz6jmtb8baxgKbGQVFSg58ivuyJHI8LYC8N
vH1FldeW4Ery3hTBhdv66O1YNH++xEQggtTmE9He+A88buxRB5M4NrwuwYcENsxk
XqcXH3tDIl+KcG/9X/ZMSe+gcne86lhonDDKn5Wu88k4uP7YjinAo+3mqjkmcGUO
sNn3IEdK9g1USu4KVpqEMS8tCPgJ54ty3WSdS+gegmBQhb7nBQ73vs1iALVVLRch
ityicVVrXux1AA2j2zToqfeJlLOFe1/uCVuxkyjvMIw9kUMLfpH7glmGVB5D4eNo
TIjYTKjUqytEAS0BdhxO8Mm/NBhrajcTNLhMfzaf1E7h1z0LqyDtMdxtyDOYDE10
TgGbGwVYhsRIsUEh5hHOVfQiY7vIKtWws70Y4erMN0TVQq3J+6l1Ao4JF/AtI+7j
pV3lSp9xoeTAqEnt6Fo/+zMyYcKQkR54KdGAR+dRygepam7Ps+q214xv05cn/tMM
f15Mncq6yfl/tjiPujZJNuouvoRdDiudpu0ccY+4wfGeeBh2w0Ln9a+/GAWZdwMa
sM9NFuHPofqsFBqZoRJFkPc4Yr5CrL+LKEFjFdSRFfHHxr9X0A/eKUM51Nw13EMa
gMxLVt4VRcGcut+EJrd/upPwLglCQeJ8dYlp5000KHr/ip4b0C94Hwuf+YdKNLJ9
F0BgygR12w1b8FeMBPFwR2H038FuXgvVBQmdHfVTEcW95uPNbxbQUTcZUJuQKjTk
ayNxDd9IOhdp5OwW9CL+1/kZd+BAJjk04V03FYwA0xVtIGu7Bf3Mdbxsf11P4ArC
Q4huyo6IPduDgAYSq7TSssghSiwMgKtTdFrl10Ucktiigc8dCXkp+Ix1fFCNBp2v
jvnJWIgLllK484hexfCR94ln34e5DFC6KnN83OKsUz9/3bs0g9VuXrUSNMLEwgF3
1jn/gGxEvxZFwLtQGqUSx5jjDJJusjGkfMxKRw7it1LeKYpR70e650UE1BnlOdkv
sUJWkWHXt0MdQ4SDq1C5PsEi6inKKhGd7X26g7kScJZSUYaw9biTMIk6q43WS7Vh
23qDORbS0KaHZdGg3RWdkmcpe2PW/r0jv9C6QWE0y7ZN9qlyUfvZQCdWiUE/48za
UHg0N3foksKnukI6hd/QitJ+xDJXW057ugS2gWx1S2eD6p0cPbJBNHINI2OBtfh/
rJfcgqf415bltyAa6Zn3vQ/RUNgRskplOz/AelcNYA0y5nQuSR4/fg3CrztskKOI
enfyE9FgyHiSmkRZH5LLjo2/60JLveGBYj0csBQ8o3i1QMRdIYhzFybLNV8I84qe
6IeyShyxX5UZtZSDkYwdTIselWqRuQRRt13akZSYExV84kwQCoTp3tMuf8LUBGEp
t76ElEVaZm23wXpFuOU/aOTyjtvVDmICJbNdR8sC1zlce20W135pB+SwsOGmWPYp
RcTWTWojrqOuecG+OSAOgqObLuYzmwPRlloavuLPW/+SuKXGmvzNMrZEJt5XrRKr
kYJYnkdxAmY5AlyAikZWGJRf0cxFbLvSq+ZFCCXLSJ8W5GRsYCvDgQTQc7/GSpIr
KtoHo+Y6F8BTqh6j+4Q70u4KmDbbrDGSP9PgnBRWgBhXQE5YMlDGsvmgfpeD3Mms
UVbEca5cig/7fbIo50P9SDT36MK0tE6tsYXrWAD2f3YPK5l8CeZAKnDoCrSPN72F
1nfAKO5r/v6K8gMwtzPlV4Ejfjv8hJJHuRoLnV6t82epLb2kuH1kMA2/zFqN2rCU
FwdJ0UXnH+yjOGONQdA3Wbd2KKY6yHBw5L9AHYeOARyOr5RE2Us7rNSVCkwJyuW3
9/4MyEns49CalgV+WHEORfxffrGqXEbOb80wcaQ4EfugS2E2pk/FcKnEMPq9C00Q
lBX2ryhHoHVvxHLnXMWnqRn2ODtntWhd5gTNlu8EI3ZX6UkHFTHeCvwgsMxDmLDW
vlxlldHMdIYvSFycJ46JpwBnotC+8tevHY+qFE1aiXcM+wR7TVJJzFrtJpqDbvn4
kZI7Nludl2toXYk7Nj5nBwx5Pt+xpao+YUS82C1EsKktwivUWu543pgzTILyNG8c
XHu4hBv/t/yPFwQyH4Chmy4qqVezAFGZ7SiGxPqK4dY0DtOYtHEKrJi67dBLGDLd
qIhbS78pMyRvRc6mH96ms9Mi6obMQs+CeERuXaSwRf7FxOVjmfIsKwCiE15C/mph
wsK4RDAWe4zHA50duNTj2HfszFnjzWMm0y+T4kZfYEzxpl00wwARTb5GDOEq1tmT
YD0BFgMS1gYhU7A2MORow11W/MFKzmUiskdjqGn8ogPwVS05jwmutLVCEZXVJ24k
D7MpaxGHuK5Td5PgpMmewVQMKglxl59BUP7tVTACRBrQAHOxJSMPLZCNGSJl7+TE
Te9pE1Kpxtsz5aMEVufuD2RsDF7EhovQXtt5wjTi5pZvIda3H/i94xJQo4EKAHLZ
3iYpprPwpsBy/EiOEn6aPU68w/M4mrNWCknbC8uOv8WZ0/sI5odQm1WQgIlcwO3b
kMWyN/tmugC0Kmhpr4574jaL+cH0LVl5MqUT5BHcNrCPygEyS5hyF7bKE/jTUI0h
DvLO1EMoGqG8J2W51SQofhq5tol47WPUlaIszqyFkAoXq+ri3QAg35r7zFxDGFRJ
OdLNAHz4516+Fbax6axed7WU97mCWTDtxcePeqLtAvko63X4aJxiifNRxSi2cyxE
eVzUvKFpOqRhlOvytgR1LgL69St/U7a/ujVKJbYIn9Z7jKvMbmfKvVz7CEHgE/Hh
3EjVPNX+3Q9oSTlAeh8ix9tbf4QhZQ/+LonmCag+9l81YqYf4l/yczqUCdFcm3vT
dB9SXijTqjgVO8p+oZajiECxGPTC3NWzPjf7Pu5m3l/qycRKCVL8NodXb+bo6woI
lOVNe+hE7dpx8ZwxmHUSSth2JP+MDJCtdb886wwTiZv480rFCv+ADPYxowscnY6s
UWqvPlmsG3L2gcld7bSJj3ThRWp7USiM6rD9jJakexBdFzfOyTiPRiXMF8c272nU
f6qntDnHw+ECn2KZ75T2zkUxebMN00EVL0ZeJvRCyJGQyotkSHRuuCHkwsxRnwVF
cC0d8ck8n7PI8hfnDf3tzTbh78rDuwfOf5OjS2gCydQOlbh1BdFDND2F4pWnML+6
qGdNHOefd8f/coA5Nl35qMtRLvVSMfK/n9BWbrWtYpvdCbFqE3C5cRiujmA6d/2+
VogOemU7LUgA/2EpQ7A2MAE8Df84L00yb5h8xpf0xCJZw8ixK7ObEZmKbDbj1uz7
9gO54tLp0DcMNqvhU43TKzluNCCPzG95LmAMNRT0TgMgw/GRJIRjFcJmBjrWGVRi
nkr7+ZFCiABPx5Ljo7yb8NpwrD6Fxc5/JjjrYczStGVDoZMIGe5wFQniW5G10EvF
h3TMyoBzoUc+R5mqgyg9PKkW4OuyZf6EikT58s2VbDW4vRmtrfOo/G27EjbPVXzI
hV2ZKSEtnosLMWK2OkBeEBxFtnwO1kpVa3Hk85OCstu75Te5k2R0eufx2ViztgPM
5kFOU4dCAzKv+d/Z23cWt04Znni+HkFxKCLGYcUJxMhxgaZyz/JGvr/0Dp2F/M3S
1VhVHdjITdwqg7/Sl2psg5Y5DhfPlnHxQuIP46WGx+4BL00sSJuPjg9JlVbNI4oU
22GTpvZDvBJaWLQwLReWJhlH1jj3pHcgDdAIrPdC9EW5zJ3suEQp18geM8kkEMNR
gXboYgdeP9AcVzAZyThSdnw3n8syHq8kwcPmkLMKUFh5pq1HS2IqSik0cFOBGRP5
gnCh9mpNzlg67pY+AzeLBkaU85GCGMAdRzui22x2zbUOcCjaJlbK48Qv9ubQs7EN
0I3LxKYVn8VsckkEoNZsE9THjI9E8IQ2i9nGtQEFrs4XM5ftp0u0422szBoQVRQM
bZSJ4ONwLjv6AnDhP7eOZX2F+p1xq1DNjXArO86H5h8iVhzB+a/7uUCBkDBTVSrH
/qyG5jXtql3l/T8cEkkSpmCUL2QdseXQ2CN89r3Etfu9foMtl4c8UCFQQ9pbpfUl
KSEcmGsKd9QQrhG7RbbjUIdqhUWiSL7DEDayNCmkh4cnq+p6E7LELKxn2gwIiOC9
o/OmwzQO6kFulyoyAv0Su2hSpCxdQ8HAOw/YFwXR1zdDcTO+CNgkr1c3Jj29wLtk
VkCGDsof8GEqJ+qte2LRdSBXKu1mHmxytgwMbJ0fwN8xbYcl5/GbZsLcokU1GDPD
22BZlnNrcMF6cH+T8yECa7j4Quhdsmth/Nb+f9Tz0R8f/T4j8Y1e0QNMEk6OVKBb
5ZBQH0TqswTcyyTs2810XGl+BOHQWdDmD1k00XDz0ksV54P63ttJ/NIbXok2k6OK
bGoP8+FHXsNxBYihBRp5gz4ZwRPs/qmLG30lwXh5WOTDgO+GZXWDsrlh36j6TDmr
mt7rDzLsPj00lpE+vf9VH4od/FBoOA1AKLTd+3BtFFt5ZAw7U+ykvUCmDowyVepS
g8Co/tJDkboc83uapImp/WEh0bV84GFxEbJj1YQjUx7PTsUK7H7QnbyXf74V/XgA
G5ewNrELhV+0tCQuk/7Bef1rtv+p9Yag0zRywmBkPDOgO755VgshYb0mybkfQd7d
qUc8ugwJA4Dsg1D39Ji7uBXvGiIMzb7ywIbJOOJEzifrwB/BvOQ5fuoixy8TZ9Hv
KvRSLnA5wli2kE1XRDsWMNgk/YKgAPhSFQ242sepS1W37BaHm6ldrp8zo1wMmNVH
xUmuP8dgx9IDYXCQwc3prBsgSzFxsQgmks3ENL7p8sAETfN6PRxe+aAhOuaens7f
7t3ChNfLUovChDZpIFDUho53xmZvZ/Cc7B2HPuvrb5kDOaM73tNIM8j8kRQCO7L4
RZX2jfNWVeMe4MlifTjfkNBYJZ/L5J9hrnZsJrY8hUQY014O5JtwF3V6B6SpBXab
ljRL6Ry4dKqQ2eKlvrAjdELZHUNrtZaurkfXmvKjSvqRqROmzFBiPYQcjXOBQFai
ZsqeHN7Jc9I8DeN3y9gK2cbkT9Z2c2QUG14Z9k/43o/8Hyw2X2RbRo2g3MDAZiSI
UvhpSt5sKRK/LBpXbhlZl/SrF40NQkeNScwWSpouviAdG6nRdf9K1sRD5eBepQTg
YC7DhNNE/poHmDcr7YtstFOT0PKMcRHOcSshxRx8Bklg0UD9ItuNlL3uGKePDzul
BWPpJx2WZ68elWc9D8Ac4W7ANQGCRrUzvLGGMEntNvTbjWiLyyZsFEPWaJJ/0oPy
/e79GlvFn7NTg6pVaKdlXBDx9JEpohle+WFIwLoFZmuLkAwHOYZai9N18l8uV+A9
gZzdsT00R0l7XCQzn5yhoM/+J9pLqOQVZY6MxQMJUWGOAclU6G5A/JHYSPLMgglb
wgPFTP3dQ1LwFciqtC3RDyfuYLsJ4YV9n8ZVWew6WFqpe8oWu5ojeqx/HUfHcFvr
BONsTvlAZay3CBPyfYsws1O98kQ+fASVEwEHfsYkGdWjmNGr+19mqddjepvyDZzt
+xvmDcRNZ/wGRIvM3nna/LPRFKCgFOknGXf234+s03npegESkY5pM3M3GlX7rC7Z
Gkv78/0NMCQLfR4x9Uwl7UwlWje5gcM2FHPAee8ru1h+und9wVONXXrPB1Sb/k/l
81uLygJlVtasDnn/4A0MG3g/gxsDU2Q1FpNRcL9Goz35nVf0E9tqfCLzXGgZw+Dr
CnL7cph99LXcTdms7P8f3Mcu1xcspSzK72hF5R/ooTjAx5LkgBmxLSc4ygOP2eaZ
tnxaLq+hZEQYtS/ZcnnLl9DprNj8CSeujtdZsmq+CgYoZACU1yubQwRB0a+S7V+C
jSSz4q7jZvGEQPbINFCJz3nrqixG0V63R6xkIHs8JZIBImH9AKa+yFWpBzKkBTip
5l3Ys8VeWUV0shFTyEEzLAQ5Bt6yPRADOpzP1Zz65lj7ZlbKTBvLQMAsBBMmHqGi
IOvlDMqhkvGCgLzpxYeWIAVfffzBgA/a7ofFit0GGbDjyJMaHOBjy8c6y5Hxfzbf
psJM54KwDhlgBLkyrKe+1+iYyiulzwJ9IrTtXj0FkYR7rnT9/zsbrMKmBUgKl4Nf
DR04j7e69G9h9SuR8eYQH9b25fp3DKTw2M8CrCCudcZJ1EMKOVVIvrf35BneQxkk
vx918O+82BZ+GXBPG45M2L4wAW5VxsqJlqbXQqRqEtoA5vyzj/HaeTLESjLE7x/k
SokYmhkL2WOHTH+ZtMFWpaePU1jgl9l6tSwly1NR4sHObP8zwKQPv+2RI7osamTw
IOnC9V+rxinRzDm1c0CylxpHM5kcftlRw4NuwHxD9srYp/p5Q1PJpGjIqwKllXli
sl8NKaw/pPbE3SwpR4BWURehT/MRNCXep4Fcx2x3pVyeiaYZbj+JsojqyPIvyIDI
eVM2q3TR3xjwKFmygU0LEBETzuGOrH1sXngvibyelIIU1n6MuwFG89VWlm1Zde29
qeROjz+tlOsCVPldLaVpeWOhPsjZz/PwAk88NBafOV/XAhhRbxOvt9Xb3ZiNJFxo
2cX2H8IEH+qC6iAxbsZiikz17m3PJ5yChdMy2J+WImZAHEfdLa+O79AR29qHADzx
gXI+oo2392Jk8Ss7Vzy1DttQar2ustpXNOcZY/dW5x2ugtt/s1GnvHyWotFP8hLQ
p4N2MOJC2AQQzT1fSf1KcqB0Glk1Awou5JvgXr7TeN1tlDDg7yK/WMnQyuma8xMk
Jp549q4EWQqTC0S2rKzTxxBDgPUpvsHomiokSbwC7nawwOPmST33VU7kQ+sASYRd
ql8pION/QdrGNDxWnxEbcJlp6C2gZvXIGxCgQjj0jiwnLeiRgygIGIjYKG8LuV6p
2kUgfYInPMF07jQzF34flCHaCNHMI+lRfmi+hs5cDLhjySzZgoRjmjIs53c+q2dp
a0xUGMZDGgmYFvF6wdewLEADGK6QyyS6q/FHswBDjiH5WwGydL8HJFSzo3ySfW/n
PvIEU04GTNyDbX+X3uTsWgYu/LaA0EmSn4vK5gdYML8RGvq7au8jwxcRQnf7q++/
4L+N9FpfAgJ+7FL0CiZIlj6j/+MPPZkoPoCxVFLIVGiICh0YXVo0Gik2xTMAp03i
+bluqvQ99bpTnevfjVNJmHqMFnnzl9I8jTDqE0evEqmfz9wbnl1LDI+EZ6UWR6ji
SZ0vYYOAYKR3Br5kXptr4yuwOpk7DPkh5Xe6V4zmbWhxbDvuk5H5zMu0+/NQJeOl
yblm2iMzc0NalcMRKd+3W6fCoIv6qSL0oxxSPbfl+Rb8I/KN9MXPjAZHEW+ki/Pk
GoMZIEhWoeD33uvatGZLLfy2nDnPvksZXA1b3wJO8tnw5oBP3cKmMENEkvaVyvb3
2vMMusSrAhjORzD0Y4+cgOCYSjktuSfPUH0ZNdBSuWR0VsAzMSnsZVErZZ24+Dp5
03itQkDKifutEuYYOG1YZAAes8d10dGzAi5oEZZQp84OAkkLF9wa9zL6f8UhSCaG
eQd+kIJl5B1Dl959ks/i7YgR6gc4lHyy4QH8556PVcyNWprXK2EhwKuCs4YLplYt
cNLiyyruqOah+ghKdekgV6rI/acaMf0AkczWwJLtEzMsihOfsGtGx0Z4xgPhUu94
6PYeR6H1LJm2YY0WVun7dRXCHMYLqbcWmo5Mo4FfCKoxq60O7xzpacz+bagHkB7X
BO2lhG2kZHZjeEWNhNsASCtAky0reTgP4YafokSGC8m8neXPEdJRfTEn6vSgbn44
yE+kJlHfYc+51LlB1v8zceySanutaBylcvVzQN1Ja6KYVuh8pJRxa4Ahpnsm0/kd
EgXYeamOmz6n6vyD6bjjLqsQERml59iERT3z/ihMAaKhyud91Ol+yKeGFZRxQ9Hq
ezd6VDZDlV4OFPVIddvwjXhkgyiH7xvsLjCfuyKEuSwqtQ/NGyTcGyDYljWVKxeg
YXuGR6EOC+1iOX2QTzw4pzDgpmmQAe8bWhhuzRZ+aC+WiY0AJ6ktbDdR64+H61Zg
Dy/rQ5j3+H/NWk5FbnHFmOI+siLSoxAROk0E6hsz9j6TYOe5ifJPtMaIZkLHRzCE
gjQhhy2fyVsIH2RWXtfN1Gzo9IuDqWPJ49E00wBfh5R0AY75laDCfpuSS+zNzVa6
6wRZn1ROUfvCH6B1Tl2+G1TNesCrUf65fghEG133YyC26ji3JVJ8+MnbLYc21OYV
knKBD1BrqEfJTbLDA2bzxxKtTlMC+8oF7LzDTPVOLmxepgrY/8+uKiuot8acnqhp
M98kVSKpEo6V9ueQ20h0wg7MKOak9FpGM9fcTSg02GC3IWMxsXFwl+gTUnCuAHHK
JaMC7MTHHIjs9nXl8QcePUcNCksU/SZ7YWEXMTug3ferVCpCqpadlDbqihCNkiKr
OrmKlXCxsu1fvejAJ9pjUEHQMb+g3vnQ490Is9MJ6o3m4fFKVRQfEPoB8ZIy1OX+
+4DCPmEOqb8XQ/UNrtmbmB9uud0YQnMcAVg+sMIszeeGxDm1ugRUkTewc/+7b0wo
sj3KN3XEsdJ9eGExcVUxC7+W++Ex2Tc3inAdLABgx3n//PE7i0VpjyF6hQuP1gbO
LypIoomg8kl+zCz+ClN5Q01UJJvjULNAQLc0Pf5adICj/cNFII+maNY8ApIk1Em0
cQNgNfNCPyChxkscA9SPo/YcOQpHdtipY7zbo5m7NP3suc6Js2QqIXwZ1nWKd/Qp
n33ZkxDXgOh03GOVjyGoa+W5d1pXonOZvol8oCUYRUloZ10V7COYjoi9p4rHl0Qo
8LmX6b3eFvlSGFsNcmCiDyRD+PQoCrz3c1KFvwkJSL6Dmb6oYMDHX9Y0PJtMSx+X
4/Aws2OFLarEzIcpfZWAJcSvb5T6Ye+wA8dd+Ad+y2d1xsGQMAFkoguk8sFEIzrC
qcmXR9aUAaw4s7SDNdP3FtJ0xWPMhjSnGiI906j3sl2CLS9IsJBDFUP2E7ZzT7IE
g1a7fSHd0hWu8FrPuxl5J22WElu5/yicmBHCBDYse4wNHCIQFpKGQ8Tz7eAabVHd
hjLRjGPFAb6HmtEtV3hfcmHFn2daEvgTB+5frB5lIJfW9+Gh/vjEf7yzgOeYABry
yVoX8aqyKWUNkV2tu/CDKWKpOKJCFh+Tg3sEV4Ly8fWR5ElA7M+LSTRJMNOmVvzx
Un4uiG0gPG+tdaXZmg80j25a45qVnD7KhNYKI15pVDX3X7jxqVvCZmLjH9qH32g7
scqx+4IWoURJ18tmy3lgw/2cM9sO2093CPp9PBBi3VvDGNb4fndqeIET7eTGlW0v
5Ppe28ONZ6kCXA2TBGe1pAkQP75H2t3fYd1cDuPowf03dlXTawMQwIkIBLp+uUL+
HQI5eceM78dLpZwcV7SEe0WOF5qkdc3ByWgTxiNo3awF7zGiiDa6DNULcsik6SRD
Mpjd44eEmQee5mAKqGPF5p1arujnWaY9qg0OIw7q4tJ+6yIEpmKTa2CKAOLFN9uk
NpvL1yq7dmvceE3zIAi025LxrB5U1n8ioHkjDgeX0ZxE/abOAkKl+zIzchUkQkKY
XH4GG0mRuN8dwV2rkIABvPwddjN5nWBElPrhk736310jioLPFQkJtJfA4HNjhQws
RjSCTgerEqq5GVbvZDWgstbmiyyWjgmA0n9Gcfwqt3Fep2f4+s+Hq38zd77NIhBc
aXRrSVczQSaUwT6iVRMMksib8NHbGsHUNOAJYt6TVZUevTW3zUlZf6WuqB5dGnBR
l9jtZuNLWpeeGsRwA0w+Q2Foae5QDMukoC+5dVr8MnFu+uwqzw8nNHrqqCvkbOn8
BjLWCwjFh9p/PgPWrkspqG25jN0YGjFxivN1gVDc09PjTHknL/zeT74HZ5C94Rip
iC2tsaoNFKqmrHH/+We8T60Ea7VaEIITTQ5MpccIOFFltV3zco4ReL3hBVRg4j3x
9kwVlC2QeEwGHPPjbxrUKP2cHFi1VRv5dcMh5VTWSlIlEQxJ7wFuwV+QRUJOe04w
AQTFxbIMOH75ylb4qTbbqPYNUxK4JrppNjlHu8BEv14SCAgTA1S1VWSlYI0jGLBb
2EKGPtAx2fBSa/H9iXkboK9ieV837rqBf+bOpt7UbrPePpsDC6mcCuVhiosrsBaw
Yyz43CiClxnzR6BrFLsS0YEsaJqIy++w1FVjQd16Zo4DM3yrH/99BqvFMXmc5/EL
TIVk8h+wc9x490sevJNjpEyKaBGnS4CuLOO4P0jmZBHgLp9sogt59px7bWgKVub6
7xFzXqRgQ0444RwgU/U4qFF24sANPwWUi1y0JhgPR6P0GQsffRzV7ZFODyjquKaa
Y65HKuQIZmwcSxOZFVUh9dLMB+lPz9rntlmrZnCjed4yxpS6+AoBvScFTnIRf4Y1
WrF9xRX0IuPJCyfdltDPTeICRNwOAtx5WDUqXlnEM8h3z+QR0wRDoMGmWtiy+/0Q
B5d993ivucnCDFLtJj7G3Vz6J28gqqoF9EqtOWkH0PfPAYYo6NWTGzWgGbv8SBnW
K72ceftSe+8ZLslzhY1V9jWO0uNickH60DZe/RegNIXF2Q+qcUsknieTAkXApqGv
lVHRyLqG5Yl8MBNuBZMQ3Pd91EVPHsye4XVieIGKsf1OqQlzmqHKRMaejQAoEhku
MQTkNSLhvHtW5xMBRGW+JbgdQyof5aGs3sbwg4Jf7adwKb7JOVpvwVzbYjOBwvet
6gS4lWMU9HG6ScZvObhdfNv6AyaBN4cdezUE2Sh5yfGoZloyN3EFSL62t6rbduIF
VvhM26ZowD79oIZLfQX7pnAWh9O7mS4PVwIFDIFdQMxLmXB/Fio1RWCegrhrc+6s
bUfMsIF8zBkB7umdSL66GbUVDXUxfoXZJGV5umTmX4Yionj8aV0mVYsDBBb7TAN/
hbpoeQdehjhGG0FmSH1WATrPUvVb2QzNXsLn+qwsoPDBdwW/oVY99QkDMSgX1t7b
vnLB6Y5Bb6+ElLfAytzKZcd0kyUu9AswPg93UPaVpIR+Gu3RZ1uIyFJcXJ3FFuno
31uXg3dKDMia7cHjDiWlhCY4BZpht9UaS0baSRKYaz41jrVuLP8tBJ4cm0xHKVrR
DQwux4K7I4eNCf1OYDiHr//Q9XdZh5yaM1FhwtPQXVE1FAaVvsopKpxrYaC74mUq
F8l0nRi0zYGIQ7sneKHl5ojKR64yXA9YgllfD88iXhqXr1cEstKGP3oMvrmJJYHe
R+C96OSo23NXakbjdq3yy/fxRSOYgE7JrfkoLpQNL/IdAEaJJD1nj7Vvj+w6xWfm
CshxTKhDpeAUk2F+7F6TKXzmhjZOgt6FOhjJAwj1IKbIiRvQl80sL7O3bWo8ALap
u1rfj0lVs59u6SskxksRPz6M5PTk/auTxIQk5I1A5GT8EwYSCirnJqdqHpfrIqMt
1R8TQldYG6aDkFjSD1KIG8w9waCTmdzROxOjSxefz6YAN5Roq5/18uM3rJ0Lm5nW
Q/rVWF7KQWjHex+vBgSaJeSfE7TDVR2Qgf2jC1p2t+X7fSwRjX2iBx+phdbxfeII
dMfAg/wIErR0n0HB728tJYIkBC/R+HYy+yV6URB7KATrmYuMQdR9yQAnyWUcL6Ng
gc+CTZ58Pa86GbdAPXnOkcwG0XDewdSI1R2pfc/2kMFjBNKxIMNtWZV+3Vte1rnj
FqAyIxJlpGbGFEquagk6ChumpsLsm4Nytebn+FxH91pbwPOibkWLQbMttHlpPUMi
r6LyrXBoJA46jYRNRm4K0dMNxwARfzEHbCV4IXxjXxgR3C3UnrWF3jfGRKnhQqVm
d+e6rK3idSetLt/svHvfF/iE0A+dCB5qWvUHhiqoXEpIJrshcvqsQ1PhfPggUan/
Rk8vLDIM+hsnmv4VCaPXPOzOkcHKvVMVIc9NrjO9JsbG7NmFoJHYa9RWZNxV5wjB
j46d5XplrwN6+FpAf+WTb3coZzWiLbPE6WDSJT/0HQlWTROcL4+g4LeFA+ofBFfq
5geqhaU2lA0RUt15h7A0+ElBVPEop2i4TyNqZC3wzObbkIMUiR1h4dipm/VgD0+Q
u9L9Y/B7vMYt1ragJLcwLqxTjIpWMdl47u4/BjFyizCPjZPXcE8VR7/gt+2Amk3R
gmjWsDEBQrSmiVhmbkLRG+ZQYc3aAGB/3EizZu95EwQaPNt8tigszrDfboWY0I3F
Xvja26AdOUbCsTXHr1wQgHgUnpKBo1BAqeqPSkHBJ3RZ1S73RtbWQRqV2DcuhhAR
Gr/hA3G+L+oCiWpHsfI714E3OjG1/DF7z5IMegCDIfNV1U312oxaB+rYPIZ8D8TW
Ev82ycYPc22dgb3r5bvcKr9JvQoWxAIxRY268C8n7yGbzCW3d4GM7Zk25IXgs4zZ
REuhyAMLVrWfmzn0j6KVesKDFVbr5t4jqXEKQ+kB+llaM+fjtBI6y2ToldBpkwsr
ZAeKmtZOhtMhdbKGTtCe4OQc2kT5Q8xEwais0we3ZKSQqbCWuchq/D2ViCpv5x/2
ET6QM90aJIliX0CPtVZklbARe4vbbwgUM6kLiXlFlU19Rn7K5zmuZCIB1yRRgJ1t
WYOzsDUwvlyS5iqzuiAZ7IIPyL83fkXMpZFcssyng/dtAzfi42UG3qiDLjF+qF/+
ffixWMHaXnIbIpH07D3mfKemebxMJDy9KWVM2gsfsT7wCpEKtd7Fp6YdMBZPJNgj
cnSh91XSklpImU6SQtUxbBAWmxqLzxucPqInABS+y/Ey5vaPjoKs0GlKqYMDpety
jX0l0tz2+T5KrBAcA8HfLiJwe+h1ksLb9mPYnlQoHSTl26wb3oXNxkDrL6uVT+Br
pvIA8twJqhFMqDiFRVmSR/1yu4MDaP9pkmTHt7WpP1OSwJC0VRaRSNFteEQB+Zyc
G06zkqIQ2SEKYnvHepMRCe03vlMu2PZNybNj52sJA0cIXiwQ3Wwm5O+ve2kYgVix
F7TaiSuqSXUerLkRohpZ3ziPohYeCP+fa2SBSWPTOxcqvrb8Sd7Eks1GxBLcRO79
6EWwvw7JGMIRGBR5iFrcWCgXIbK5+E1pSRO09pr1r4S5qMiRYL3P0yeo+dFgyDJb
DX8wDe4wSf+fL3Mgepd8RQAcwLYkrz8SOr9l1v1s1YVJxy+PllpqoSWb0UHS0gjt
Kb31XAsr1R5rgQW5Ok5HRt8PeHYKHlIXbZgIEgL9o/i4x9xDaDwrZTsArCxXPQxW
AU0MbmhQRIZAgSnemSWFzwJ/mKyvgalcq+c6B7Mg7AZ5sNgj8uaZdbjNQqalJqgd
MZhbPnJl7ZFajGHOZ80lYunFmsif/Mf6MmPSImXYVfMkHbCFqaY0TUft2a6o6YHI
munphjBd/2l32ZrYBzxoHMNg5pM6oWz3uvLiw7MlxScmn5nTrd7FV0ry3C6RR5QI
aOe6+2tSm7cqsKdhucl7On6akn/6L0QGAQlEVVCFFq0teuZ+wEl1qB4LEkKJcbfC
S38vDjnvani70SCXioFGYOr8/66oBscIs1cDsFHcASux4xZBc6TYPlVU6v5B1bGa
39UVHO5SBg/4C4SKZN3fxxnESMB5Yyb3fPg3OvA7IaspCfMxL2nNqGTl/wqTpvxG
tAx12+7O6UBwH9lFKh9UVGHNLzZDq61SCwhwkwUwz1h52lM5ayOYVToG1Dkuo15r
1sMb+CqJUJiSgZeArfURyYK6nO8shAXykucMJKmljSaeMxop4+5Oyyy9I0wpDg3n
Hn6qRPGgcC91vWpW4W1fEV3dDi1aRWkB+oS2CzmxV8NgWRoggweJ31Ntg/LDEQia
75JJq0hKhy8qvWF7H7NKzCei372C3y9bplR9/UHe6nDYx1YptJOn1KjRCVBQncFs
vAPTLjAxD85lqCQ6pAtbTYnA6NTFN3111iYFevRiqJJJpu5bviSJDg91m1/4gvVk
+ffPSFDRte0qgoD+qoM+WyQmHdvEfC1l+8c9QK3n2SCEkEQTXuXXSI0Z/LC8/mrP
PML7Dy9JoQ5KTeIbq04JUHjMQeGT75Pw6+ETN2L+IKVEDSGsDkpRuLGwt4lB80Gt
WN9HyxZEzswjG7JYoh7MbcbEPpQPnufgwNpa1yaMEfBTTeZgMFYC4dQW5IIlHSmr
UHf/alJGNqaPdn2KlD6KxlR0nI6ejxtIG1P5w+0kyHcjt2tsrmH/aoHiyISDcQxN
NEH3TarExq9YodnPIaKmysX+D6rMy0uDdDE+1wcxySMN4InG6nmJMhDeOzEdjgMR
EdzE9WjX+5y6kK+QJ903tFwCfU0twwBxAO4mnKMUsDtQKmI/Xgeb/VBPpO+zoN1i
CLpNJXkx7/Q9lI3nZXo7080Jb64Y5tPvAPwTBQEDM/jYCWN4I/fvqOZG0F72d/6i
E1MQVdwS2j2pev6rvA7pOFy5VxeLGl0EqQB2Sj2e3qbyIgOUBQvIUgjPQcfaBrR1
p3dQBBlF8c8P4vYf4OOkTtfcabDYDq95n93S4ivj7+x0SDZEAM451xTGYNxrH4Gc
m5vH1520i8BRa/8VqQ6zdSCfFuMZ9CIZ+NoXIOJbSlPA5QKQ0tpR9HlJ3vJesqbe
V8uIKCLmvO0u0U+Y1Lu7tyqgaOjyUwVVGoNFSU2GW/XAN+EltaJ06toiluMJ2+FP
z5mRFjqh4S5Gs2I7P6dmdAp+j076GkAZQJRwe4olSeG3n3BqZMlGnoQ26CJXRTW0
ojg1hDVZmH1tjakUAPeLHQvyAOGF6THYqGxWgqZWRcILuK+5GLw4WCdzaXxozFKp
2lhmRzuVz1S93ab0R19tTheef5XKMy6FWCVWeAJc5BV4VMpnSYGb2Bn93FxH2CyM
JradUvnPofB6b+Cd8kXuY4FjZ6Wt85sjtEv/bZLgobWlWuhxRAnk6BuvFsDx2+uB
BNh5bsWlvftyvtAdA0ICbApn+usKM/V4KPOwiUl0euO9zTK5i/lGSEdREgeUSHxd
PcgBJ1ys1aC3SoGIYjc7A5zTEC38hKBZc3FVcwNXqxmBM7GGBz0iejsFb8YI51N+
0rzTCTc/XmBR0JPj1y7tBUFXbM+ljA3/f/XjDbcxKjJp/X/8QXSVlFZa2pb/B4YE
k3jfu3onAMa6LrIDYZRFFrgi8W6RK5fCOfN31d37+HN6GmfpPNPQkastzbxoFSl1
c9QiIts5ruSWzdMwXTVIoI2RMpwUNFiZyrxYmdLzQNaG+7jqeHE+Qu8HeYJfRLcN
oIXXCu6qnepyc7xmiMdJbOctKD6/+8bJaVGzrp5HjZNgniObUcgrLSnixu4KW+0o
/9nyoJVpz6R2l47Yx4/K1moJTz124XPYxYEWELqQMp3PfFThbPCwWk65cvfQnOQ+
ZZCkq8Cqghzo/1hnks6RgvIR5tGiA6qNDroux6FZ+Y9PUvrSZ/cG2vU0XliEX8uK
c/DI7bykZLEwz07KrblNZaDa3zspm1lhfcHIxZTaOc3dym/b6FIUkN8x26evtvw5
kLxq1hKG2zOXmt1TyXYCQrx9mzl9Ya0L2J4T3a/JdcDMja0djs7E1ChO/TCMdBCX
CyN4x+aQ+hwmwxHbgOy4c57RgvDUVjcw6uYUepQXkwr7kU2vQ4r+UPbu3ZMWSeUv
7xzYdS1Y8rIj54qdZ56KhPlNh/c3JdxULv659eoM1aBG64LU3FZeRcoB5cPrCd9U
7FRWtlDDY1n6sMo8Eeeo/78I4l65cybSIT5YkYsQNdp560F1E2EdmIPy1YfU9rl7
i4YvPzHhvVOlk3FaH7LUUYsl7oDKHIhPtWGpl786lyNfX3aagbXdVt72z9QZeCLM
iMvlM59sq5lJzUNi7xb41coAQZ4tzIdjRLaXm8gBHOupsQ8Vruu1fQU7pyLny76w
sz/bAObzCq/phSbVxLuzWLZBe67Yt4dY9kCY3My9OXuz7mP6TW6+IlAqtMwX3aXJ
TcDJI9BS1At3QcsXro1vx+tHF7+V5P7jwi8d4hUwVvUlzKCE1ZKBqjacOlDUvD4X
ERNpvpuZ/XsTzVUcszxqc5kWHl1qvMleG90r1BHXmaaN73RiWjuxyxe+a4mP+Tlo
RGHn6oBYLQYdyVzqur7Ho3fUC34ZxzHCDjf1ZT7VUH+7dRZ2StuiScyWIIK97OaS
SM3+8oJVJHO0BntSADCSKOpcLUaO8GlYNuL4xiE7kP1Zr1Z+1r/pWXv4x3ktyYNi
TJzmziO0xOknMYDUnA5rDU0K+JobDlDmJRXRkScTXvWI8Vxjlh7q+o8vp99PWBEY
bWrHa9OSyFi3V9sUitDsOm5N15BOyLqSiks7oz/6psF2o8C+40VRz4MnVLcShVha
EacLXJK3PL4gxShBF3XoF1dlCd6DUyPRGaV+6rcI5BS6D9DZ/rPw6AlrIDa1+T9W
s2ve9Dx84lIfsJ4fWMRnrIKyLdXqYGVi2Ulsm2pHDH8y6fgCHc9fkp0WSTtGjYid
ZG4bYsxmhvpBtUeDaspJ3CGqKUf2UY5S73vahbD5ddiwGIuiMy5OmeKU9R7t+X7K
OF2uwhzZXnwxWL7KrPwxkZxYA6FYzuqrwt/K9wa5TOK69oOMt+4mX/XpX8Ckovvb
i3cWSoYPx58eta307MgwdAzOkdeKRzYFCGSoN40fT5HOGqmUQvxJAIgWDsQ1SBOU
v5UYCLo9wvP2LBCzTPREkhGBz4jtZVftBrpBIqPSi1cAaEZF9FM13LQFi827H5We
B+DxFCO0zPhMek6T0+JNzOjHIG3zmM8gZMssS9ArELhEvjNLfyO1BGg5GnjFiAC9
jDJzpSpR2CpWkKRyfyeq2GgbY3NMSwQSUub/4vw9ygziQGKdkYPdih1ahTpb7FTi
Gu3BNKpV3Pro3DbpsO8L2Gl8usm0FKopkCycLgAbYqRZpGOtZOlRcNAMxRVydMY9
G2mMzesWWH+LOjILKiM5OXemA/PrcZ2Ioz4BSNzjcwwVQhwpOQfXYtJsIT3770XC
HY4vDn3AUTftGv3LEz0H8PnXgggqGtFp3b8enSEpz2ujeluKGM79DHGGS1dyH96U
iB4NdweE3RZoHpsjD6RiHMmcSiCa8nA4685CRh8ul0uWz12NywnkAltrVlUwhkHX
i6ZSgorA8PTSOyu2GwN2fVvCLk3+rZ2ZfJaP9IpjVHm0CUHczPsdYL+3k/TQRBan
jycZgTA1XhOrQMxDBDFp+/IMVra7hQomkIOD2COxzTUeGeLhGmSD9pa2IwLlE0w2
fDXTXcL7BIcobjSlBv+IbjhSaMUCcjNxqF0e5J4nIbL34ieAQLL3QQkEDL78tCgy
wao8McE3z/zHF/9ScMuQaE9k51jGNoNqdRKX+J2HNZndWdLL9d/8I/ywm95CWQIY
TqP9XUDY00PF66baCVap4A2rIBN2XFnnaUW1YHyc4DPpUl9geosPPRFoCX9tZ25b
NdEfHbG5mQAv4/Fg7GTnv5AQn/1IWx87ZNPho8MZBx+Ia02xOgqI7tu+JAFmDxy7
8q1ZKJoIrzT3a7wMPzPJU0wzQnX15LZ7T6QZLloZOfGky5XdfL3lfFa7jhLjFPAR
WyK32E16HEsXWvvYIRLdFB4URHRBMux1XOvhuMM1/iruGfWQMoqi/y9gh80Wzw0/
Oz5I4cPYo45Jfm73YALUtXBDTERSJEE/4j+yVFHLRrWrTVa6Pl9fM2WNmcOfdAar
rj74jSM0yNf3kCnFqLATnPxvKAFYubRmJEthJt4wFc5riaWbKkZmORYAIZEp1rGA
QGcqSggfWX7dBRRVG3kPhuZ6Oc9ywzdTXv9da3wot27RGB6s4pPC1MuUwCGHoCT/
XT/+f/Dl47TiGe/rbUQv3QS6I6lpuOSzQwTLDyeue6ZFnG9Sz1tMtCTAYziL+OLy
smU0fqiykaRMW9P8MO3KlW3e7L6liBkbI1R3/tXIYhagdt3WUIyV/hOi9yKSJPto
LjboFQ8o8rVJZQC8xWkCqE0aZYjBjF0kfDbbujUTczS7bs+6HMTZ2utegy+szIsk
dWJ0my7kpFHN0mtnZ2UASYi9QIJsxFV9Kz/quFWPGSYdRPCF0A4ENOceQaiYd2VJ
i/h8j9SHzM2TnoxuEl9nkhJul8+TqBdZ2A0LuViTVzL5y4Ar1EU5BEeadI9++QqR
x7PSXNfcoPDk8OLH/9/C7sslRpoGOSbjpQEun9rDoWS70g0z4TtkmPWA+fNwJnSD
CSK6nK7k945L7m2Kr3Zuq+98zgG91uDb8nupfs0Wxit0y3ZQbwFJvlcuR34Ewj6D
fs3srJTkKXYFmThwQ4yUWc6qs4/YOyStDuFGBghGN9B4Lz0jz7LmWGFgKoFba1e6
KCUV5abFS+aWxEqkaUfUjJZsOHko0ae8kj/FRPM3s2m2RFLmCsipsXP8pGFUhSe8
aMu0SPqpJ8fa0Qygc1vfFjT+FNQvHsNURhetF8ZUMdIvcULthtVyzFtsk7NjQkjB
wKxmdWFYkTXK9DzdlvoLunwcYY671N1SBlrGzmATYZB47MVZBN2Ii/LY9D8Tbcxp
28VFqxr3A0Cs4TjJPouPs7UKJ7GjpIWyJclOEsjfvgyZQtf/shPHfDw5F9MIVp3I
H4TLVr2cxJFKSny4F9llYFMRIOct1kpR+eM8qClEcXh9VoElPxDG/jd4luXP5uBE
zAnIU50H4I2vHyHPX3aLptNN32b8ZZ9HYdkQZVNUJB+GmcZESdJr6co1jc4asOMU
7BDI8mTzXif/WTypM+yu+G/L3cA7OlnUw8dJ3H2fuY0JnwrYbI4Fti8IdnkOrrbe
dyxierXewUr6i/BpKROseJu+OnZBIdkDBrt1gtyQm38ddR2CYb9GbeqIC1q0hp1S
9nEESkF/aoMHBMTwL2qw4mD6b8MGGZW1Y+XqYfy6CW7FQCn35OUF18U9cMzL9bmG
5UB1WPKHwtYgsYqQsQqXZODTtJGfxCN8jifBMmAhY5jAgDdJlxrHAoBtCV4zp5z7
86pH6c/13OBIS9zTBv7FHtEcl16TrOMSTGUj/nVXf/Bn21iKq/oEEAD9u/K869Mj
11KXsGfzhFaXsVuNo+P3gmte284qtTAos6BJsvamzcXqegtbSiY75LLbsMgUzTnN
SZhgm2eauCfRTJihdttmKS11Z48jZNjvGI8zzI3ql1NxZpdWmUk2BQ5oXDM368/r
uaTtBnNk2Sg/tcvpr5KZKfAQ7uAZxLDsDtCEA7XrEJGtb9qtMiV0zdWC1H2x/XQ6
Q0h6Z7zOLxiGxSAeVZVm5IEB6x65jjLOeBphppvDXO2SzejPdDiXc58thmYDdPur
ExRQKeq1riVlo9CWDA2QWiQj93Ae58fyjbd633diNJwVZkGR15xdVS5gWlKMRf9V
xaWgs6Oh9iFhPunKGzpOOLNx9MsPmm+hUypE93bh3HMVJJjqYtF08pPI0HRszrOM
VSxCM/k8Tl+0yVmjC6gb8M21N+vPanA5t+TOaz1d4AFeQQjAR7SwUuALO3rMfK9W
v634mMKl4tI6XjmnQXe4RE8lI1PrEFdtQcJxkuBm5ah6V5kztEAFJXV9Bf6eHURb
tstk1R4ORERdyqGVhtFQzXFyuR9svtwfIboDayygm0IKkJqlJlW5mPML3XPJDJHu
oh8EUTsdSgi1BU6XQeDdYex3LLmliMt7qS3k8v5aaP/j3w+QmEzxu2UiqwAvxTLh
DBfincSdSP0Z5SmBSKfbdu0GIf9ELaa4g+6KOnS/lPkc2Hhgl5KGFdDCZzCst9St
H3MszSs+ccAi993FaEwn8G14LlyQamuaHZPmx4ZqyPmcsEI5Xtb/HeUdan2DR50g
9hg+e9Vm0M4G6ZgU0si1ukBctt358p7/OQ1HdMxFLda5O2mjZVm5iTYklHeyLWW6
uZ4uN8wb2GPWoPrduXB5Nc6uV9d1P5L4yZvycUlYuzx7DDF8skGte1nCDATqHv3g
dquU5O1wXGKpiuml7h327r8YmDtIEA2NlO1frbyTBrDIVSA4MSytj7PHk/maL/O0
aB9ivlKcM7/2DhXNM/r2Lql7ZllsUxTyD15pknxzpkIccNgAaTz/Pnif7MXBCCW1
mXhnCxhjcmOzV5QwVo7Qn5f7+R44goNqWRQtWkGHJcZX0zMBdkVMAabyl5Jgh2bc
aUvrmnGAZn6ymcn7sWEAjDtX1vmKn3FrTnVjh1r1szUdmFijEPEvB13mlvbAbgQ8
UQnCBI5ij40EBVBoJcncbOVeCpNB+sFlmRo+RsfbRxm0D3/OabR6p2O2gp6i9H5T
qyjIoe54pm/SHTZk/lZ4iUnhqCbSl8x69iof+oNlgdL71RheSNXJ1hH1bfCt31RU
oEwkAadEv9yB7kfQ/gQ1nG0+F8YSrCKP8UcHFsjDXywtaFD64w8kdGncjfNwYZnj
wjkDd01mJB1yos0TNzItT/s+BpJkD/AfezpTIY0A1D2GBoIm4PNpCpnGTP2UffJF
t5wJmdxjfFhBQBelE/6uWjDBY2WPao4BhjZSwIdIB26dO5ecX+pwfrNGoS0YVrLc
j4Vl0drRmeAUd79edzB/95jgOlbO70bTcDHNEj+Ea6uoKII0GB+5OZFJabEiSDlj
2NlmkSoxh1JkliKyIgFjSyYlHXWjXR8tJo2c7cRrrKMuotT7OVAf03OxQRpch5sf
+c4pfSyZRpL1BaFKyd3SdtAEP/Pd26nTf4/B3WTsG4mIM4+v2bS/QSiGNerYXgSL
Stylia54jUSBJjWU6R8aH3/lCInW1e2mJCzWXsmHOeJVSDJ9ppeXkUtsUwzPG0yP
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgXReg.vhd
`protect end_protected