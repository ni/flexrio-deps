`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlCMmAdbgklDIucpcNMr0PlKjj5whe86NDV1akweuzlZs
xF/INWXqONPgaUHlHdQyGhHp57HCXr9a2xrGaLJf94NkVTA+j0liOo+87xhQrIyG
XGS6XsohIDAcssPONbTn6E8y5nNNZ7/SFt9g1EkH7Dgg/I8KmcofQH7GbiS8mg6a
+JMd9vwHIFqYoZ5qD8ZbS8dUM0SMtqplv5VP6oWApGwWP8VYQPLEPkWnVjUoj2o0
4FpnZFiyQihNNxT5rUT/rgxgZMbZ7+opJRmflZxmihgZDB8FwmgN+ykf432oGWxD
1BPlhL2OkgQ9l23oMTmq9Aah0PCKcaZV/9uB4haQkGohkqg3Qi/+7ynKWMhLZPU1
YnXT0QKpkmkN4BQl6HUXyATUI0zoCcIfh0nooIAndMPtR8zSkOu0P7+jCla5rIAF
0u2Yk1QV2ZKb0X84vedMeekSv6f7PHhu3XQWm8ONf0jF3DEYMdn9xT+a0d9IYK0W
wHk1WccoX1ypR/RL3ETUDpV8X6kVKb903rqDanBBe8wPWZ2dBtD90kW3CzXJMOSl
QXk449+rHWTKNOd0flx8iJvqazpY3pcLDPDnI/UkdDANPNYiDLAFE0pP7vVOsydv
JB7S3ZwoFcDCKW98Vh23bwgFJ98kpQNIfE0KDL9DhfTJgl244JTlBKozYOfGxzSj
C+oRKYF6qbF22h8dkVMbfRX8pngnb5FlvYLI0HFROWKQJXNHusrvjBep/E5tG6Zd
Jr02m/4qRaEx4/gkDoa5qBnFB2087ZPwrITmY95pGfDwz4KZU3hLXjwTQbYjd7nw
NAFMba4AgXpK421wQZbH2IXYoiTsEb2nIWYdSeOIrUYLHfSby4Pag2t3nyw0Q2Vg
ssB/o2mJTRgBhms1WpMMTImVuzGBm9L5rr+NuVFK4CFFzXsmmsE98J49prZryZfV
ERCrqvIFecuquGHxQfgAKsb71unj3yysSwH3/khPntBbUWw3jTjtHWlhJwcd5Y7l
NGrSfiZ2LELMSPWOVo+iXL26Q2paKDa47zYZ6gtY9HDPydQY24dNRU2ntuM0QqLL
lIYiOUFf804dGoWg3skFcNb7X0q2hUZIaMp3qp+/rM26fxWU7z3jf2tkR3ob5OUM
3ijKIv9tRjL1HJwVdAPH/pg0BH7AXxZbF/eGBvMpeF4dKNR6JIOwc8k6kjpJyvOi
Hek/OoIXQLdvH5QnWdigyV6m8+dOVMKvMRd4b1UVEIdsXPX2vr+Ttb8RV47aCt/g
5xN34HSPHB5ymWlcZbqCv98Ss8v5X4Ybyix28imKyZzph8ulC/h0G9jk1syeW4Tu
NQaIGg3CtYMLa7pB1RPe07qECgHRXdouh5hQTJLQOzSwOY/Pr73gekIRDJcIGRMO
SOMYxg/oir8lu00S4ft2u78gWU1Btp6+IzVACgGbRr1S27cjFGhcyhdZbtNLf09K
uhq4W/r8dnPxRFgMKeHKOjH9GVcYwmGAx+oVlzYqgGaYqMePR9mK2KYXJT1T4Q+Q
9X6HwWPrCqZ4YyGSJCVcWFclibsWp6ZTpd8tnNCaiBvSZJcSI91F7U45CHOC27Uf
ANigKkk3XKvgknQ/j+0g8l7Nu8gOiDu9SpITTQw8cVS7RiqoJwcqmVfx/a5KPa+b
7ZtCu9lACW5mjFrHQ76SdZSwzfNpXH2U8gi2QcqGmnloEq98tc0W1CnXmbsdvtcO
OZuld5Q5PDcZeBrnQTaRT82l/+I5jRN5NfrI1vNMwB65bvL4vXuSuIPLd1wrXcU9
SIrxsWOw8O6a5RbkkB2vn5Mf3bsmt25NW/jHWI+Ej98oO6GieInckdsiHegfXBPX
ZE9UUdzKeOr/lrwwg9AI4s1NNdpbORNNsq4rFuHzTL20hblyHmchJDC1IfxlBtGA
NZSmtKgK/ZAUf7hqt8hf7s8wplSlXXbCTb4hUz/f7d7y61OAkv1uroVI0vy4Mw2r
QnsDue4jEzZ7Bzx81SceC3r29lfjx6HZ+NLTDeMurpV98Qvbd968XMstQzF10dtk
mQBUGBd2g/GoVBvStsq2o+FROa8fjBhM9ywy6Fqs3XcvAygQ4j7Cfimgrgks3CzB
TT2xkppuTMv1b0Zcn82uVxi4w44cS3+A/YY5LUISuzw98jjlTs1vDV1z7t6osOfI
VSnlQxn03n3Kv9/AUQpR4dkVb27Pd48h2KCg3A4LI44fGuoDX3gVbrLH56LuviuJ
sAE3FZUF6wZtNEU5ifWhTrXWvGqv5qBT2nOpwU3Xli/qxMJZVnNGT+oYzMHUk0dV
j6v5aVBYD+Gpvt/U6ivfY2WjsABb5bAUMSyjUcOYXaKq/Kbaf3Sg+/Kxq9hSpIpb
nt/52Q/LdrYxSDr3zviMlfdIglgf/VK6HIsPrJ2eKC1SZoxchzajITfd2MoyUM3e
sbFGYLg29CGU8ERR8Pru7QtCtkrUTZAHGw/nzan/FHvPJ8ZLkqnh4uKU01DTLajv
JECoQQVILSZZihHhm+FpfxOp+w++Zky/ROJ+1RxvgU0hR60vy+AjgPd1vO1YtArV
lTJ/KZY4NNA6PMAiwQheV8D0ZKggW4RnSC+jWtFXcw3ylX2Op7pwbtvhIJY//VLl
VG1PbNzHN4qM8s//kDHkPZJwj5ZolLM8PyLzHH9RFQds9Gvuphv3bb0egQzEGO8H
e5WZaxjwlH/NHDQ1PXMUcXrYKto5T9tJKeQKzOYv0Pb9pciSmYd6MyghXk9mmHHo
XR3V3wnCXZj/bi+p2tsveBq2zRQrH5N7NhX7+AXHDZbJ62sB0nXiMrX+/mhhXps2
8Vhkgegr1ZCK8sZDy1eFnHqNZafpYL+Ldmeo6ohUk1tKbDWKQz3iUOFKisVAQy1r
P1KFh26l5PWkG65+vzIYmF+rzC5jo2hiY20LVKwl9nZnq0xEc+jRvwoBNHcLKwDD
LaRBGuQk+qVgF12/ByvRPhJDBOWYmlnBZ73EIovk38fnhj+p1wghvVLC6lgHpwg+
WqarLhMDICP9ycYwCEBppWjz4Vj6nndcB4casCn4Fj4VtoG5AS7dLDiSlMqoZtgP
sHxqzitgYjJmYOConq5U09YM4UG4SimmDmBE4ONYZ6R2X0mWTmhngJHX91tawgWd
Jqll5B9mdoIDzbJhuh7bVTI4GtC6hHa90H3dekDlmuxzJ9RBNoiP1m0YS2WEdMtL
evDCrk7VplE5SSRM1q+ZGJSjGipv056lKvxQgg7eyoErvdBextuUYLOfjI5i9SFz
ITMAh6fw09yNT54Up3D9JYUzxKbbE0gAg+lzf07GYZ4wqg40A4ChGIo4QDu/Rp2o
iLKqJwPrBaSXzkpi7MvgNHn/whH2Pc6vyVilnDF0ruYZXLNpmfNGpyu436g4ReTU
Km5pBDToR+ZZ/Y88cfLDf7TodIAPFfnNmdeWoqsdRw5+CQW5iJOJ2DbDcpiDMnyg
39bniyih+KIGnFXVCFuZxbDTgNvIKWq0mlT54e4UyOgmURpkwV2nSc0Tj+GLOLgw
Bkf5s2NaAMYdCghYeyisV3kThM+wKY51DfnZw2rWInR0+DPt2kLYX8t0Ul0wWHxD
gQR0vaWd5dv2lOLkbCFXxNuKYTjgb1JnSP1dewoFtjzvgLr/iQ5vWy2h9QiAMGNb
sZJ+nDV/LjWyV/+gHUR77GvF97rsuTm4hcOrGHVSiZaw7rNV1jGlujjqvNZmyEE7
UZz7wYdUlq2t1i5GevFtR7SP5D9mDVBwL/JduufexJD3EF1fIDyeQrrnczIg86Q9
447t9FL2j8jMKnFtlNJhkOxllj7tqysDBEGxb1Qk25hSBdscsHSuw46IAtvYtsqv
x0PYeNjsdMW7JyzaoM0aqmDM46tmCxa4ntkU+NNFbjZCOPOgVg0G+ETJIaeh7W0t
1A3ZBQOVq6VdH9nHw6+SunusuzzD1jMvYa2hqBNoTBeIfeOxB7+T6yGEgtKVou5r
taVIUltpZCGyjN2TNAYmbYCa3ouznJn29McxqrQ5qoHLThs/GPYAD0PQmDaMu4kA
70MFITR4/h8JRhpNY36eG9EGtAIZQx7FZTccYwVBsGsJZ+AKyhGwxnE5t1rgu+kq
vnlGeOT+4Mg4UiK2J+wypM9AnPAvuasJiHzm/GdDdlLgjb8srcdZB37qEf98X11A
2BMnWLxI9J7H0ncb6SCAwcQDAxvYk7TeheH2dqi9inCIlapDyEl3+Im4Vpxjmrbn
mf2xcmki7dCwpjt+b9NFRNEqUV0t+tNP9WCdPZBIilVJcB8q29ok4wCj47NJ5uxs
rFalN8WcPhH+ydr1TrnBX10UGU6QaRih1OF2RfIh8GrxdX1TPNICwedZ3pHWqN2+
L23g0pLsdH8udOM4/ahjhAFatZpk8OIbrLF0sMSypEG5d8qXs4VeNnN5I+AXfPis
jqyX+84X3ph3KmdBF+qtb59d27g2atel/Gx5GD9kDHJfUnHOw+y2mRbxfv4a689e
CELe6V4XE/yZaSesXdbHQt9AyTdq0uYX10BZbHEC11kJ+h8XiEiUFT0VNMfhNZCX
UTQmrbR/sxNp1AvXdCdnf0QgeXNfsWdIlkeLyxGXfnHVVMuvIcyzK/O/f4xG3Iyz
wP4DDOlcUeDL0ZfvE0+6Ku6Aw6GMJZp/sahdTJsvhbpHo8MwBlTCtpcN5tUyQahO
1W/7FANURsvcw4bD9TM4vWD0k69Dr5xmeUHHhHfLw5XSkHX8HYBdQxHoAopuAs9u
rFT8T1zfDWYCGg04RCPlxAeujqMLIMETVGQpp7IcGMDg4vhfGziQD7pELwD8GF/u
OmGN9FoB+p1TmzF04NpzsyQdf/BbmK/Pve/kGeUJ2y0u9jyGuAkRnGmHLiMDrFZ1
L58JxbpIbSnzqnAq5gKCwg0+mQa8Gvsopd3jApqifCfOUxp0ZVN2lDBXhqZT9JVy
kO+5fm3aVbLJ7LI6g1+UJmA0AmTmic2zuyOEopGkfg8AA7p8C80CMlPbA1i707Or
QURUtrDoLDWVUuxHwzYYlEkgQBNt0IpGum177OZp8tm5DnahRuFLHzDHDCO3SJmQ
6R7aEZXd+C1pz/DnpK/GG83jgFR72XPeyx0LPEVpG8yLM2KpuMn3hb+Tzv9uXiNY
cHDmah0ITOmct1C/M/jcVb9bc/i+USzvlmy+GH6cTCZhkMKQwjSges5A23KVYKD7
fCm4IdeQ5X+zBo+pIPTglZptixKWa/FMOVVwHz5V+QAosYuFPksgNRHQOqOqGbQc
caH5Gn95fIkbsPIni2W+n489Qvw6yZL+kh9mF+0J4+z1akn1iQ5Sq/lVowsb3rDy
3KBIldrKQbmF9PzVhWRxLMZp6igLi0qUY11JRaW9jEfbfg0fqM9KFsbir0tdZs3Y
zwzeKL1lFkQ3GrgoRN4hlllyO9WgC6f8/onNYuWerqWU60NcrhtJJtB+FW99p0T/
iMMEh13oVrmN1o2k5WmrAzqveXjQldNtCuPbD7CTRkuH/uiDWlC4d2qmyzxB49IG
5YSrhnT9wZ75bHYGfC08DDifsnetPOuI/0vHTRIb7F3JljZWz2PoEd0JN9L/2kjO
mWwGwiB/iWU7OkCosy5P6LuKJFK9hE1x8siMgic4gav29E59MX+NjBZem2ZNB7KK
we/7Dk8S0m6u2AluziqAjIZ1OskMNv+ScaTKLmSlvt8R+B1DX4nvy3TR5ea/2GFL
331c4aWzwLxH2m6oLiPI2Hhm3Lev8sFlgEE5hglc4Bl5y/Y/vauVi9M3qaXBQBqi
FbPeg0ips/P0dxbnH5CEps/LDhk6KjD8ipATCn7hZQEzq0oK4gg4wXe1qZFfmgDM
mwSi4labXqEgJFEPZEfUzMCtLZ7ohhYeru4mPzYz9D4i18q0PJDxtUhy7RAh1etX
QU8SQa2ivOwcI6Lrwp1eFS6xluPGfmJdGSmHCNu3SDsLoiz9zbTrnfqJ1IFjKamc
3mu9tn3PUb5pPJj//+rMARXmhFEfLHU2UKdVb1GHML6Z9d27zC2HIlMl9vuRIdQp
2ilRqXwIfGwrb4WAWzfbB/nsex8GMUatoHhdaL7k14+EbNtkcG9TxM8pEEgVpDXG
nJydvqeWFgjKT19zp1hIq6K+DNFHqmzR+XaHkekbXMbWJ+fQO8q0Mn8pncViSnX8
OfBR/d8GwRmGGCy3DhmpCZfat0peEJlI0J2j198AmOXMOp30eDzZ6ZXrzcNdcpSe
o8qvH3JtFwZOkpOvQ17EdC2fFXzdcqSsiEQA6metHyN7hL5PLB9T/TCyE7l6JGl+
EFVBA5B3d7Y2yXriikVvL8lsU0r/a4Dk6LwBDM1VPbd7uAVSjLpmgFLOhvs+IemA
oXBlOGZeM6uezEzCFE61oriZBgwOo8hMi/zDA1iNO3tLEHQgFp07vvOx+bbVql2v
atpbiORoBz3XwrENivSxqXFtCrpTLrfNkl8cJGmzayw7lpIpvsctV+/BZgyTaaEv
PFe4xToDu9eoLkwY4HbOcXtr/vSVb3CAt35qsP8NTOaThPFLgT+3ZyCfyjWtgqSD
N01RrHkWHVN033gpv5Rq0VHBK6XqLHUW42sKSbCGGZSsSdRq5F4QVF7S5k42Sw0S
Ds1zWC7FbyoHa93hEzIiuFXmCkVgSTk0E+LIJoPVtejUcdCLR6HxUDv+A3eVkDu+
8xaKm2XaTbW92Vylr4ggKPKD0/ZUTkUrXbjThEm6QFVSpj/rlXke34x/BlKjABHc
29ZX2F2KhVeTrWK63V/0rgp4lGJVtJoe+I1rpO8Ux9Wc98b0yo4XSd2mpqZ0GV3Z
G1y150xXdtBRsvLBud3/m+3zD+5lpg11bm1uf17bhy1PCWrAEfEnM7RvgyHrvsC8
VDgO7bswgpIWx4FbG8Xk0mgXthpehvlxhT971vi6Ijqy2/S8u37lMIx3vVU1CXiG
kcn00JFmTK+7sE60rMMEpBBS+7Pb8uBRkyPHeRFfWtBW0+mEzaZYKMzkmxhltfOW
ghUAPWooUY1Rc/p9se0lW+4SrQ/nmPdYbvXFkB278tQpMOfC9b+bzyuUxQJ7wVqV
aRGBkNhjzyChKW2x13wZNob0ElSJ2R99nZTw8MZvBGeJ7aupn2OZkppBEraLfI5H
+jxwWILP6UH4wOSLXgV341jiJihkf0OEN06DIc1HsB3QOyk3NpM2MEd3yGvnZK31
tHrcyKCDkabRIwUjfcHj2xM6Q6qPwNX5+6GkJnR5rLfcxKTQAWsxBZcrmwgIBWl9
kHS4vrd08H9pd+9QEcbfpPHqP7H8ZBLSq44Iz3h55TubAbPTAh9T0OMS4+4xZ1UJ
LLwwOPEbVFb/0kHUUfsr339i3reoRtgu+bPn7t36PcqBWihqfoDNTQXLj8UQU41T
fzMHkqxmmg7wG8wYbxYsKdQnIemGA7YlRLyNZcEVUUtEd0BH95ai9hX9CWF4HovH
bbn1d1DFUEJQQnXIEkqKPWU91yqS0m+AC/X3pTImF6tZtXnXVvKoLn2fQlKg7M7q
AfdKq1AnDfx5ufiucvYTgW8p+qrzUNmxcIqS7yhH8K6w00eFOlXfUyvqKGVCcztr
PL1F6d2rpluuVdUD8kQhtZfCNZVneI2ckdWJB/O9tj5lo6KmKJtv9SJxKOifSIWG
wvVb3w1ytrVeVAmKadlwnegctG4Ef9XBh2YB/W1/6C8ghXG5Gtex9WiWg8MG0hnJ
/0dstfKbMbbAIB1hAclfoq7k3nDljELhuaJLkXsLJxt/LVwpF9LcX+CoJOX1BEEZ
QDpRr2u4v5JmUh8IyWCZzzhx4Ho6LB1j3weIFOqAD0PT+qfcXpWoEUxxP+Rgj611
1HYp07DQhGY6ar73J0tYdVzULJgAcdCmGaloMAgo9Ec9kqEG+sGoBaZyHh2If0ne
TJvuD1K5Ax4wM7fUVnkw3STvUcSdRe1KY5F1h6Pmv40Os9eALRdhED2tU1TwrZgh
RQ9WFqYSt7GI+BLCqkVX8eWyr8JKhZG0d5l9mLdA7CkDXYybU1wAlbeyHlfLqlhw
snv3UV3nepQJKVzdn9kfgkPCXF95+3yBuFYHdrqRbq+7yu1DSuNS7Gutjl9OhEjT
zUa4aDgu2J+QkgGx9lF3vAwr0+wRS2G82JS/xcYRBdiNrGx1etFB1xDNTmsU7HVx
HPoBwua87mcFq2w7ovvRikv1h3pPvARNVUYnlUVu0WdRO2UiRIjSJRa0OghSxci0
6wRgmXH5ZqbP9TkD7Vdkjs6RMtqxqTGF9L65NNRhwme+RUrH0TomWuCXI5fguV8h
T0+qx1YJYjslgCCKRtkEmYdqoOtjSJfHrj2ets//0WEAHRYHitHOFNHdgv8j85QI
VHKYodM7jeCQU6oqahP/CdOudfanuK3EbDtHfUrJ4rT3ppIR+hH6qxyXzYvxV+sf
gpJ7CiT+9XZEZAI9mvHHR/GFg3azlugON5F/c7SoiurjZkdD5vYvZEToES0Es80S
5WeTps/JmYEyQJwRPSSDP0mUnjyliu06yhhQcTb+j6Cz1tcA3smhtK40ARBiW9U5
owj7Q0TulhGKQGxwrDEUtAsL6NZf7wmkdomJu1wkuuLQtLrHmeIqCr3D4xV02X6X
LQBBDOUUnHHDQsUAwbZftR4tBiJ/EUO7OYmYYjrwOaKtW2lifE8rUL0izV4ig8ZN
vkRzmlvrBU/xOYpqirCsaVDkcRiDk3/Ng9DdIxoXDeb8aSaQR89zNrMfwiptTGTD
NVrT8214UqDNgdrkmpZ4QWgPAUDnBLI4JkUAQdYqZyY8F0RUZudl46hSMYSJcShR
A0CUBYO/YFmBIbJ0Z5+QAJXGey770sisQWOjG+SFFir5tuQzQ+dhnYhmqDS3rXTE
zNAuwm6ksUQ8GqH/OksY3Gt1RyPV64AbvF/mseLiJB7GazSptc0SuuzGvLJAaky4
aEKoDZWo/df/g4lo4MhmYGOoMmDpne6H8k7JNNrI/vrmVfSIhxzE4xkfgvgSmtyB
4/FkOaP/SclFGXOYBgVao4unRnDDKPYhIW4iup5T9d+6aqTbB2/nm0Id6AUxCMWI
IAyma2lXCwA5V0rutFmu8rR1IxxdxNvOeYAlifec6oxdJJfaOTVR85A10UaB1ofi
tpv8lG+KGWmJjbWLf1/TfzEI00RIrYrUKhaeunuLEqrsUt7wWTSiQPKpcuvcq/sg
H45E7JeRnOzunNLmNWsHhEopEDdbt9ryuFxyWdmU4uReT/pjwlhdRZqW9lQfcWk4
V5df5CUDm/uEALJv3fc+VhksYmkFPcDy0jiyGqukzIsdvr5bjKJ41eywgNOZdmGl
xl5WY3J1J3AxzasnbItRqR6mMUiS8TyRJBpO5yv9dGW12zApDNdukG0JBDpVfOQ2
+ZCgZ6ZjdG+sNxT8XURKnOUxS4mYETKky6Z21Jk+0Akz4+TjlkuFvwOdHLsrzEUq
5B9aw8dkBUtwq+W1Uc3Nkb31Im13+TUJzVY/Vv/2WqZM2TmXipLMu1oojzc7jAYU
lWWTL+PKwtv4Nc4l9JVmRjY463mlZxX3cn0WPzNT23328uOw+BrhDbL8FsGExDWV
X9fToKr90JexIHHQRAKvccm6yZSi+do0uyBR1SBDA1iMTaG5CYiMLVecrfYbMCX4
BfrnM6sRZ6dNdTBf1EyEkfJoTN1EiTpwvTEGZOitN+ngZagZBSxFtBPCNg4/ANTA
yucDHbe15a7mfM6OacLlB89HkY4vVxfcSQxoQP0pEDAv112wSrcUEDZ8HtF5EDr5
L25dDwsi+WcxJduk3uTT8VmfZbK0KqZh0LzL9gkUevY9uqtpqlFmYyM17bRtdLCP
i4o14K1voN8A7hIg08LpIijUcxZm520IZ4Bbw/I4IJ8td1zcqvFOkjjSyoAW9lHw
fpviSz+XRhO4F/LoWeoYTJhxDXNEDVafpfJ06Y+37JbMMjNZ7SXPqd2d7PEhYoW4
Yg+kOX3WvcM9yAIZZLrfIvExBhShBrOQJkrOxHBeMlwMiuqI77TIWEtLBbvNNnUw
mgnBgbAXijehb4bEHUZiqgMhtCwOUK+tngoYx/Wcx1dx9jhBJJPeZqHuBGx1+Ozh
IvCJiWC22kMlHJT/2dnyNoJ9a6okcfBllxlBRl5YzsA/Imx0gvn/PO8dZnF/fqTq
6Hh88n+x7kflLtPw1T7bNpfUiU5d4tUbEVxpBZmli7CO8ShBcd519VGHbIAgZ75P
3PldVa+X/nNfxZo33hyk8sAipOfHrjFS+WqyGErRvC7QN1FNU9rJYfD/HO6k8q7j
tcVPP2NU8SHlT18MbOXydCM27pAr7NTbGbaGipg2Vl0f3nR5VQoxKzVns3f5Zdaq
fcFKFKRpHgTTg8K0FKTgTZLY3DNjVjY8lTUJNuuMaR9MeuHNbAUkMOr+uc+LDyPn
wXdQWTnL/L+x5iLJeawZ/1zAhMQ4GzGZ2yD+0IL3s7EY+Kqx7yx40e1g3/BZ2WpB
Uub5NUueA8w00MTEG0pLRXIVO2QLFI4OUyyYpYhBkVzRKPrCFXmn00F+4HVNYdG8
7xCpa3j7JggwzH9MLIgOgDK9TQ6kZezvpKEUHenU0Md79KL5aQvNZvuSynm8C/85
sU3j4V6YWO9xo+l318ZZbMqb2gIBWVnTVOldu5h0e7RYje449FN1aXLYTmSsF/xR
G1iepXyoWSR//y7N9rbFukilDT5sFmtoKVmhuRF+MRuWhjONDMDNeiMahQzu8fqC
7T6yLgKQOXHboKBs/hYr4bBYx8wEXbPHBNqIXLWKkkh2HJFMVclKK0PJZbBBKhbH
nwz3AqvjdwDEtDEiGLhV0qpOS9nuLiGnQPihlnxLzoIzNEU0bsdoy/9FLaTfBQ0M
psZISZ6lLurX1CYYGSyCxAa/LwYAtuj3FTyb9+5xAV397ohO12RA/W9pwN2r4xZM
Clkynrv0mJnikSs/7pi19+3pCBvms5NZTLBjcIr20JqmzvbpZqPtR3ccTZD05tV2
7uPGTf9gc+iqdpGy+9gP6lvHi/cNnyghImGyQbHFUSoK+5pzqwe5qhTjojRUw4kU
FnROWPlWC4NxQiEXBxvmRWIDyrPJvX6SaqtJVHoeScSajBK0qID4nlL489rkb00D
WzPJ2jF9UI4+0psSUJzrPleM5OEm42Y2cBjyuvX/6SdtklgYRQn/RrXk8AslrbyN
6mPUsMWxz5+y31I6T94MME1vXWk9LO1forpXRp26ZYbbq0kqnfoTrCfEqLvx8/3d
7CK2c80QTuhhVcEIKkFaB/NCNUhzjxQVPzoN6DLXIlTVB8nG+SeFmSaN/4E2ZTid
123oNcSysJTbpxUsyLl1e40edStln7MRi+FYi1gA+XEGUIRF1QVv1OdKFc7ZnaTn
hLZ3b5i5adxZdICuMMj+wCgDq90Fh/TWfhmdICFEYSAiU6TfGOwA4DGYFHfFTkZq
Tpw+R/P4cC7CwWp0ntlVa8c7idBOflt5gO64rsmbwAh0q0tIkCKcWkHIEGt5IGfM
jZnxWimuNwWiDqPkrdxfwrhcReEmFKhJO40Ya/Qw43tw12HtX7ErcfVO03lT1f3q
XJs8iw2hNals5Pff8SHaMe+f4/fYXD5yJ6Cb7IFdv3I+4na0EuWq1ZhJzmPOjvek
bdwCwqIWOmSM+PrfmewJlyKskaA9V/SxJ3rH5brxqBf9OlewlQK1yXkXpah03WM9
1HkX/VVzS2z32S9zFjf9DeGTkvdEhx+Ck4r6ooUTDbmJwFhPDWbi+/pbk9b0itIY
6HrxrKC022u0cv19yx0s71a6/YpArUifsT7fa8G7hAje5VrQHUYB/i9eHFc46sxl
Ce7RbNBdAH3Untd2o+nkKcffKcXN7s6RTN52Dw4JR8LnQz9k1NvFJcZs2a7RNuRD
uUyWNZggQ/F8S+ddQAyNoPzuLZE5moTRJw6vmQ4anJRs455RDMaHJbovQ1NCphDv
q65BXLlWf/yeg95ObbBZXleBLeUzBcElwzdYzs4d7zuTBgbtdkA8Kxej27DzqL5e
2Wi25VbXGPDIFvIfTPutBBKgYdqaqDbVzh+/NKWosf60K8zwDpg3Z1O+h5Kg1NXK
nVj/a4MWWy7CNqDLix3vUjxHfZgvnVnXGjb6gUCjJmrPJwb+rnMe5AKYYl3D9Jo/
M+otZduwe/a/qMYorhyo8auoDWJnDbH+dF5uQeLS+6qtoEZQIFHu13WbuhZq/09x
U0YdiiZRpbGVTfjMCfwVxLmpO0xjs0KspxvZ+a+9rVze9kzWuBvUUG4q73EL7X06
ZZV7loVTWTGX8PbCLaDlQYlseTi67sZuXqK4yoE8j7uy+AshQf3eU/0LZ4eUJKuI
trnoE84A4UesxO8xvieZ11LxTCRhXQV+mWu5ui2/QjFBpki9vBw1JT4LD7QiEYz8
eyZU/Y95jRgTRRjopKx+nLZQz90ckgd00rKbPifvExgkx9ds7Mb5gkdfhvYvxiH6
53sRqEQCtLKUqSuY43SfcoBOq3P2UQLUJS5BknK1gPPHzZ5lRMWGZmRn6/4ru1jx
a1NHboWjmMz8vIcVcusLICMW02iCL1nbpW92PKl7JsIogsUJC+DwUKkyhmFUBrY2
wElHJUtI26WHALaZEsitdfD+b25QJw9cdOfsJ6F/VdewfS6A36bEm4oOO/X36FA0
rxXvPFH+NsU+af7yJBgBFnKnBatfDiJpqiWR+iJOzujcc4y67Pzda4L3pzRDLlDQ
fztK33qYgZYnx9rKAFulKSYansStwDY0bmkjU4A4hH4dW7WL3YAHsyDJQEdfwFox
C/wQUhQIpkZhypy45VEiSINyNzOTQpHFUelVMO8S/uYv9m9IBFjq7qhCgyXa51K3
1EDgzURiIbiGecnRTcn8W2idhoXEsKOob2DWRQ19beVuq0mWmUmOByuLsnHHaZIm
w1lW3J5BlJBWPcVZhVOYmJNsgLWRr8beZe0QrPIKVz+6S/4FsdoVhdqFegmc9oJ/
GLISipD4Ejh0MDFVxu406GghhkZcQXQME4B0OYbG9xaOEGnQ1M3JXXkZCmfAo3nX
ZSQ60ahjmTQlEyB3Rje3e8DccNp0ceXzaq1qa5n3B/asn1u/7RjmgzA17D5a4VIj
z8CqWsEXGCQz0kFSbhERUr988jyvGBIJCs0WxNcDoZTaqQVcx77f4Gd7lzNtIjxk
xIpj1VRQjl3UDE0sqLpkQzWLbS27zZLevfasQZEh2z4VyiboxpN6mnPpx9q1hxxE
oxmvX94AkT2r1z6BKJ8qx2CDVI7yduh9Z8a8dFMOnm9QJWYlIZEuQThzueoIMeIq
/yEIbYZEo5KeyfJULJW4Nn+4y+j8WLo/ZPZtjnjNVHd4E+47ecgunhXkie9uPNef
2nXO6ALdlXuj5QILFnK7LgzYUoxx7BI0L+G4goA9XrDKdEuumvmZk+5LogvNcVtL
eWnvcIxHpAluVaG0bAZ2NcOJqbp+ogl1pUEcc32sE+Ugj3IWVNHDpmM4rKnrrbgm
IWBSvH2mwK/FTFDLvIYopgrjjvEBc2pLTGxqQ5mk0Idy00jUnJp3NCDcGvIeVYvc
F5Hn4Y0KTsLuavhp5F894UcqTKTL0n7ALWrb9r3DAJXB2xisC4VHBjoJ+H4Pr1SD
OARvUgGK/Wl7qDu2x9xZTVyRBZHv4Bw2HDeRm0mL4PwMiblRoh8ADmIJWY6/xrx6
3oJ6IFQWTMCyR5IDedM1jQmMZ+zDF04zCWSY2P3noE9HamCibfvSiheMJ3fh5YeU
N+klYlbQxs2NNWr/xAeQ173AqRoDWVm7XRFo4MtQb+RdR+PmiV1CXxfB438sHRke
pe0EFZx2sIcHAidudcqYX85YXIz0VJb3S+xFrNAiSvrMZF5NZg2QMklvmmSMJvrO
QUIRADRVsG6KFE3AmD2DU12i+nwzg/WqntLJHSINZ0rT+7u7vTHSgyCgDmKG2hrv
aymEg5ibcSNXvcrVPK7lLpVGJE3IPgg9Xr6+1Ar6BxQmzT/8o69RNapfjWBu8JzC
m9xpTpa+AdHGFjtQhGizV0c8YWg+JMPP471Q7yxo2UooMeofY68L0MkZ5Mm3sGUl
M3ncBNtIEIqRyot7xSIujJ40gBFCg7VsibtQE2AKMXD/l0hXF/RGilSEz5O6TkUJ
cvw5hVCNvKbsuou7lWL9zFO3f8hkGsi7BFYqZXjsvL8s7THHxFpXSdwti93u0uFa
bvLsh1kd1uYWivtyQOZr1OksgKtV+GZyseng41jGIja2B1II/GR4R3SfsPWoNsAz
8pFEu1+6FNGbzZHoLOgOuQTOVNSCf4BLHtwbKXYo7y7N7L0WGlfiOX1/kPY6IS1E
r+CkdUmVwLMvGKxpdKinbn3842LIi6eEUADdty+NsBc+DL1K3KdQrK6SLEHUqA8d
znlwTY5y7uHh/yxaWxDnfGL2UrhBreU+ovEOIJ5M/KAsNh1N06zYn+leYFo6yy9q
ZMDuxGYm0TckmKrMk2ypC2eVqCWW++rKL1UHrG7wNnqrVMZiTAcVmVcxkN+y3AJr
HO+pN3D+ilQjNf1UCJxEo2jNheIy8OECnp8HaULyYUbFeLf9DjmDvA9HOkP9uTZC
4xqKzKMMUUKiFT07XYIIJYfGuI0JjWXrmCqw1/Y8SURcedwQFkRnwdQUsDAnuCZj
VMw2919twt8GPEDyyF1Y3a+0dIV1jcT/8PqbQAqqeSBlCTRVDGoUG4iQRMU94qMu
JYZTz2G+4EPijhtGlgDlm8llheOLigvSei+/kWJXcMDMO7QvygPOmpNmRjIDKz5F
583CVOmMPy78k2R+ATmySXU5paUumzlJezYYy4zm7Zqo+sY3uJgfLqHLJi1htS6O
xF8lx8lukZ2gRC269qs791mhVAMKvwZHBunGUaIeFQrfpE/6mWFSVGZWVKEpWg1l
qeWJ9oyxpqubZSLkO2qcTjHnsnSD3LMzwM7PQfxXwcFwqAvOIAztIldzU2Wsg87v
i5LCLZTXpq8aZUjAjR5LNwtUweqoE+rxUVUJJAsc0JxTxoYaJJSwDZTYyk1yBa/x
tPKPlByv2KLCd18qf8VhhaD4CN5u70YdLa7fycha+PTlAmO9/C0OkbIR7hb9kyfx
S1kbOaLAfUOwW5MTgwIzlY/vSYMZ8Z3KyMcWijz9u1JEZ3ioOP318E/ghWVxWl0B
gJkKZd4/xWWTmiYV5Q+DlGNa5sBh4ZvSP0ElgyCKpz55ln1I8pie0BIU/8XVqJqv
W5TLPFaWtDq05zIuVTEIXyDmjdeE9BNPmE82cA7K1AB9O6F51408eMBy6okvs0Bf
WjLBtMc9Q0c+PmLatf00u4PInfQ6LJG6QAz5L3/0DChBueOuxcPIr6FgYvZRpxdN
zPbrhPgL3dqXQkiDVmPPfyXXDq+ocRu+wPQ8+tSTyrlxP7Q9hn5b6mpnyQPSjIVX
hDPSci+GT4ey7oWV4INWL314puDorL7A82IG6kvOlA/oNNeF7C4MSEmLbOx+wtNr
bfVia07Wvf2SVUU9RXayaT0xFtS9d+heMoeKoczDa6p5oBcciP1O39pC7maS8zZ5
8DwMr0679WhFV+YA/z3ar27DG4WLdZUhEgq0mUjCfWJ8avKpKz2O+XZppz7Vv3lJ
AXlMrAtc3Bd+5xDiGS2quCCn0Ln8wgyMqYa2I/z5Pj51HpV6KorWudWDOj4gG/rK
qMSfJHB44cKHX8CleSlXgviOq4bTr04ltFPdoea5wxUmunv0TzzDQadxsCkKE2EP
A04sJ6pj7vMGHStqI/FONoaymCPlKI01M+VOVA5oJJ9IojVrVZeRJMpPOnIHIU0H
u6/VynWhWmK9tQ3Lmg0+O2CZzlQ2EFp7ipOGdQrklwL6EfRK0o0JYFZe3jbMO9PW
lcXKaIWn1a9WBObW0S9Pg83qvgRGqN5KeTUWZlntG+AcQBt4cpnakEXkrSL4vBkJ
ibmI7kyXqjuoNLGmCiTwc9t1rYUHhe/N4xr6bULB0EApPNR88kMoJYobRJ9un8zP
CUDzo9KCMBRcWW64M5VkjaaByPiTRKPUIMzC18XXxsYjajcnlKWqWnlUG8h2tqYh
xFSVOV52mNSYMV4qyw7yaTC1IFciXgNqbGiwPd0otXx8EyQW0jD//csfw+DW4Jm8
Z5uca2YlgLiDrU20ztttGUXzkVIH2EWlvzE4ib0L/zGPnKR3GnqTJBPNs1kcQQpz
zN6Al3sipcHWkaIXYr0DcPT2MLlwX4x8Dmb239Fwqde8TbtiDYiEHT4A053aTwT0
UKvXz35jQr+747LZ3RJhXSbsI8BSF3DKWdoey5sw9VjtzmCHGqusu/26CqtJCUOx
Y4Ax44821stUg2N1dGirg2yOqhpdDTm9IM5XWOX65cGNM6kMpCS1g9ZgzSmPBxqt
6OOqntFQtv4OY4/uF6CXZ3CrMq/ZVTlCsm/WFAnpTZ8frCEn6dS3kgudKEaPwj0M
Ob9tO3gvh/WBRgL2Xux3SnZ+0fCAKR86FS9QKwaWg/nojkT+Sd5H/tdx3GTWlaQP
CGNjm+hJY0vlFRwPgDL8Pop5UsGpY188DHSSz6LXv2X9L4ot0XyTcQRqE9YxhROf
lWl9q1U/dBnGaOS/mx9z2tyu+mZ6JTp8A58xQc3UNFj6/AkbSeS8P/CMDRQy7Dx1
sEov13JE4Jlf1MYlIf9K9byQyMlrF1jgWy1Srn0xDvnWcLJkfCDjgKkc79PEJOcH
Fzt3Svvt6dbfWXcBKikwGMddocEx4hNM8RLGus/aMq/kuN/hwDAdXMVbo6BBqjH3
yi7/XPB9TjW+Mo6nRh42USZL+7LpP/K1IejWwlIiVn6TJHFB+2hT6QDv7PJEh0ke
o6bM7Q3gGLgSEF50b1fvU5pQgpYDtn739vT/8y26weFmTuyKy4wiNSx+o9pCEIzy
mVeyPvjfe+qRTnf3Ct/8QZk1vJu8nIjk3/WnTGkeyukej2WMy5oZ23lP9K/+UlCp
aqmRjMwP2OSx8oQUAExILLFS9m2fna/D+O+ENz4TbxnBQmyEp+yno2ehj9cGBfvt
5DvJO81MggMnsD6vn5CqBc0S5mVulvQnpxJJ9wq2VGrjYqdpafozdS2LNcgmjg9t
AO7cGBywFTL4uHFTHGo++NHglPEazWX6BmgFGtC/7ahmUdJDAfJwRqvAq3mZNJG5
lRXoJVsOpJyyAtxkAHGOzi5P7ki/COaX/aBLxZaeHB5cehJq4Z3UkEFyr1ZseGa1
J+bFOTjdOQ2/PXwXBANSnCh0Ev2oeO+kIWsLi9e4x3IdTqjBBQHN9G9KpiHl4IPA
H4cq6GKILAxHYKG3UYO8mQGjry1Dpxuddu1aEqAyRdW8m/d+FfCbd7rSS8BVL/Nb
X6BarHVHE5NkMsoPtjFc4cwFRCjZ8ijeSbg3qNRE1ExSY+XCCC4+4dqjacrvVIK/
s/43tYYL2l8ufWKor+B7zhxds70uFuPScN8zBtAkOZ4Yi17YDZtZBdiGBHVXDDcg
wLrD1961igHzCw7K+d/2jKhdOIv/NKf9Td3U1OWd+pFXRVVZGFW6qZuVOMW0IkjG
4iQRNR3TrE55RyBhQoGwHELFcCF8/iiljCJLdsVuhXP3Kgvs/PGtuRDw3qe6UP5s
V08A1M9/3tiZkQKbCLfvqCKq0rAZcOF2NiAO04D9UexUjdJ4W1gv0bIz705/DCnz
474AeFnQ1KafsaW/zQBzKKjBiSbpLKOgYHXVNE2cmgpavUJKivn5D+7Oh7O4H5C0
VabdYh5tJSl1alaTXKFtflgOzgwtT8KRiNuIVrZzYdp6sABJ/HQWBi7rtlPsJWw1
LZBfySI8cJ1dbAfuV9AkCn9DCm3av5pxA/3EM4oWlFy5ZVpAwsS+a3SBQywsmkqo
lRUFDZZKzT22PW3G8cuYKrpSJnUJtHRu8kApVqlYUkZWUt6Bit+k0bkQfmAmPnBq
7k9zUmiL4nawjjgnPzZNxHJ1zHKy4/RtHfsqVzt8C8z66OsGMVQ37wPDUQ7LuaR4
Du7XGniVF1w0lZEI8Qzz1f36Hk9SC7s3HbjOKC1IYiFbk9xY4LjTzsH5fi0EWUKQ
dVoQD1nx63e/TLaEd3oEypNPyu6bdqdvGy39MATSN1aKW27wS8PQnSBbOK2wrY2S
uwOWiFhuUS5hXKKpa3cCwZvZI3N6hVJ4/7U0HR7YXHr7fzW6m3AzcFKftui52BTm
XhHIUw6E3ecnkWNpnhFEfWIEizgryrHKPgwWOsTHbt2wL3zJXmW9O/ciMJlB1Ate
YmPeVeb+0jjT/uel2BvuzePSQxrgoBfjDf6RENuA3vL3dNgtcleI24FGz1ezZIID
cPrMTlEOn4PkELXaZr1KG2W5UOPpun4M1Tih2EvkqfrfuUK1Emngth4IYzRcsVqe
v6QQaIDQ7eYtNPKNLYvxHb4B5zvZ29fWXlNyjyvqgE9+CrJ5YtS0VR3ZxdC4SaX/
RXMwjQ87eK1kkIeAQ+vel4e+NUctESbYyXdWLrRrDJ9/a73OFt5YhvgKw/NJCV+5
vsoSoeG7SOIgNRFlzkYBygTY8XG7qqLtr2hZ9/Svj2rB4WOWMw9j/pz+7uNt0W/0
8aXf+lQstQ3KALbL8YkzTWdgUOItIF5iFT7z/hHzvaYt4S0qUaOYZaK51vDiZMcJ
fx8qUYcfE89jsE681WyOdpO7j+t/hKVJOtN6hxMQLoxwBScWNncCf4X/h8F2+56d
sHS5oQbX339VAwXyiJ3Eg7IKtmnW0EUhG780XM1cuN4Bo1qIoqah45+7SYiziPfB
D8K3Nd8GKq/XDcpNbMu+LKU/rFZ61q6KVzMZI518uUf6iZzuGjYXCUkwbMsQDmSu
HiV06xvGY0y0U3OCtd9a9Yurhd7bA8pCzzDhlzP6jBHDcl9fR47Ov6TECOLmL7M5
Xd6WYzbPii3gClJqZy3SKGvFaxbSb0yCQIhA/NAxo9fvXOm/0RYs/jxXBEQjAVDi
LK4RSHCItzFzRfJ7o19Yn0TGQZSXaJH/LHAb8CY09KXzRRw95ACGDaF7dvLeQZsS
H+r3HSnLUEjDMmdCVa1DM2D7Q7xIJO3M0QZTnHRZObz1BTh9PcshjTXt4dcFdNBV
qoO477zXwww3qNmVJuKiRWGrQOg+hGjzyZIqOnh/VGIl/c7GQLd2DG2FwBAWCBhh
lXFGI4miEHR9l5rOlTUaQYiyJ5y8v5xQeEetIH0yePkOudujUJ6RPHJozMVCYeIn
s18j1flCZKZUGNPKMY0uYMGIqfGpVrl6GsOpQeSY86NcExn2g6FD4078i/271kCW
WxhEkagjA+5Vdc2j/cqJK1KD0Qe/PrUe4Jl9SQIxtJOhFHcxqWk+PZO7JxGJbo67
rnpPhG3hvTjY4ZRZQcy2BpT74UPqIkoo2YG3yFIwgDjT7d61vZTziutWXx5h3jac
8CEbVxrLZqZUv4xc2NtNeaHSlJsvWJcuK0ph1BRpy2+NdotL91sZZaPeourqtq77
zFDqAFLm6kaBK5qv69geM4bTlP7U3vt7MtAatRAWUqCx+hUzJqpeUzQp/XGxSjp/
ZUGpoU/aGi1QcCHF/HkKird+KOnicIVuJTuh6jHeCq7k/EzdZBZhxnorDdyIyGOM
wk2CLoRZoZbbIXowZ+u6LHW3wO4VzHSsJr9FHK2/YLcGVNUWLae6xjZmpYcS/daK
m4Fg8j5I62kI2GTvv2E0aqCkefoNCzyKjaRFbfgcKAKvyhbmVtoWwARtIW5xRCTW
DqH+u1rPhYSDVGuYgLU4o26vbHzo+hPZbGegD7i9PI9zRPfzjtxt1q3rTBt/n4oF
6DXT60GaLbunKsaOaTRKl7tY62+b1TbRkFk6PVN5N/gu/wr6OiJdd6iE9JAi7IWI
6jNCp9mNZv2CC0Z0dW8OBvWiVPZJEUCNftYNMpLzAIafFtkbjjoAX18EDzAwm7Op
Bfsc1VxBvD7VmrIJ4bbiRM/6D/jfeSVMxVUdhwEboFPEecByF7w9cR9epWSdCpz1
59DnLtHnEAfKBtJpzMSat7xZdn5v8bJ9g1z4/rcEMx63/+/wqV+MQCc6zm7g3vAR
j9T/UWW62EO0ButZi19mx3/zPyFV3YGailoxwzUJQ0XTsmZNsR793gJNwoFLnafP
gJJ7tkhLqfIBzi/eYG2mdZncE96Sso3d5AfjPfbyp4fk4/ptLvtOFss6S/mkrtCa
ijfWPkmrpWiZRm2IJ71KUi8KefMlZXeWGb16cb4MV6Ddu2pOnlBKW3ziTUGvB3Dg
DZaEKhuZVXcUVwZslzfM2RfxtCiQrl1v6p05kRuv7/dCIB1VOxh0KEzM9RxS05tf
RQY8atA5y1mBeBWSW9jnfLYyjhfWnquLcoi61VRLSRnvAK//qM2XoI9JGQU9lXdF
r8GaGKSdFKlx2pJpbRwuzMkc/DC+OAmq9t8+2LGv2zuioM90/ryGXRiUWJTC63cH
GTwyZmxPFA6Hzc2vpCWZ8+/2qWbieCRl4aWzbSOwEbhRrbQVSmeIvbkcnYUR4bG0
LsiQcbjA/pVMuX7s8OcwGIZJY3FnQ0tlL+qkXWeNsGuELI5E6Y2UwO2SrFOnymQp
LJQd8dkbNjWZFQRJ1c19dFD0Zsabgi7Uyc11QfyPxIlMlZ7iXuFnNO6gZb2Mlk2t
tz7XjRoLWPD3wB05rGQQddKu3fcTOXHRwKcNxcPIqpwsYlQSBYXz1TF8DDdey05G
8v4HC6X8F+Sl+bSBusxfui5V30GIRsE3R8qf9nmSVMF54NxT+9daOYWi/fJBxc2d
RQP8zULmYht56z+Ap19ooDwoj+W4ZMxx6XVPpaytXDfnXZPgBxwmmeVKVz5dXCsg
fqln6o8rlCYR8x+nnKCcAaZ9lCLeaG5SEBZmdebEkPhnrr643Np0IZC3KYlJ9kcF
nNARrNr4tefH8yYHbscUmOV8TLqnICQbqVpwXTwO5w/Qph2DSo+0KXhOpvuVRx3s
LZFeV7Ko5anE3RHTpn+Ka+n1XmlCpMaOGdqy/Swu6S16ik5mIPRjoxMmgHu6RkDM
6t4SXTrMRCnfIoD80Sk1eTK0xEPzUGCWtwSV9kG9yt+r3zXkkaGNJGzeseRgngix
8LAfFWaTVSNylDKIuduehRVLvWW/vhrHw5bN7elGloXwwAIjCaF9MTB4BaXeUsxI
+NT25rzJo7nO05Wh2y+c4Zto6PttEDEJLgg7TIkOGVaJrafjHDs+jtb+2tHBgLLR
qKEZj6FEU91HdEjohHOm4OHSW01pberJVicc5dvjmJXsDqIIzlURfoeLGWbwrSKT
LJJBir/g9uPdu5zqj/Bz6qsAScfMiN3nYkFEEJRM8VJgr0qypBaYNnM6QU07CuNp
EsQNRt6tKPA3+QUOWiIN8Kqr0Z+j0hOzedY4e68zUuskUhRNqQhpo1DpD14F6VTU
1r8rsBDpXJbMo3lIYiWSQTE3EgBXe74uzeSth7C80+eg2+4qgkzxv0iK+4SXx8Du
QEnEB20bqdtKL6hOnW8MFy+02OTq/9c3oj8sFrIHO+R3ZfAw9pdI0tluoaxQhbW8
xRdQ+3gevXNmwD5pjQ63hRVRtZ4m0F1ghZMaCIzcZQ6+x7Z1ZYNqY96/Cz0BDg+p
IeDEy52C9Q34kmUSopEQlOeUaKmuZLMvDZ6wF9J8nwv/MkZngdmbIY+5l866b8HU
hvol+SVjlvx2eQ1R3oP9MlzVoxI2IklRmc5stVgA0JRI7Tu/z6fn0TpLZCLYAcmo
rY4DDowi5o3p/PSe1UTy63ETeIRev32XK1TyEIkm/3csC4tVITtfwQlzyiek363x
X5K8trujJAT4B0MsFm3RGqiRWq64+d2LzTGYa51osvuKRIEQ3ng/XNq/0jjmjj24
dP6/FXVvXgoIeHzKiLYAVBrVUP8JFy4SpCp/N3Z4GYtS1lnex0tHVmgQ+/s5vcTV
lT4MyfVrYf02oByNctV64/TA9ym9F1ZKe6Ppx0rkXlE2skdlJZfQYUWMGg6urSLy
ic8H8m4fXlhzLizZHj6KdXjPzwNBRQc9HybdspvwF8ygElvzp/VU6pxnffWL406v
6sBWF1NFTmUQA/GtndzkHoWZgBsCGPXS3bmWCrXy1GRDttiklViFc6Qc6434LSFD
Iik77t6vnjunLhBB11uLSPX/5R7YJM1BhQVul+dQ7oHawBizvJQmgnkr/y8/5Bg3
N/lQ6P9oHvXBXPvOKQgKcGEcvQ/jtrQ5dumWGD/fJyjjcbLZj4Q2NWqVHBxJVlSu
sdQ3FvEAloLyvViO00p92weqiJ6buNC+jq5Ej69yqG2aKw97Nyjh6CwcJdGVvusc
TnrybLBkzSvNRv+2Pq7DVmJyFPtR65NsPw6bgatjd3Qk5QwUDNJBxRu3I1VQxqWk
C26iYk4AwQhEmtu1J37BEOyeBY6t3N9+rx09tH5pADTWjB509GwAyotkTo2WOSuN
AdlvRuiU3YiGNWtG6cciC1Oo13ArojgzcFFdWdWBWbWvCYoqMKAeC4g1Joi7QWtx
wQBbt98Aik/A4h1mgLs986i5rDW9g5CTjOOGFysXnhE3TgTiHwo5CQxnmK3Tp51+
7gPHwu1NA4PHylTzhvrdhYUY3GmoMC9klAr434KhUWDFdmreAR8zU6Xm45yK4EE8
FxcS1/R/SGyL/PD+kAJ+UoywywNjed+58T2O17JDGMA8qpUcIW2z85iRENJborVA
uvmo8bi8aE4RdZQT4rOX4HrRbnmS1x2ZqfjZPjYOZC3sjVXsnW6kWLVsxci6X1rC
hQfsmVgJkd7Z/CiwnRr/7wJ5j4/xhJ9tALV+lQ26MMF4OPe7ptmDRXkM7HlfDIuc
gpZf8/OlqygMYLDisZurVxh5JkF6YBLw5qxXuYOIjUC1wbXQBpQeDQZy1YvmNAXV
cFyskOAZIggVYDZtUYutlVvzKz4p/gO07RaVa8cLU3i29HrZ7YMr0sRAo1HBnxUD
ek8cxksOqmnv26+Ztj3c7pxfLkxVw6UkeI5eJSVX67IrViCjco5pAaGgHGeDIZ+D
N8p7hN+lTgp+SASguPtygtbMKb+e0ZVYkznSMO+G55xhe13heaKqE+m0xxguw+gK
kgejTo5vhHtQVftcAVawbiaxBk3hYwTAt7/ovA+/w82TBOFqlSkZehvZJCrCS0xK
1bQcWoh1SFAhiO50qw7p98008/C3T8xm+8SbRH4Dnh8CEFS2ELd/RsxBqvoJBuli
/1iw6wB5KsoE1UBFAMwfWi21eVsYZeEzFsRCmYAJhOqMFWmr5ppbAT7UFM7Pk/W4
rMeQRKgUtHL2nouATRiC4x6mkP4I1folImOn/OKeQjsmRun1AMO/RgP+gEk58f7P
jzUKcFO6Zrlt7O5KMWhHsOIQinY/A52hrHl+nfSiQEVrI4BQDv6C++eiD0iUX3Uu
hoC3xSFARwET23jYJ94/8wOJ1KxJEjezgtiaEFqWMKE6orl6LkNhUPBEU0XAsQeG
XeA5PHODzWk8F21hWpYeAcdqOjWO9b4awEZpD4dWGpmWQhmzDrTTIA0PFnnjDyPH
9vL267iXVs2HEpaMYH3IGVTKsOc3WIPon9Y6UkOJ40JflZnQIE6+/adDuW28thQ9
6xnbynab8h6NqgRbQ1Ij7cWLmWkFMj9ThhfSZPQmmjSRIO+dqAYjNBktJSWfq230
HdD75be94gU08Ymi2pG8WQqwchycTsB1whMosRRZb+23pyPXbhoFliWK1poTvfy0
q0xaxTS8R/4iRsh9T7uwD7Le1iHSwvi68f3FCVK6FwYvVKCV+RCc6oTH2o1LRgFm
gDixpnM3OcD+hzAKFbEPj6Kk1iIOA0oJb+VCuVOK9xvgZ4pAVX5KdLV3hWnyx/JM
G97XgLULkjlShNW5yb6GzotL6mtlySC1JttVS3lnzZht7eiQhv3e373Z2d8Av8FI
fkOUwPFAIPRYHaV++7X/YRD9Vdx29rjMcTGQVO1gQ2nO42VuWoKBLo4drktlp07j
alq6k9/wGfddfOzxdRmax31Yu8qBKJfDPELKt6BYxmYxe0FWUTNAYwCfpuQApt3R
0DiexnNsyR2gfUYku/No6frSXMDYGA0VKOriT8/lKRjVKi8bpD/ByR/tyEWcLrA/
ctf7lTDGHTg90wohRPucMjrYnpwT9iZWdgf0fzgzgCOBG8Tq6hcOsVFZsj1Y/cGu
T9JiEKXOrqhCDKGFM7mx32unUGYrojH/w8w09hArwMiXooVg+vQ9PRJD0++749TR
c1k6M++r/bINvzUh4eDFMw06EBzZsB3Nj+YNckZrXxN74aqnbqoB451Y7mXfkxSl
z06cJJ9Rye1xHqNeBmIzaVTO5hvzvG1PeoKd+Z4Nv4ZylFcYvwppTrXI05Zlacrd
1C7tf0H2z5CDfUezVffqcGRtyo3Gz/OFpmVnIX57nuvGTJVfIa+yIda53kTk/YvY
wS8FSpz2K/itAqE1JN2+ngmaMtK7B7b/ZqTt9ZCbyB+b8JHxmFGtKorrZrdqFr3l
WaW06UwSzaU/VeHiIpF8O34bPC7McrmkLrM2Z27bpCGDoOJrU4yqxobBofyNdI2l
Huy3o0fUWpfcMYTlqLmHvQ8A/Tsz042otrKK8hzTo33uvANn2/oZwH1NlW7Y+t0p
JRvJ6e5ML4aU5RoWD2K/M3gMXKZ8ADgwER+H4pt6JaBIr+6u7LO+332k4KlPRxZy
jI70B5UnSPHsJbe3wRfx2t9i1U1Iwr5HvalwmPn28iwxlM1ddSsgtRnQIQnBYJD+
yAZA2BubL8NpbBKZNSLx5IQXgen3t6ILtJT8ilQLmTIiGzEAAgIvx7ZTD0Mzpf7n
qGisWlgfZKhmF27k/mDhSYzxch4OVZjm4KWk+LzPIbeZKIm9sdVt/eJFIhT+NMCH
Vyus9t8YUvr6iJVm627KnNVdBintUGC8JDiruh9mJSfBT3Q7+pBjsfHN0j4pW8q+
6f+uvv9M0t2JNzsSo09bB+59VEhP1DHJJeISpQxq6RHDHRLl9t/xZPhRLdQ6Kd1A
npCn61Q7kOLv+1RhERyhiZaB4oZbqVL+Iq4cLfudPpvHmobzvuLq5mDQwHXo4jeZ
3d4pE9Wfrx1QP3cNtOqiPyEjBHZmiXgLEWcgTHSWjuM+VZZwC2J0/b2t4m4jCyzW
nJP2NU2gJq1ckI00sLZQrWOYVxfdbzZhHDvLKxMU15kTKeSnZYZGYjyNi/L5zAkW
gB7/Ar9qfniWXeN59q6YPKeJAkKy81dbLuKF6mD/MRrcYKJgnelFrXbE1WAojA6D
f3lkdCGqb/8uXdIcswiNmoaFVN75+C8eMUt7QH1gKEuhG5Owc7R4HaaOaT4syTp0
bZhTPMetgKSEJfCIFbUK22i9l06UUMbFoba3ONULSQef7EGQyosJE1sErkOLYDMH
krAdRSZ75NI+Locw+KxyD3BaprcOYF73DBw7MDWoHOGNLxtqGyfdW7DwC9BuAHVo
pn/jKGAR8zyIanXeYeoV/bAvAWGoGO7yQRDK7Vzv4GMTF2ndCbJnzf8RlmvgRaLw
DxGp9WXxdxR0DxNs1vDcjM19YZyIglmUMGOOGMZdq0HfviEqbapAGjWsqE3cg1qv
tJs1I0cIBUiJJEu1Imd9/amtX+uhJPSvTZACKMSUb/KCHtBTK90ue86sx+c8F339
KURPYNyLoakObihcazZW5RlEa18IvQIrUFmfU32GH0A58tQ4uVzqXx0KbRfxjVqZ
bJPSb6cR9VGu5U7k0FBU94C77+lsf5SIkTpKpJG0y5Hdj5ATVOH/OqfoYRABmZNR
7lMjlyD4MMt2RZw1v8j4jSbRCjPYfPjFUOOZZfbD2Hx83sZ1rLdy/Qn7Ji0NsfGe
An3ZRalNViiwfjPLr0+JdFsph3qRcBpMv3xIhHuVhisKjRu/GTNJc2dgC0d/idM4
EW24XVpgagYSzZlVnZC7tL1l61owqd69TgrlpIplZEjw2msX+0evC279v+1WYG0P
Z55AfjA3OxqNjqivIkzb9W+EuX+AA6o7Ltz8Dg4touQwnsWaqFe54wsORr4m3Bn0
rex6bedYPcFsQ8OpyCqVp+VjX4yqpCSFeeQjVHLy9EPqu7RBv7Vb+Adg1qMw+Coo
R9B26lJ8nf3/NVJrc/8RsV+Z7KeXBG707DIPAotWTDSw7DApDkYbxZrUJqV/LXZO
lNytu7HT4iOWLwFThQKXgdGWDAt/sPLv0GpBnQInOIUH+QLX6/ea4p+XxH5KLCHm
KKfpjotoJ6OdIxUO8hYdCgVl95yJCScDbwCOItrhxjdUseBdSxqg6Xc9NTxiTJ2Y
7qkPO3bXuvAHkwydc0PUAXjNztdTWa5TqgotOvwQ6xm7NrV9eF3whzvLxVg4Lrdk
tPG7/L8lbB3layfkZkR/KbPKrBGxu9L2+E60fViGSm8622+a/KBmkX6HNY9+eyuo
BwDra00pIX4+s7ecB54LmqnB5zY2NIDqzufffDZAkkH70I8u0mIn1opjIyLUYWRo
NeiKqyM7Zbtp9hZbUWQDgSRCzGW/XrZwKeahkeHKaI22BqZFgzPPM9XlGO2wNaby
xuZIYGpZ99+HteSddgjS8OR1nRUlHCjCXHR/Jmm8VGc/N5JDA9CsMuujN4DEFJqG
bYi6p4OCpFhbYWFTlyfc6lqMTBDuD4nbWAzG4NOqY4iIcDgftOx0XkF8+HpQ1HK6
CbjL0vKthkfzmggRuAIgN2T3iBv8fjyajAwQPP8mkfis2ahgd0XLWQM5yhCHavqX
8LtaRCDgLQmwu03TPI/Zcyt9EZn4s9WzWu8UivQdb+diE0qsyVuadFofSYT/M5SV
sPHYHvxjEzw5BmssSUNy3zNmqBLhIABfNFl7vwqDspVkWB3oIomWA/2xy+q0MxVF
yvUs4IKbjQI3Qttb4e0k+7pUufTzDClrUySWMs+JQlM98TmdIuuRozEmWrvPB7Xp
2tBMbiYeK2+1XKlcxmHxKrl4nK8MtpOTMyiH9ytzm7oc2nFLZVhHSCwyJ4ocR1Gi
/gN7vZw38hmsTJOZqDzikHyc4xftewOfzfTU6vmzy16pxBsT/4gck8esThVrsV+B
1HkC0oJoSOAJEgxbGm2HLn4Qk/93ZATcU5jE/VWFB26HStf0SFnognE36biYjJyE
9Jm1ys8KOBEqAXQP9c0pi+vP1wW/OZBy1JqoTA2VkzLryw45Lgu/VO4W8dHtc8Fd
shaA5+3RSua5kScwl0R/kJuQX71ULvrf8IpdAgWEl+koLELVigzpcDV+VRZvPBBU
rnXi9X2QgSyGJ8fUbfR7CRcXeG8C5IWs6AR3H9a172ZeS7vnCqHK9k4BetId57gM
9PSBVhk8y2D2pRw/us8PkPHPHPgv8f6HYFUUIr+WjeIPMkdWBkzJPcHdtkr48hHm
JAj9UVkFjBpI74vYkdFHXiaB+ON4c/zIGcQ+YvQ6iCGViFipF8lLocHeGlI5+XV1
GKwrroXATSJ4Ao8hLwlxMAo1gqyFIiPyS4eUuiMZQ9jPIlcdgU6CDlWCJeyDtTvJ
ykhdhGBB2ubqMxcWxMPkwpmtCI8hDsPPRztqUK90A+hH3Bp07K7tovM39dQpoQuq
HJYYuscw2z7OIn6iG7xmhDgAHZjDio2tV720tkuleW+w1nnBCZaQlN62HrUMB3Wj
dPBnqjnsSHiRHHDki7PXzwBtoR9wFigm8OGkgzfn/vOptgNrEBRjr/bV6rltwOi9
rkFDaJpb/T1wrE/MKK5dAbJ8UnQR3pLrirfo+ThSUshrEf/dqHYOkv1PKpyJssMA
3G1ZulVC2eJoJwJAPhwKb6ACduG40rxzzyagKPD+MHfw8VUAtA/aLv0RFaiOkxh1
d/iPhlUGUrBeAOvDK30+dByCKl+zj7KKpXvh4lRo8zuzjk0CY2qUpRJxpE8hjg8H
kEHzMYBH1A4kaIS29iTRJVwOtSROC4f2pQ4hTRFjpFgtPZImgpWWeUIIkaKj78mE
0jF5A4Owl6NctEiN56AwFTUkQNImn6tqLOt3bokHqeLhyFuBAqignbTOBcD/1No6
3I8DKnt5A226DRYMsC2RD1ACocNASwuMyaAj5FSsuKoB/So9qAjElh19DyrgC/p7
b+dbf3Sir/QyNZQ+HyT6wn8fFIWRmWhMB+T9IWeraZ0/hU2VuHp3yJ5UGL87aXj2
xz9hk2EMDYRgr2rYzIq9V5RCyR0PHJiOLtuk/fF0wqjiVtp0mUDfaUDLiGYe/8QD
p2TPT507GzAC11b0VRu75hCd9ZET4QuzO8hf0aMo+joAvXaxG/ehNmegb/jErl+g
FLmwI8F0g29KIO2YpHuCtffZDaZrSlohdOhRBRanuFxgA2sPUFKbTz+Wq7Pm2EWq
sI6VXQPkWHuoXXkXeLzlrRYyblUA6xXPF+34L+ZH/qfzW95IYqHBGjCZ0xWn4KLk
3cr80qXSK+0rfLSgZbUHbkQhQ97oqtpWC9FmnH4CyMuIwNJ9vwPYaZOqFZrOHZDx
3XYFFUGXADAynoqNyhM/c7KIb4mV1kI7v0YH0zEzXGiYbz6ZbFdapf7evx+ciT3p
f0y8Ep/eY9rDhLjYmRGE7ZHJ4y2kx3Fs7zIP7S3l5cn/L9aMYnF5HVfW2uSxgD6X
MqDLg8fBY/EHsX3gNbMTTtDO2zRiTn2A45QNrFj9DPUyDoGwa2F3VctP+Qrn6025
8ABwg+5AxuosrGCbS1yt/kbaTHKXcTY1LMvgmmxMSfVMzLnmITv9F5ScE+S8xP5v
9t48eUKay49Nmw5ew4cTA1E5UjMDmC5mBvBrbCxWkMrt+D2RA9Gx15kdn010I7kD
65/Ygd7UJiw4K/ICzsVS6zXZ/cS1DfvupzXA2QIYLMJxOq1HioYY8KApjTEUh3Zy
vNMpshQBXhZOc7tzeT07gT6VScQC7qySx+UI5ssvOh+1m0vJRviy1CqJmyE+b+uM
wCSE7sSakLaArmwZEQifQvg/P8GBlmlYUALx7VJjRq0QpUA4v2lLqS5b5xVN38ri
2mXnRwx218DbIQ86CajcpmqrzjUr6FuIJZybUHCn6VDQTCjE2Y+vTk6Yp5zjd6J1
EGqAFlxjkfprOLOfhsJ4E5v/40wVwfp1dffwwPU+7jvvHegkhrj2xgI2/pXwcvEN
DGJA1zEEAmv2NB/DombUkybzB/BEMjROpAM1B18JEqD0IUboc7XoerCtQ6fWkRcw
IH6sspNWfZmOtXvjB2gomyN8UaWK2KvjakBhCChLnUjEGHExdst1lzP/wOcrLxaw
Afn04UAcqFO+yNcXiARqtJypc1VfAptr+5p2C82r1jqJMIjMAjwZs7EnTxfpZeNp
FZFKlTStoA65NPEbstlswiX5SpLaxCX7nT1z8WFnC/bkSoVXJVE6JOGDGekurVwz
TzDAt/6IzvvtihQ183z4CBG99eWJg4lihu6pfgT00F7kaR5K6sQsrirxqWspln9s
4tssdAEHXyUnpqZrSbSSMr8hZL+SV3sK8X1X0hm5TKQkIPhGedXflQX8jbmYyLbe
N+j6ejZRwwY+Sb6eZMY2bXtK3v8ISsofc2AaEXDWjlx0BcDHPjrFHGJZBrxbLV4S
5LfybKgaZ0rTkFctUUfqszaYDYZfPLsdo2YpPgFqBADzStsorOQiq6TA6GPQS4I2
sNH6JWk2xJ/gx08oPCzF2rjh5v7AxWh8H4qVXWNQK029AUIpfBVY0XiSKo/HlzTC
AdM3sLkiCLR7TSbj8gziC/VDauNtrY9oDRhTDikiATv08DoVDDzy8gTBXAQzplZb
gJ6o/nDZWs0WzS240CHKtI5hpFWDnrnaA6/gxpa7nEYFVYXqO5zTVeRajniPwYmG
pdzzrhtdvO3watyX+FFxFFgqx7AZCl/rN0g36DDTmaO3iime7Ys1/6oLucqCM2sv
z27n3RjZtqbyGTEDycCyayPRStyFRNDQC1QAWApoE2gpGzhMOqijCxhVtN2Xqul8
170cJGT8Ieo9qZCY5qcM/jFFCUmr00qpGe5YSUuuhJ88ZKVpPob/xV9+faOSgN/K
YnBb5lyeHdd1TcSI40MRwi+dhzfWRuKUoyKXllDKEVvV96pioaMK8TYxtGKOBo+J
fat+Nxmhxxy9mInUYZcHLv+ytKGNQ2U5sGVpT8uQXyQ8j0GmqJRPEcy+qIrxSCun
PCBG8/MCq4/KPxdQ36IH2BwL+AEN+tOCSmlVIc2+h18QXLiGad6YeAZYjokuW120
yc8rJfBR4D43bR5g5aAtDZ/l5ffLR7a10No2J4mJdU3EXlJClK7s+pEjp1RhFsFo
9a3bm7ih1SNVrLDyNYmrwGVpMdUyQBvCdIVMJ6LsU+RInwQk6ZRZwG/hArdNLaQE
yR8LGUJxUArFeg45CIrN5kULKX1fmZMrvthtRgTYGQid/RTJsx4rqhlE8Cxgd5ni
wxR0c+mSKTvPbJh2QV+0+Nwos71DQhODWYN8Zr17hkxBsobgVJ0/5OhREFhqCgr2
09eaPvM4ZBSXjNXvRYSFyEhZsoYX3AI6CxN+QQuaIUHorylGdp1ZQ0TvuNrE22UT
WwP+JmfiZSSQ9MmF+eMQvzzqnH375DCk7+bqKUUBlu+P8Tjih6yOrmInSXrvswf9
GvkD6ciNPuYxpR2357s5uT5klcNP5DaHQa9d/O3XL4BOcnDshDA90lo6F9Cw2YPt
dXBRk9F/mWAjTKzqXDSm3xVFqM8vteC9TrOeLIczsmVHrze282gNy/5RazmwRJpd
J71ixiSb8SZCMo0DsnOBa5mQ6wEOtsNlfUkJ1qkZtZwOKJ/P6pbkKd2GvI/gaNaS
BQ0ZODn20J6CmSvtlii1vDSqaJsP2TBY0IlrPAhC70uY7bxxn/jMZeRcKurChKO5
y0QphVLo6mJoU1DwENquepOFljyylqycQyFj2sfXrj26WOpYKnG+0dBqee7W5zYj
0/Z/bB93MXJneRTTfkVdvEX3pGkUxJB0OihRcFPh6ZyoaE1v2xxzDk/HP3P7Fu8g
ypIOAmFtIn+MW8CcIPH5iR0wnXsOATEsCs0Wq3TMbE1EWzN6f3W+2aSmT1xVBGOC
OZqlSOUGBjutcpUUMFv+8tikIcz8akHLRcTc6AX3yfkYR/jmtp8N4gPK752+NwRC
vPddb0Bt+zn8pw2L4K3NCNTUR14Sep1pMIhY6WdZhhDhqRmT8WETUYh4xyuB2+UJ
vKweR2XSulcJicHb0MJtV16tFqPYvCWNZBWbSS8U1t0aH0xwObGHhOnusowYl9GK
nTrUPOtfau/gVYKJfGrCy9taPAfa0SoJsV1sxC5oBgVLvBJ/MgcOfm9b5/K69PnY
xKRp7Yx5zQIS1xM8AJlunVWdjDQ8gQE4SsAPec5O8kPEZsXuj47Dao9ajSyHbQmh
ncj3JVBURsxXLHqRa5HEU3L7Agq3+/8Q8G2LZHwT+7erfaVTYo/s9HsNj+B1X84i
oPoys9b2DZ42lqz1mnljW5tY5IIitf4cO9tlbbUjfBmbSootOj4UKmQelowXcXw+
lw/+bpDUrPQzBQ1NlYafdP3tjqAgyFiYIEDa/gyeaCbzkVsDAXQuYNZT/0eC+Kpb
HW0iGPSgDeZcOCdmvJzru8lLL6MysfgwR8cGVvGjtq+m/+a13msm8Du4X+2lqhrJ
EVs/sEw9R9c6UqfZ7MVGP5kbPFC37gTWTwPBdp75/Zk6bOz30V7LNku4brirhmzj
E/n0xbUuHjjI9d/mDFbBMa9eBNutixQUNsPUrXcTV/9G1FYTBK4qhUombFBSRdh5
SJpEAEF5xKSLIAbexubAW9CakoCfbjCSjuAbejj/oiLyry4i16n4PwSYzcDGR/6m
PQzWutxcsUtOHNjTlTjNH2cEcA91soQ4QvQPOB28Sy9V8j8QFrgfsfxk2Y49YMa4
Znuvk+8CNoorgbED433Ol5XEMn9jp+zVVljP1WccoDxqkebzE3KKFIkfPb1/jxPS
DSoOmmAwlXChsJzKEDzzBEWmnZcVxcX/xWP1LHccM2qnt1Eqg+hYuMVu3ivomsBQ
6eAeqqgXExs+/XjnphsCVDKGJiCeXuU4dWJW0N/B8QYYozBf88FVpX7YG7TysQTD
Mo1GnR2dTIDeGXAPM3NgflftX/zeHEaxNH2f/fPyX0jnCH/ZKncCOIOGHmDwP1UQ
cv+//jlT5ChdHOWc6KKwkMUUQV+wvLZP7Umd3kZCocebimQRPJ2fXTt4Fn2RqUWt
TX5XbY6Sa24U83cwlWESS3gK2Oh6cuxo4qs41RmtK5SXBvCGihr0Zlue3/Rn/l8W
5TavvIH1vbRNqlL03ldvF8S9pIGM0gJogENrZBA05DHE7nZifiW3X4CNnMhxHSDg
wLeSVLXxjtxg4ZJhq7XsPV2ygyuvBL7IahoMvFlxMwzT+lvRN7yHWfrC9acDdAhY
T/klBGDPirB9QvAj0hoDYCVVYvKA11lH7wzIN9aF4pb3KzOvXh6BxadwXJNrXNfF
fygbpWcuWeW5xELIZ1fb8oRAg4klKZ9gwqdGAmNsdCEE6CHjDJIlGdadTFbuv8jG
jq+znrK5VeaQ5i2T4M96Niic2IVIuT/RGcQjqSoU6gEaCXa1x2oqdv3CFZFtGn9t
5ZKOKwxdMh/AYF4sWZb4FKarULhLYK3LzsRdU18pWYrIpFiZel+kOLNDQm/dgw7l
7qwEbcpm7rj+0PyU/L7ZOr7Jesj+eWT0MiMrUnbrTE6mSN3uP5gWwRxA2vq3nh8r
Bdqk8+ZeJJrUR4Ukyq3DxEy7p6nUvEY/4wJuNhTPPeMLmqbrc9XTGTdI7Ia3yYvQ
7mkpm6iTmrzgI45XFcPmuLr6P9A6YidkEgpQ/D/2TxupEVFlR9tI3rtqI0iiSXvY
bxcJrd5lVZ5BAsKzpPlarIrUaOH69j/aiPaCiy53tztqoFRRtslr8wXzgpHw1jcy
tJJXR0C8AoztsKJk92McE6scm0c+fz1kq3rsbVcTuhQuyO0IcalJ193y8c7o24Fg
xj/H2yvs6gjZoXQeQCuocY/aizwm4y5Y2GqRMax15S/NZCaPszMLxeGxxmydMg5A
lzP0k5BrdR4HdQLWeA3BT0pRZ3k05Ugm67vf/7T5cRMQnIa3w/BR74myrpIRbEiy
N85BMs7Epn0WdwLC6BY4Sa0bprYjWbMXbHZm7RNN2Rw7cecBHTC3vHYF39oNAzr+
c0LCKIfQqimZBZVb2HJ5wHfebi2B417yXhqtHajNTgTfBTFqiTi3+v2/rUcNZFCw
RDhrFiuUifJMLHq2ZrvaZR9UjbLNjpui40N0bMHwmMZPuam+ey0GGVYHEUyOiTR1
XIfBSIuCOuSvT0ayxV0hTGPB11A58JYd0qwPwLRdeIR+BZXvpL5PzGz9wpChqYEh
h4j95HvemyRwMTv45M/JuRPUgYfoNZvTj+lItmh2nJ4Vb97ZJUxvdVaCBxlsfa3e
G8eHpwisJxllYt+JWT/cRhavxcY1kRiW6800FWTn0/JNkYXlFb+zp04x+7b/v82l
qqFadGHtjxC0kMB4pBIctqhxQDbiV+XiyWa6FYwIQm6h1nKr1ftq409M43yRenlU
mnbtK9crywuKsv+rHjQn67vKTaBbySy4nnY8wc5mg5u/ALzAS8fXmt2OrbYXruTD
dizSMmqYJKPkhBkXzGmgeXSVJZWnEOn0PGHGWYzrQtagHr8CrKxXj2UFcxySamMY
+KKJWMQcdsuXZ08ahicyAOZiNThixYc6wLTy6uP2nhB+BbdQorpxG+g3ep5VWEJq
356j//iIHbvnP2DWy1QTZ8YxVGUQp7uxghsvGJ2z9M+cUqnVauh6RReC7NG4EgPA
fFSnMOZBh01iuCAcxpWErxU0XrNoP5+LpjhxiniIZgUIfUMNGkfRLG2xatinaqdZ
yJo/0uWyL7GZEXviqGKjflzrL48CvBR/VV/MK0S9GwBNBMMSKuN1nYjC4j99gtxv
l0W+R74SF5dLZcd+hIFRA1Tlo0IrTTokaXdmdiHS+lbj49XbLvGOWi0OPCWHWVJ6
fOGquZo9Bq7XXu4qdGuhde5V+thl43UfHOywlhTJ2zKuuVof9h573hGUDmZ+Jkrb
xQmgH9dMzVeLPKz6jaM2oIQWEV7nzTnscnHfJ9mZ6o42LxxTl9JpjKByfi6Llqsm
TUBEKhzZ6Qc8BmeMnklAboSCvd8iZQHwSvUJiTXqHlRo5wc3RGvHmlO1IZjS3REV
HK0ADUumyLNbctdY0uKUSIErf0YePhRgIZXwYY1oRl2Y3NA1Tw0inqUHZQdXtRDP
iInmtbU8KI8bh5FCO4mshZeqGwz0Xoj7ljcpoY4T9ukKnRXckfPQCZMBQkXyVkZ0
66Md4udxOnp8FUazO6kNMrlTW0xzNE3CcvB1VFvjAe4LjikhP8yc/mWQCfKgQ+m2
RU3qecFVRBS/tpB/N6lykofntp03xALOFQjEm1iUoaUPCrIEXHpxvAoXVfwUxphC
KU7Ur5hOLWqojBmV2724Kp0V/ZxeHnpVMK78465+ADbw2lEtopVx1FCmKA246B1l
wZ7WAsD1rTWkotmdMlBwhwZuFN5hmVlKu/GfO116yJjhUTh6e7ue5ZatH5CE3Rvp
CcukdEROF5qrHhSK1ZRoV+IcqXMgSDN4A8KsNv4cKOpvInlxCgG3c8bPLODgYojb
s44ADZFnKGZP3lpEAKp3K8N8RwpqHaulTuoFzjNOsKLzAFVHuu9KeJa0FC6OLVnm
18hJJxCxGwwfv7NeMSn7dV91E/n0dxh57SMfD377tGoT95Fm6CStt+1TW8vLdwjY
iKop0N8XJhGCTrYQnqwnX2ovQVyhUTuUWLtZazHrd9oRH5+duAgmUOTRJrbE+ADq
Cdyd3il348al3D0KOIh+oDepM2NCm2RBqGVWe9jGjpM0q6w2IzqFUeVQb2lXF4bK
bT7t3ZzjPHXg9Gpsv46t8tj0XecoRh+THW2kjbHKj8gMR/pigkrOZ7nz7rD68UXm
fhHgK0gTNuui5VaxJ3U5NR1Aoevwv0Be3ihIgN1zYErn5CxDfJsL1szxazSnMY3e
bYPF8q9iITnuIKSR/Q/MmI7D/sZkssY02efBUJNh98flV5/8IzV9noTb6ZF1AgPO
vpZKr+qcd8AGa5r1dFgfmUJkMYxhtTyYXWT9plnfIiFhtLVlLSp3P2F0A7ySIOr/
mWUEYd7SrUZVC1cKudbEP0jA7h5uj7DHgEuqWepNAvIMRbVTr68yqBp23hX3eYhT
ZS+IZPQpr/AmNszQIdpI9fV75OIKWNYiuC8PRCvydQsr4spjy9UBvGOarDN1Wque
9x/EnjiC4m+9mzyO7sLJLQrrfA1yY360AicG163mqTCF5nXNfcsfHaQ49s/vbDiw
vaAEZ2Qm4grZkmw462bTmhrCMd4fiAVsh2mKOrWqlB92yzNuv2X7WFbKGvJh6qz2
zXpMN6jpPxlShA9UHM1i9vW2wDUVeapdFoIeiXBNWPofxG6xZnhIDnzWQFpI2BpA
PL8xBYzAyYaJGt0D6RKHuPyR91rqvM0miQFbila+XuJa/dWvgbpex7MFuRnPm4Qi
/C6uhxCA4RDowN6nSVQ5F/pVzg6VZwfMnfOv0TuKR6No0Hr/KkCtP7QfKj45UIHJ
LobX0OOMKqTFu/OQWd+g3O5YnlFKgfsinAkTNBd+qaYDFxAZ64JFOtlI6bSJ7Rea
Of4UWXJDBnqVLnxGopG+YEw5m/jSNFicn35A1PBOGevrKKsJa0soVz9Ona2V9ius
os7SK6o09z0D2l0qyNOjdWaxHALBCEJUjAg4Uc0LbwHGFO65J6+f8c58eRVQYXHj
0aNskp9fU7VzH7aDH2UkH1Ay94N/JfRUI1sBo9M+gy4NZVr+s71P7i02bpOrDwMB
eh5lY+8ULgmTXqh+aaCPPILln69xCeDji3Wolr9Gp24J+wurTA4+wHrR7wxcaXf0
4BYk9G+KUgFHlE5pDgh3chncs84aq4QySAbE91/n1Lsyti6BJzGCGeYOq5ZH1kgE
BjDU/wHtuQ76RSgVqGcaK5lBFcCY1/vQUSMTsLWcOXbvJwpHFTyd3W2zUL1zpwfq
vGpLLhwjR57M3q17597RcLc2ViI4qh8cDc++G6sBU1wbySk0CIwruf9WaGXfp3Wl
9Mn24K4l+0YZmX2huOjANXEXf1ZG/jynNgHzCdkVoZ2mYJCfrvNeVpFlr9jbx9Y/
Pi57KGd+ijDsuFaiyCqfpglN306Jt1LwB/eGqB1o9KRk1fVAepRc8YXf1DqgJusI
q8Z3oPEGSRUFy76CD9EE0NNJiMUrB7Dg/shLuIxd7GDXeN092RkW5CQuUud7yENO
tKZKwDlHDl8od5lC8OIICY/ujw3yclWSZA2RfR2oku0EyqxJGavuHxNYBeK5i8U/
M70CeicRX45usc6D6qw83+k7hfkxwRDVPiNJ0Nw+VgV2QS0Flq17T4xWWTDIzW8r
htburOsGMriGqSjm5oZkxx5NOn6OnEQEAWMP/kJyC+aAea4xMo4M9Lmgvs7/IBXs
vmvr1jUw3YHTMnvlQcOEhZ2M3hiynatKD00DVlWavMNvMrT2etS2ACPu76J++Iwz
x2RVBSckFzcEaKdEn1s7q7rAmGoHwIeuPV1mb7+yl8hQdtg73MKn9Q0VxRx98RQf
+YPf5Plh5uEIiZQOiLqFhrVY/8FSbWjjZQ84bE+Xv2ggHWzMFa/aN/utnWMQoK+v
lbTsYW/xHgU+j/QzX47sSmVjDw/w/ia5TxKt0AaWpNFXs/NckVY24uTPoXe9Cv7o
Y2CX+iGs0+YNvTQvtKezEJKw3kIVA+my9Hor4aV14Avbz3LR95joZyRXo5epuTE1
aAI8Itdwz0xjv8jk8sVuKENQDUsxatEjamybL/xpAyHikW9UyjgCOcRTxbNiPlYZ
LAEAQA3iNfhkZSRSmyK1UvAsSJSnqekUjNpATCkzBUOEm/L/uTV/FH/3vc/scbGy
y5k+1OXBATcP4U87Lu59PJ4wpyS1Erc6hgWijiXtyN+78NhfjZppqzqJ8no8pY0g
saa75itOQmNleaNnGs4+Mn+EX1X80RTzVTqTI1uCANrrcemrIUGwNIW22AeYt9Bs
686NuVrOtdY7pCYFYygRCuDsdu662BusP2WGkdtJUWHuwJrS/odIAzy4F516C6bi
7ddJirOwJ6wmSMiTPBfEraD5xhAfUcgyS8kRPnqR2Z2/Nx7xfI3cZQKcznwvTs6r
XoYhxqhndsBxI7Dw5cU/K3sD3NQb749oFPi9Xihk4oRzkTQiUFwxqYrg66AewgIy
UKtDrDbNpN8y1Kt+6FHlXfImk0VLoB3++ITrCqcYwyeQBNHi0Q3OLEY57TbnHI8I
Uh8F0kjvud5SuotXnJZGrCukDnNL1eV9Qy2SEwmz0fHcnXSzNSot3Hcvfyj17Sk7
io5MyFTZhf43eZvU8OqoYyDhVgmxv8PHtVxOSr+/6k09lNBW/DYDYXWgJZyE9Rfv
/0eEX91HKFUPVfNNFKv0o+PeTXuR3cu31TDl7JoU7Lr7/SuahxDlsAq5XRIqQk5z
LnFYb0nO9aajLlR7VOBUte8xyBvi34oDS1W/QTgYvrlOMLpNzyNRwAkFOn9i5eze
L8OrR/zj4qFSmrSyGAK9tF0oL3EizgSkrIcxu1bJ+qLttgxNeuD+6sl8F8AfLsLX
my7tk6wLRpp9DdxRMINf22AZ2q+OprL2jKJ+jdFRC0ugxeGp+3IJeEzn1SpgnFJp
nYfamjMHvk4IdrxH8R6PA5E87mB819iPG20Sko5GzYmD1tn622bcuI0Nq0Cj0BFM
U+OyDmSPxXWqB6bp2hVDL5Xd9dknY+uAb2+EGzHz8yf2By0wtKAIeW+fZCmkrQk9
RsKJm/A8ytV1EsLgpYX1qjyVg0o5MBMmQlHCr9YGmrZB/y+yrbvisWbWmgOz7i6Q
XRAgOp8WalPN2IZbk+RvbIFZExaQJ+t849Fc34ruZThYMxdTYUYEVpqu/vTt/I0G
bPCAt3t2wIipKGvO6arKvXNR1R/EolpfCm5kpc2RsWKOUSzl+iFUeKG4N0Tk4cIL
rdzg70NMikG+PvPh3dOUhvoe22pM+8zphwds8YgOvNpAkN560K8xL18i1r6ACS89
NXH1V1vi8CQiNyRrHFivR3UVtXv4Rl7GwOje+KGsS8QP9Y//82GGBeHvrS/jPAPY
ugj9X3NdQn0HjfzTwO6pQwOWhpaXysbh/6S4Q5CyOM+23zYiWISscjfaj5VSednS
SAEf7w0WtYH/uKx5sqTBUkwfKOKESGDbaPolpG94bbKuZ6ac3Awfez9mI0x6yAqG
ly3QR7ePZWN+m2/0ucej46AgMU8AIukXxQT1SxvZSi4JjqHuzbLtNIdhrcP47xVC
nExKtZfPW8NfGIfrZIOxpgWNqA9fw7geEIHittx7p/ybK9ugJqIZBv9idyDxOtKx
s+HjsEVB69Lw792l09DcdlDfTWtNywZwt4Bf+ilLd1tH97H/xQurWzXXyOTZsskQ
hkDYlpNo63fM3fH2bS2/W1QZGxkB4zTuY6qk3L3+2sk5y+i3/h+YMlp//IdsXpVO
NkkvNq03H1iPfiJSQwmAMY14LTkHJ64Jlvw6krfris5iG+CE3BYwiJiVr8WKzDZw
sXDemS7brmEn3anlU8NH5ZT21f0t7RzxPNgdQb1uTRkruggtzbxz9+YTFUaE+diw
l/tdUeBjLTprTKHsmGicyfvt/WcXZmAmyyIIQUq3xLm4RpqMxCaVdDgJZCC3lcPw
EZiauoCPmZoF+K94xrdtj6trdvUisRb6lRe4v3taU0lFOaz2O+6rxBgY9+3+nfT7
3FPzL4co/o0pioz3qySkfkJACzIfY9Ib7KSVPv2fCqSrW+uBk+Sn57uRdYCWI7RB
X3ZrO7IqfKc7DEvKo3NBp777cRf+iGeoFjVx4p+9opZhtmAIhIfs9qTzWaboPnku
duHzBmuhxKNL2S6i3ifWIUVg8bN6bmgcoJ4PZ/jrMV7Hr+8Kh8RCtYIQ2RG47hgc
oT352jEEPCnNSbfX9MA9tbHMQ2EpxwxjnkIQ2GszEBEZNKdGuocad4A7jPECmkak
ACeaxHVsVLZj3MZfU5Kr73sUZagKaxVpY/1H6GpNCKBVKF+p9tWoukJ8XkpJu7fr
dS3ehOtEm7S3JhdHIaMZCBfpSVwA3qXWGCUSf4bujLkJYRSpfWW86OARDmhDk83K
+8/S5uemLAaRoAg4R9VDJ5/vipu2Ywt7bnZ7oYRUiuShZrmoGutE9jqfGtcUnCIk
HoFMnwzwkDaOVnJqvT51lgHsgaXanvwJkH1FoMdfe9Td7f5RdZb2VZboty7xiDK/
sQzBO7iphZ3IOci+oH5sOBt+imuUc/p8GGmXTTIxggyIJHgAl8iqKinWbMlPbK8S
ExnZ04LzccfNlW6LfInkKWDmo13cIRmXrv1EJjizZFBs4j3qZKv+1zX0AomT98N8
kzw9kCNLeNJE1oYwsfSETftE3ktvKSGIKEZtXgftn2MgL32tfuv+bsEZU5IWpNbS
a/f1NIt69glJUuFWhB2FoGychnKfKdRb+aNZmmBDtnaCVk+j/skV9pEJ+luGAaCB
`protect end_protected