`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQbJEbp6Y2LeWNjLkF1rdiIel7RxXHfKEuCDYOSRALY8i
t+t1uW1K9kECgNZiVRHBc20XPUeJXHhK/LxviEQZ9igLb8QHp9jfGEZKPZYguJqu
JL5AHWa0B5wVwqlHSAUNlVGvGRAcsM9NptTWev8gM7Fdwm8mlnZV1KglRtwsyut7
C+/g37/1iiAawmpooYGeJwqUkgAGMurLeeFWFDF6ld09XL19pZBg6F3iL9/L3qyA
4RqFtVsjMiiN7JXzt07N0fnhxqxhuxEYnByQaSwMxwEwa/SApIQGm6pKbqVGNlv/
oFjyQi0I90p8nUITPByfVA2GTSU4gfFr/s+JJld/DHr3v2ot1Q1kMRg57yQDaour
VfiTOugx95bIm7RzQqaIniz6UPUVmXn7rsogzIRoF3a5xxGBkQ+jXV7vUWp+FTYJ
H2wvq1YpqWbvxazuNmGRwqcLFN1sV/rU6znsVptdDChOWJ0pYNIE31OGnchfL+IL
LyqT86qa8/bVH8cLcXiFrAy5tNjr/S7UAZBHVbW0KFtD3Ws8Igg/JMEnpPcdHfpN
nYljag9fhc6QR0njYLxt7zX68yeFFYdezuMx2LSswLTHkz5DqbLMuQyvGpZfb/Of
uI8Lbc1sB6cJI3K8OgJOg1cGX4KO6i9Iw5rn1sf8Qnc6ojEfINzIWOLihKuDH0n1
Pdy9im3vBmip+4gImD74jY4zHKA5Sw6C9f1qfv32vEbLlzefLtCCMBqNOXYay65x
Bm9+CekcuUgMSpiOh7Yz7vu4VKC3rjAbChXlOvqOltII7IGW7ueRGTehZ6ZR+1jv
FBrj/o6aou9x5ikoymXYNoSFasHzfL4s4ja+mTnE5ff13xe9FC/Xaif8F7pkiAK8
c6432a5OEoeaekUuBTFeTP5S7mTvH+tWHBttLCU6XhoUnXu56hs2ywW6Zh2Cl/8A
oDnbpJfKuJdvr3+p5FGshW1nu4/n/vYk+TkEJDp/sDShJXUM2OtC36AncXq34yhA
eV52Q9oKpH1VFn0jHnkKYnFctcRsub7jJ/ebpa/rTx6cf4IhHOG+NnprxIR+ZAKG
0YTRCGrSa85BF7WsVxVBwXsEndSEyKnQZwdLLdHDoXFK7jceACKKM8LtbB0Jc5Rt
39GHOz5txgScdnwHEGFhrF5PeFmdCHtbOr7LfWq0vLRkdaJEVYiTRqBYXuFTMFHQ
e2oFIh0rIz+S0Bq1RskCFF1EDtZLexOTxRF/iiS8uAYUzcfzUOYPb3iK1AznvYWh
D5vmF2woABepRF8c5LP7mJ6pxhodQ9tuzCFfPPgbLnPcE6/RV/EhVAFBsyBMhi1b
Yz0WfW9tNj3llVRRM2Mjm1HAiL6Gmpy6IPKHrLe287WIAq8dgjFS3NPHTvMFz1qm
FXmEY2ouMYX5K0SPWwM4sz3Rncy/loy7fzif8//xDViWB1fEqx2qlOgHgESMaVxt
DYHl/3XsibK2cOPzg4wXErp/gzwdxysAOKR7f2vrbsSeFaQfJbvCozc5BH7QFLhp
XhI7OY0cN9O1esvbLwVWne41GppF4EoVNG4MiyWxm5qpNMYokFv+QJk6IvjQX/7U
Y6ASadk5K+tLeMfWQfOZsF8rMSu1e+KMxkoH+hUytt5SiTdolPDes+jG7qgOTEDw
PtXJIVCXJA1GbY5x9HalC+oMxt2DkRjihmm2v4/OfrwLgnMX/+hQC1uWY+8lRHJX
iJqGIJHf5kW5d73KX66+kCmjqvLQT8rv88BMxApJYcv69xjATC+obPdxUjkuTBq6
VGSYjA4jZAFRlAZ8z6rsyMUG82RefxVZ/dP7sMZa5vU8W1M8Tf28pNripkK32WI0
w4NWHEjatt78ojTRLMmBTwXD7rl6/v64zUULKVQ7OjVbVSPPBmiuC7a5qsT1Yi5t
DKW/gQojankb+7X+3EUGQx958M6/CqXd9X6vCJOzMycEt+ikPk3OPx6VwwojpG/L
ilfFDami1AXGUix9SAS6cruYuTuE4Bcbmi/edQgTGI2YXsP5TUdJ/+t7sdwopCCx
o4DEub0LUKblowZLX6/BsRlTs/pTa1YnU9cRryIpc4Hp+lOWbldixAGCX7LS3eZZ
d6h/biMucsV2BFxBNwsi17PaQ5P1BZWPRckYJqLhxNR2TORp4RgjsVoNf3LveHoV
mx2rI6Iwgz1ZLzdClsp7LaKfFOdpDz/arDP5qG6lKEUD7ncZY1gDm/ZpTjVSlpGd
HGsIHkuwb+grNvFjrKLmYDy+Iu09fSrqwu1sJQrmjGmbzYadHWbuckihVUrZplsB
8jZ/tc6wdaTGnqUVEWRqud2VsVtZOqpDzaPsS/1g8DuzT2jayl2k5B5ctU866TB3
n/Rj9rcJrJT/PDln87e960GLHGCUpu68nlSzY+hsY5LLkUeE/FFF6fCxuU2sPFkx
C733R5KA6BRzOnRn1bfuG8dvuoTWwAVaKkjljNOymEHhxbTcrux1Om3gpClnX+T7
q7Jh/jYXvTLB8nYontoJfg0Buj3suqD6rmulmdYIoOjpBsdTivjXttt+r6GYrphb
nVIlDI9FT1bMuAb74/acZDbRtVRZk0QiobIP6oPOYFn4jrltYg0v8ZgW8ESCA41B
Xy8dsynez+Q3VYCX+ePxSbk8znUylcFjDgoaVoIh5xvQl13Sfe6cPzTBjY7QKCJ0
EsT1idy0hJPFZlwUK7iFqiHqwDGWQ5LuHj3Xr7pffIoufqAUvZiU8x3833ngvRoL
kY58lRrUQlUThaId+5kgxfNuwYAOmA8DOKJ/+QOfjM55Kky3QvS5nkTqleUVV5GY
539sQ8HBCNeYpFSFHLW1wTujB5PK4pMKY/qRhitMsnJODHPqd1DBHGH/zpgrK1qK
6Q7wNlBvSw4305nytMEZePHos0FfWK/A2lfXyIbd8CD8yQPIFkhmiNzbhKTRikG6
rXGSsyesnaNscgqNPHloowzoO0FZRotR5NwH/8GYVyOgmI0l93FBIlpNOjIxabfI
KbSSL7GC4GwG+lpFAqag43aRsJ//leLcY1kzv01GsXnWdfDbxnC597QAGz6SG6tN
y8idSAhTjAmX1AgWmWCqR0MzICrf53z3t3TA6Bmd4TFucNC3ssSnswntYZekfBX8
J24ICKdRYKWumonqEODJX0ZNzTzb7XCeF1Djg+KbGlM/yQvxe7RjTR26uno6kZ/H
Wu4A648mVxRn+OmAwX60TgXK2e5lMsUadNV7aqdrhFHaKR2lPyxRAXPycovkVap6
s5S7abZJo6jXQy/ysqw+O07Xxjd+4ro5NT2KafpdARfiX5diF12qXgtD3bPv/+jk
iHxvJl0evJyMKg5wQgcKMEA+kXheEMNIn4ghHjOhQHgde0sNd3kr8myjKtxiFzWC
NzudKXIqZN0sDDGoHof5MBwNI+pxIWbDCbuY34fN/iTxoqiko5cot5VsulcsWzXt
MfhVBqJq3IfvdfifJDVcFqMYzs1wzNui+oyjUw51cLN20WCYok+trEsgS/qMTJ3Y
sv4ue37jwB215mSMktIdXh1uzMw2OxId8hcsge7qxihpUoK0+4ZhQTH5328le8Pc
suYRHp9to3WFrM9uCMgFeOnLM0OPsxTuOSxEyVx0wVaNyonQP8xdVlgIyTiBATkh
mfLknuRTmNZHxGt17MeOO6Kt8DXP0sq6HO8FvhNPaME9uj2KjJTsQUVkq5lgKbex
3MRNot1KxBDC7D+3USyYUo34dxvgiWbLYZ/4t9dyVzfapc7q3lKmup23ikRkteIa
8+mzvUe5kp/iCl86nZhgA23jKP4aPYQQ3BuhKyMU5qEZFbdONO1Nb8VHdaKeHXVj
arszmxzvaz/FJAyGa/q9hVbJ0ib6vVkCeWykK9UXRjy6by1RGlrtie8E4N9wq5Vf
WgcnZCdbmz/Yqbk+++mIlaurQqU01xWzlAdkJJAD7j/tB30qHokx5piGbxjGuIsp
WvsIunp0opew+y+vk51b51R3rvRlluv3oVE+L/Iwf/1bEe7RFbx4LWAscnd3gjGk
hfS4uxhULe1SpT9D5+4czG7KXD4qpxujg6QGGdupmc0ziaTmqE2OHnctLMMHfZ7H
jqcFul2FlBLxz5wQqxdDpSYgOtlfcuLLVh0qDmvC3mmZgy/zAgjLvXx3QE67u5xZ
PmhsXVbCSUBuueDgO8Jm/EEYJPtDEp7y8+D2T5Pj2Z/rahL3KmQDYyl9pUgA9YmN
v80sC1Ssyd0eqArzYaUgk1wxWqgwZ1Kht3S+aSoQZKpBj/SVG3YVO95YV679KRkd
7KY2ZfF4CNWvWRi4RV6vN72+wCQNEsbjmWQUA0Xlj4NbiTNco9bTRYp4kPToYYS9
IcvBrF4hjjGOkfK76JvlxLS4baMlPHCx6oTsKkCuS/jug5ki5Wmyhs75GRcmCHuh
MiVzkA0KMuNTr10r+fFGwDrNsKsjCd+4/LZTbWq/1W0Fl8FCY01HJ0qQzqP9zwxp
BG4N9niemk3ruktDl7mQFG5m3ea77A2d73NyC4l1u66mLobgNq3pwvTDDMHhKIk0
M3nFT6ES6LuIxs2Pf3v8loFRTF+1hm8iZk8+obwTad7QYZeS3ZwJ7jOIfzo4p2ts
N8JGdH6uhKsRI5S41nMN2/kw8wH8Bo+D7Sp0Xcia/k2OVY359vu2YrWP93GUWHNT
VH2fTvNiu00CoBFCbttEWNND/c5FGa+9FqT9fz+yDEDDKDOmi8iREeFpqeUPfC5d
+JvckPJ4FOZK9IjACsUIwHfyempKTB7n9lwuKQqlAGhnzIN8dQht+xRzeCtnCUPw
nSus3AXAN6E7Ieiqf5uaAfKdMZgnpDObJ+CY6G/+C9kJ7w7mpgrAaQ5cIzVdcATC
L0++qRTyNwIDCi9QKPADOFUCVpoQPoHE+UlaLg6BEbwEm9kc4F8YpwgNLgsQNodA
+7/+ZUeT1UUlzLCGAXtQMtN3qQsu1Git4ne/lLsMhwxpNU497iG0LC+c1WE32ftz
8tcV0u7LIryPfj3kA6kMT3ZAM5N07JznSjd306bf6+xPf7AKoNU+PZ8S8uRxUQ1T
wTOaQ1inpsNhdtSLR9qCPbNvdcWEX+ykVo0fv82EWwlEIvBPDMGNdJJAWRRRny89
0k2KYdVmWmxk2Q7HzfPz85WGeGAnFhc4df3Ya9oPPbhlLNeyUMu4cAhGGy3WsxmC
klxMA8hXLGqgur+yfp6dhEd1xp7LBtU1vmefezmIL2bs6fOUjGdWWxv6p7QG8Qns
GZMtFPj3Q/UpDLk0maYRTIipLEJT/ZaIVelvqJN3niof2nAMhO1qrzQdd3cLqebY
umKXDc9iByvSRqupa+gTg0JZw1GO0x/iMKKe7utfg3oe6Xt3d5Al27sdRrqBN2El
5N12+OPpAY7TOF73joushd3LiQYVml6jPnCbrJOCg6OCue/VceNqfW5n8DHm7b3l
pwFmR2Szb3io3khskquFXXRB0dipVvGuMZpsSu8DSebFv0iElIW/UisE7xywGnCy
ylWC7WMpICd2LXdbuGzcOLIX0mow+YHxdzYcPklF63n3bMnbVwVKItvCJ0Xl+kJe
Lrw8sCa4dulNaaizu70nmC7Oxom6JtIMQofbnCL9CWcgGSeuthj3UL+KbxB+kuJH
OYM9mCTzrWRJvRb5Ga44B+f8d/zK/8QlyQ+bHfPtHS85NtQDeEIXmPICozbmQ+pH
WrJsNyq+WpkotZjQMD2kzxLsYEx7bRroJ8CsG71xqIkVZ+sdd/DbkgpdOe2bqA1v
129FVdV65DiYMWFbq+rF6xr2xsAT0OZqhquzCu+P0Mva1ZpOEKtpuX94cTDpUMyZ
zp+bBQFxuOfoerw1wvbBluS7euilnSFN5QsLCgYMPikKQyBQCvyiAWVozDX4TjMY
XlJZOF8f4jvg03GwJT6yQqiB0XdReoPwpV3GGR2bC0VovzSg9CYR6fmV7P+tN29C
x6OmFDouXxiMbtFQBIU9zfZ1v16s9F5+uvHsJF0eB0aKzb2natIspB4piDCtSjAk
rh70E6ShgfJu2kruhpWQyArBevursqso4sQUykhX0tO8qkyS/DWgHccwChp9kQfa
68BNKVfNDhrHgPqpg300adR8UepNACrLeTOm95uSzEKb9NJ3RU0oVorDqcu3TCBT
h2nIIyH6Sc9K8B94g5Shb0zZFVvhqxk7JSnyQBCudtLwf2S53HVg0/BGBmvEdotj
zlekbavcM3qOIR0RSG3PiHjVecH/LrmAgUplhz+fnEAOkwA90rbBpEz0XBPbDDrG
aoU5QluDakfbSaCZ6GP6dCpy7gO8VE1jkereFxjIr70Yqxj8hrjolleXYiXtHFpt
mod8u0+6Ik+kuQChYknoWSAE7dgNWe6rtDtKkP35Ih8VqEWCHoW3SWyprB6+EDdx
fix4n0TXgHYf2JTQ2/aYjYGTGUn88naPQfoe9oYvI9gPLN3VbSGFc2O8W+twWcr6
10V0R91qwW3UytoInoL7CBocR30vC6pLqJOal5mRQ86uQUo0UeqJkwgkYJ0mTp21
7yBvlhmpUyE7lgFAzpZTAY4Gc3KGbAuNQu2UP9ldyug9j2I3GXvj5hc0bsmUxUaK
izwtkdUV9JMOpOF/hGfbATintI1kO25FVIeryDXOj5eu1lCGlCXXCVKzg5LH7BAK
0dLxzVJ7CnCvM5Pr2aR7URhiWFsSMbyiWMFXUdQn9D9v8Wzv5AnaCqa0RW8ikch7
4wE+GcbOKKo/BQrd+MN4HRuNQBdJq4MDfMVfr7UtQGlXLZyqzMTcAh1vbq16ksJ3
bd0L/zCCNU3kUzPoVP0DrNmiu4bcHaW53tZkblxGHLvMa9NIWniLv/3SXRyYfdvI
JCgblg1KCNF600ggSxxBwGXk6E83LibgaTCWlYM//5iwJekeOpy7MGahdlUGIMBD
8BNpU4WUyO5f5b0D8hBRUVkTrPmxbQoL9NhwjoR3hXAMimhXUDmLBEOswHoQDgR9
tj1qTR8ySBXS6t3B+GTTJBohucHdVUgNLDCx3f2Lgl54XraBisqc6TNXKvUpswyr
NDGxXDT4/LcrIpYX9R6X+wvlQ2ZJn4M3YAmro+uTxbvAKM35gpd7JOAYapYNjv/c
NK5s39uEsT69gaanTTUxCtg+51FwxTX/KkiAFQTSnGI5vDaSX7Qhk8LQBK0xuiPv
UlyPOIF453xdG4ITyREXKChlEZKYpgGygmeN/ZNB8A981GEXgTPC3/MeX51d7k5F
H+5d70Wiz6bApYI24c+Ya99uuug4E3eysMAeaO8zkjlAQVVwFJE7sub+Dp8KIcrh
IOSGvcUwm+2jeFis+TOjJjjxCE4HPZJ5YAXBswtrM04KanPaX7ggKElLCtHyoQbE
MOEVFbSUPWMp0xduVACFeOlXpcyIVNVDsweg5ioTiDyXZxf/VRkLrxrs3Z7w2kvc
eIQdV15LFYakKZNqIwfmzAuD84zsBpcywIdUatvww38p9+K40/u+uoZMwYq5vWcz
W2a2wPHS2Ajn7UPRw2wEtA9SA2nI7dIVFbA1bRcp+CdfJnKrMaQP3HLHiMgs+S9T
R7B8y2V5nCm472D5Lj+wFju2VUbOyQUdMT+s78d1X/2QmvI+6EySsLnHvysDa/Nr
FxHTQ6M9V2IJ6FPGBpVsIUlhJ8UatcMzXqHrhX3K2OLE3G8aPyagMH8m7NLkqO1Y
8RFeKU6oWaPR/9ZT+Nf1hFor1S0QlzFQgB6mx4jb9HisuV0pg3COYP8Tdu0UMcj0
oiIVM7PGbQQptqaimQY/WSmPA9IZwKzRPJMqNunwpPdzFRgA0NzVrZjpD8mq8bh0
zqBsuCmmg1vMeVA1YTxDnDFcmLWjQ1iTAX/wcgMvjtDcEhrv2FoD5RI1Jm0+jWp6
voucQBxOnKa+QyS0XlQamyVA+9wSRPdGinluGadgVchpt0Pl7U0thqcW3TWAufZo
YBXM7UNWzfXYS1PdvHzFqeWkKsUzbR55NE84yGBgP+lkP+ISCINVtIl0Obvtzt00
naYbSYghydM10q7w2JuZqfagTp2L13SwDWiKR/QR0X+zIQgR0rVnfo/dNFDb1NZE
+yqqc7M1RpdnccwshIxVOScmjManUrVRayOCZmygpO6AYBAU/Qbc2BhJSYSBU0U1
zn2mTACT7OzIU1W7FSbogn+rtt3sbmsAkANjaePAekoRUvJPCU6y8f6OC8gA7hbN
7l5RxFUXKMhcieCE8FSrFir+kBK2ePSJgb2p+aEDadpqg+uD2HrR720YUmOweGeS
UjEzzEJLNq8drCAKdmSg5wlnHyLUP9QScoRRpicGtw4h40oOyErpooGrT+Kv4IUe
jFAm79qJvou8Phj9JzH/Q37rCvqOOl2nqEUREpgUXi7uGnDGVFS7qz49FKeTQTgw
mgDxYB2E1RgQ/MMLQj1YVLO+c9AHb7n1dZtaoq+GqLLbN0X0l6SrKLyauvQdLCYZ
Sg+oP4zg7QEBsACr5dWo0DPd8eDt8nJgQmugLpzJ+gGh0p/6OGWAPPVGWOAHwsCX
MBXcQI34m6xQyqNr7gzgq4Oq7+SYFzYizRyheeIJLJZ9VNQQ9Zmk/6R6txl7YxvC
ii/JEj+LfgR2DqFp72tEZQyBTlyCJ00dGhENFqukOrQBh9W6TYDji0dJ4rM79vmz
7wy2WbMZLF6OQ1TrSuDZtZj8O3MvMUL0lMIU4Q4i+J5x/BYmsTjGI77PjJX5I2Jc
Y2YHh6AK/cMsHW+fNxYmC7xjmkOQui+Wn0mW9cdswiqOpvU+PB/tr1RDy1krUZox
WFfsRZD6ZCmtDlZZtEW00XTzwKPfSxuyed+NN0Y1WzPWEWIdXEaVYMj/zkL/t6am
pKnrKgjBzyAcYk5cQe8typO9irxRO1zEie0+km6AY7/bCNRqrHrmpvdjAdIu8ZPZ
OSuMJw8Vpgd3WeIoItQnjarJzxl/pJkQ46lXoX/BpLbMeexkLBKD9tR3ctOq7O+8
mXUnU8K46GUZ988tkB68ZzBhYPVCgKjfcq7TJ82WatDsv6mjHyRGdtgQ51m8f21b
x1zzsnnZUhblEtE38IhpV2a+7LlIbhBNP3q1Jtkot4Af8Pe7FOOyLPfRjVb8AUUg
S7kEWWr0lqEyNowpTN42HqX0RyR9kT6Q3QqbLKbUPG2pX6+RRf9UUgGTfBLXsu9C
Xo/AiiuuOZvA5G7osTBJwPrdaji3dvJTsvYP9AyiPcZduXc3iWh1KII0rPGaD9nD
kWY6+F4G/AQm1PDPmO6VcCMtXrymnpM9M9Mx4Z/XGd5whCA0JJfdxOPxLWPTqb6K
9XHhmQdNjqEZTv+nULvfGHVL4UlGctk4TT7YyI5J7s35On4NFp67tECatohaMINL
0PLZ1vGnW9R7534JHG9XMlKaf8+qCGRabHy6Ej8DCbsB8AVu7qFnUs2EhdVepAlY
pgTeNKeKUsZPe4XDWprJ+3pmgHeX+CUIYYBiVuRsHTyU9Wq2MyFNiD/SIoezL6ds
7h0RZIxPIazUzQYhyQgDNZqYHYd0fazQnxWaAcUovFXuaEyNpOL4Yo7MTuKIO0io
9BvxH1t1dNHUGVdNv0GFzET5nZddxp8o2la2s3MdHx4d004dBkBYxN9rrRT5ulX6
GdhUgKXXliies4Jfw6WsSFgMqqrKb8dc1YXO2BlOxLGNXB4A6ztOjDmie5GE3VMq
ZJO7o03v7DEfWKou/yF8wQbgXSAzYRbToZ4nq5Ilg21ygAlpTsCRvO+J3zRqbr3Y
CiSf3SJwoLmJ6NQ6qTOpqE/qmtLhlCUML9oay6JbI6WwldOVjvw1DfUzKllD4q4m
IQ0mxQht9hqCwU27SLSf/p2nnVkffBrt59A+CoX0CmB7+vq2njKrgt+nsINmHuPG
F6CYJfXr0064kWchA52yV0kDLj5HLeFJsutpqmHvAFaGWbzs2q02jGVk7gPfLYur
TeJvznSAnVmWTZdGaTnPl3MNISt45oPy2/7pxY8h47HRf+eRt1yAilNhxE2nE+5G
rH18q9cQgkwt/2+9Z/ILoiQTM8CY+m28bkMjPxdLdLl+E9mzPN7clQCIYNqK5SfR
RzYkIr61bKZQQyyQK7tpZZhzCuz2+A3j5g4qpONCcXwpt5GgcGZAqyaNbSvCKNgG
5lNVV/4nRv4hOKCBq84iY/0kzEBGm9k4FsE3oOXHYnVEbG8vXJOyn+qoCXiE8GB6
fjaA6SsMWus8vd0sU0jmRy5fXfmohXJMebvFQMdX7F11Rgr5gZkMwaxO50M0I9MX
L5ZaS4ttsOvJf5Y0W2eWK5igSGFRophnPy0FxOaKe/Eatv+1Ry07M2O/KP7Qulc5
rQus0AqzOVniPs4SC9Vq+jb7ZUOWjHHixuKWeWoF19gcxvO2IshAqOjtRcuAuHCX
5O0M/ElSP9P3gd3eLzugEGDaqS3M6ZpCd4O2IE4xwbdFN6qzx30KUkk9ROL1RNxl
Q66/QTepG9Eae4AmveS7nO5PVW29k8TWIhVgH9npHtft68V32+LkqV4kZp1VGoRS
7vqG3+Ai06YRKh9py8J+jbEt/Jj+Q3ygFl937lsHBlUU5Q7QaZJ0rR7m/+vZvZmT
lXWnkWCaFkEb9kDKf88WcRnQBgny6zqUEP1mgLyBLQCPFcG/k9eBSi1sbYbfwF/Z
B7xONqlX5TjdlMuud6u5Nw8ZaLFcxKdmYIEklXRqhT0QQI0uEuNKrDFnsqv1WIYG
+dXOEoRvxgqOuBaaGu39nATH5CnYSbbRjVL2I2izQ9iFdikQkkmAp6VNHMruE4iA
zwil7N0bvSoIfLGKUvoYQ4FvneetEWt26IGEspUCD5OC1zJqEoyx07DKQ25KOkxl
FH7u906vXZl9mWrzt1epi6P7MweQRGgg3FW6RlMSHViJa/zn3KZ73aMDqz/X8KnT
woWNa6BVrXmV6PZ67uTW2YXMqs0bwa6wSjdSPWzYEd+MMIqdNjMb2aUw5FLu0p9t
iS6aTib67l+G+RDbf/WIl+JFhaE6oHhmj9/h7/m8xrXpV40yja0C5XXfuPWbrTQ/
YmvyBp1ca9QkZu4ncfcMZEqpEDJ+OljCWCwqs5J08QGCxsDTKbBFPNhP6DSNMB+/
sWzxCrAORB1h7SpeXg2MLeBRqYSWWr/GnN9UJGkcAUiQpusJZx8ARg7atLAMEQKH
GKdGPtJOr5HbByO7Ty3RGvtltGd4P8c5Z8uzize6pdBsS2fgOTBJvnARDBSBAOjn
NPQ5HM2kuEAn/+Iswugu0LfvidT5u4tHMwsdiasOOhZGdf4EDxPpobKOwLKa4iMx
mh4PZr5pBPajmbEgGmHAg/1G/2lip0ng+ioDeQf9mCTnpEKlU5RhPV3w2rnkTZLw
u/LvEs4tPzJouDskrbhyYl8cP6lN/L4U/1qTeKFnZEqp0K9bkIR1/5NaQAJQhM7t
gH0+9qg/+HPhtryK+qJv9X1tey66jxe62JNxM7XdOa/B633YTkSi0cj4d6POjpg+
VB9Iir3i+K3dvjLZmIezPZfNl756FPcuX/fpUHdEnNu31nfnRGx6uw2QoHM28Zl7
DjXKHvd9LCY9DzZHZGGVAKRiBR03gURJuBVFcHAtUpqKjj8lMAUv9O6hQEjz1lp8
MzLHbGrRq29BfkSjq/uiYZjz/4fSapn8Hrs6Rpgnd3nStzHU+kaLh5TgEkWjXfAG
glYz8HfeB5PAPJHmyJ/6FWAWRzO0cJulKh0bd7AqnOvuw5Wo+aaiJuM6Uabz4Wmh
o0xwuyh7kdHp+nKHuANI6lugGyUOCP8smrOaLVsfIAuz/+U7dinh10uUZ4gIoTzi
TtJuuYa15Q0Wd1CR0hX4ic5a8CxCcJMsO5Tz4va0GVNnOelt97IoA9nqukkrgacg
cjgDTmr6++opHXFyIjyNpPZEy/be18oS+fjb0Nk1nppr8mGLX+MIahXOPNpbekJ/
rKs14I96rgESk9Ed0UXwqX218H7id/iMLjxcTg9P9e4TdYodZliPualv7b/OEW5O
2u5JDDjd8bTs6kvHclo/x4qR+VeClKCBIwDx7DD/nzKVUqtdePieujkxmNcnBuLT
82dU82UbmjJ2EI6ixoR23ZgVqP7P9KaBt60vjTJMxXhptZDcL1k2mwAjt3dY0CnO
5yM/bU037oZWGgig8Z+WcRia9Ieq/twEk6sTvoMgq2ZJWB/2/zNwgqrrk6o8KEVG
2nbXW4/fxHN+VdUAl4qp/0At5dcsHbK936Ok6TIVzkgp7Hzmcw94pa263kY3h2rO
ZIFwmVTYwg5+LGf9JZTERY1Q/pPiLI8zGgbTbWx6U/rMZGnbDc4z6DNpgSLCFbIA
L/gr5xR/Stba5SZeW+3Xb6+GdZbhzJL4q4EvY2tkhl0gDYTa8BrU2dJDzZkbF6dq
tGi4xhjJmjwHuePWJR/qqSXxL98lQrVquIudzYBzd5YP2fRkFs9UCogTFdYPuhs0
89crBPXWmPIfbYMEJrD74TE212pLbyPcGxzZmj+Oa7JtoyBoKfzZR6GCVNuGTygc
xtCk4zDinDHTwc2BkZWN6YxFyuE6/+dB4hbTP/l37gB+QogtjdT4C7zll13Rr1Jx
b8+DdtuNkjy2YxtGs7UueWnrg87bPilmh9FJKKu4J/xZ+oFL4FPj88IToMgFd+2V
KaHpuXJgOPKPbAWdxZ68ZAnXyGOkLzKWMWdlbYnKUdZGJRaXUjp3t49KunEenlXz
NJZF9bec/EJSNlxvvJVpanI+gyjZbANKOI2rwVkNcpXij8OTzL7lJZBSaMSV9miS
KUegTNk042zX12gCLMku0RMEX7ntz16IeW/IVdW9y+wSn9Nhu+PSqyZlHb2JJ+4u
tXyp2Hgkd8RKnYR2i5EkPKHVJ6AZnovDFsyMsXpjVTlUaLoyUft2CzcKrd6Y65PY
fp6t58Lf7ASvalkt9RJE2MTupGoofEWboiaiKpDswYYVytkmaZ8Vq8HPZesuXRn1
YH5R20hoOlLXR+dATvMSpdJpvsv/IN4vPRbuh1ySLfdmFm06J7dZxwoYFEKYQtwD
rTuGiO2u6ifZFSqFba+NEztBKBnHhLTp3deNJAE4GcCTsVtR8XIicyHSZb00HpsO
vIal+VskCC+vDMR95wPCIH2B4YdrhCbP4HKHXRD2WjEO5vXB5QAOMNTcWGiegDTH
g0UDqNVSAuUdhUZlrgy5Mtxv526VkmWoxF3T4cwE6q6Tu6PA7uWak8oxG/CyD6OZ
eLppGvkmNn44+A2yfpkMlIh4t6/cj8VWFjhPDRluRkXdEkNIzZr9FE4DwMKIj5wc
LH4cCTLMgJuSkLCXZssY3gCNbVtm0nsVvq6fHRgQyfgVHpPAHJDIetmEtXbCCW7V
tbBMJhbMP1Pi5X+tzcPwfr5eLYbfHy9lgBaHiwp6vCnwyuENGCGq24tNF0IzCJf1
7ZJuvA7zg4MJ50zLrWjP9JO5ks8JHNWwAUd3/S6ne3DuOAuFl4piRkXx9XHfBkOi
pC5hzFwitj5ewl92E76FWiwbyK1Z5sqNtDjFLtbrhJpnXuGSJ3qgI0o6tQ2VzgBY
u4/YJ6YAS0cj4dH09IT/wHblHlFfpodOTzdhpeAGW/AFZ9zy7UhqVXE4sB1x1AGU
eqW6KTExaXE5GJsGT2mmn2ftSIUs3F8gjnu2vXmM0Nn1bkdk8LakLmN12zicT+IS
EXOk5s7uBVWuYiO7Hs83NyGhruG2Hu3r34m6gl2QLeHDBNBtTkgxHht67cEZTXuq
3UpXI7YttOTqvWD4WlzwLXgD8aaqHuBVnCVjBugkj3W8GV49BAtDqcbQjpNiDBFB
wO0M7L00oBmYv4vG5MZ3rSHfQWZ78HiHtTrXUsO45qQkKug713BrcJs41fJuXGAN
wXPUL6Twu27Ef36AkygEwIYFyPGJg5owU0zXEF3QdGUZJLuvUKdpG5WuGqJTX5H6
l+TfIHzT8oAAenbnQCb0wj2SKNGUeuGcTZ2adSk6QxqM0ITXmgXb/WJRW+sGbrSA
15qLTr+Kd+BfGcd7++vWcyO4hdDkfAntTCz9uA4rFozZ+YM60Or+MT3Gc9v+/EUi
mK6OGJfW+Ijy9glJTbl0eHGq4+YVeEoDJIfHNxxrDWpiEk7jizrESEZr39uWI/+S
1BDokVScMG4DhbJ6YQDt8VSOoG4SX1SVO/DlZp3s8WPXekhZaNbqN5AgOocmH09U
X0svoJD60RDrGlevGuuSPpin/L98yRtop0jSdotx9s8YaubqjudZEhVKO2t7hUWc
GRcQi0428Jn66j/iFf9J1ULyKa9Xq6pnHiUZ4t+tl/+pIzJ2nFwcAr+FPFVjplOQ
CbEIl0e3uqZlLXj5Iice07CRepvrrLz/gjUqaPuxWetAyYnUrrxqtQ32H6sC3k1S
LqGCezDfUDympmx1JpbxWNGQ3LrrcXWSWA0H1v+16zMGm6G2TuNrG1/TokWLbmJ2
UQw39Gj7Doexw/h4Y8jMwhdAo9K9qSqmtB4TjN4ir9Rk6AmNULscoNPlcE+WVU6j
hpxvhzCA5aA5Ut/FvmLweLyIjL/Y7/GGOjsxROD1Wgg6M5X1VERbyKLJAjyCtP1R
NBdRw7UZgEMn462Ati7sw5cf25wAx9SyliHxG7Y5qIeZoOR2Orhwc93V4gHAzJFj
nkDQGINrvcN2Ldq5GA2CsQip4XP+3seMyR0rpvkHKNILSSJOMOGoAMUsbJ/9bE22
nZiVEkV7pj6zEou/j0Pb5QKSs6qD5Wg23aNJfynpPT05javhfN2LstlqrbghPnQc
EgoKxJI/ueEQF/qMj3dFJskDEa8b9Hbs/XixhKZNMZ/Kx+aUVkPGuzwppEzTijQY
7driTW6kduEUiKVM2jiO0q8P23ypAfXcwD+AsHlEnUaRxvM1eKHhepcCilNpckgx
34TFSME1DzZI4vQ4KEj2MDQcGQ4wJbMJnBiCdETXX1qM3QtJYdznKc242PIlGwxK
EFtabNPGLIG1lMX9a7mCw0X6uD8Al/AFhA85wamkfN8iW/ZV1Ime7/NLptKH06yX
ptAFAOBB/2jsyPPzPFApjQNekowUqrI806u520swHSza9ugvOzNi88flDbYMf8Gp
R2ba77uUxo074NWCVXrjHPjvgKGxn+6hi4CQ9ZUemtEWhT0vzUQ9oGN1pvEGq87d
3Rsg6/0W2b3k/vskdFOnM7B8p6oTqxVwV1ZJKPSW4ru9+f1w98S9AciouvO6Vga+
VS8Ha0/6ZWIT0/o+82B0TgoKuNfywHQgRYLdDwoqAyAoy2nTSaDHWzhDcUkjMyIG
ES36nP5ZNXE9MkWltyuY3nik+xeN96RLw9vV+qLQuEkLy71MkLrUSX6ng2np4j7X
UcbzqDTGuZGDmJxhxI48Bi3XF9KffFDva/KZ9kksJCINxEYuqvyp5r/vrD8C/fqO
EnHdvM5iAhes9B6QabO47Jeu6q034viVF5Dq7QNUWcoqZpBSvTYzMKsj7ZU8BSRq
75aoSzDXWp8QOcedeedU+BKZiKq8paqyllRpqbjI3pMpnZMD08BkPYw3vQaMMs8U
GtAozjR3v88r+xs4K3Iqg/7AMAbbFNslatDn2HS+QyXvApO5DzdBW5IDVEF6iPXt
vAF6cv+P2avrebiCmCmey7sv9rGXCRSqHswQND2HbL61P7+5ri5RmbH1lbRXv6fB
wo4s8yxBLGX7OdR4nn1JTG616j1vYlpKbSICr3ZPKQ7Q2Zj3OLLvw/zepY/zsFLN
o/HhhTzVpKOOG94U0Buo8na5CV0UfSUmk+CSDVfIsujugOzbvNXGJaOx4Dz7afqW
KVChahqfR5v4xD2VdRjFNPgAt/kA2yw6XHfgJIPfdDN5Z8nik4N2mIZo0/0qZhW2
lireZiESnOZ0+Wpzd7fvtnk6hjA4ShOwGC1wkmDpEkG5UEs8d8wnzPxd/wIWUud4
l/s+zJsxb6HKUweGBeYDL7xQCD28bhiLXiQWf2hZwEC6Q4WOWvpEjxseKzfmAbRx
lmrJIVdJCl/5ASpWTHr5sKs7O1M5GkXxOdqNmqPr1SuXddRuSJTMfBwOQ4DyqOet
IEUSsjm3p8IdjNmjMruflHxoPsh4oT4su+vJHaBuaY3j/nNHTIgtES8vjIM2E9JL
RFL/zLGvdaEz6zmjYN/8GIsYxwFGakqbusfgm+CWC/cxmN10cOO22EZ8ySwHowwG
fYrsILdv4uRzTKIXZDO+8fMx9vyZ9cF0R77QDw3z4W1pFczPqYiIfOusKozSzHVF
twe+cMFU+eQdqhfXuI8tdKIVPItMxv/dfF13qaAFwYo3KCMwIr6OQoDj+7u00flM
opi+kGSLWzUhb3WLUNAiLUiFyNOazYD63N5WGuxCI5e9tdXafIOTltNJw+eLqwbk
RAHfsKZuWhWYqWdnXozvWMqnh0wmYB4JAMoUezDizmh/JsA3bDG8sLVz8L719y79
B9JybcQg4+seSUsPNqn1ZMGQh1DGr2uhI0W/aqFhBePz1fOTFZ9zA6U27tr9cp0f
6Oxe9acZFdPyR1YJxRIFxyibKYRXLliXbGOMvl8KELw4/HykrtcUMJIyRi9C/Syc
xSmMa7eeB/0znW0KPenwpXZqO2l8+JIWViLsOsgtRwg0SN61N71pt9Wb748Y6/kd
mXn+TuVZ0s4s6oVVL1A95F9Mo3JpCIfrOiEDjtKM73XOvsMijrcmSUyOBRcEbUjf
PUwtbTdiAoqF1kEs6Yizx4BljWmLOXmMTi2fEtRysMoeSCUmOv61QswndXzKHcxH
+x194wtY3x/UT8xxGqbMRlW4gi+ZgJ+wbAV8uODDARmxtOcRlgdyvcXXpXaITF4p
2q/NeHdjCkCyRMKuKvLFCQQ1J+5t2A+hJ9s0Mg9Gd760OOpU8LynMgjmgRg8/NVj
9WvtqXfrYgzqJdLKfwcbzF9BiNW1ARf+WPrb9QPPWCxZkWFwsTXnf1nu0Bj83pVC
MSDzMMGEsf/qJSMvB5lxkA9vdd535U8cEhloFc8cgXTu0WxXdLK21DcLFAsuA9j0
WC8WYKcBwj80eLkBugvDS0dREmaif747nQNIlIYgqMPe9mJFccU4+dsabPBSTtZ0
I8WFQAVLfwmgzqR5iL16mLq8D9MEN7fUdYdR1X0Kv9Yd84I55uiKbY/EuCsBq39O
tEeZG+BQZ+IMWCcFXn0JfgRSKYEV4bWnp3mf98ixBvA9dRd2BtQPLBpFf3w/J7uS
l1kxKGV1VhVVNNMd/LSfb9EESv/H2T9eSzYzjN5sQbpad1/Oow3twqVtbZlLnDIG
11ihO8LldOAz+yI+dXPsa/3crL0D6m1Bl82dHiv+jR8nvCjFWEyjzJBi6Eb/MuHb
ejYA4nkasecUmBw5wV9kGV0r1fCtOgOlKvDZSIa68VgrgrnAoGY5IMwk5j/T4eUC
6f4Lt/LOPCUjo++9mujygDvKQb95BQ6s14xReSJggLEa1j1VeR4Fl6cDAdjFhhzC
bLymIm17S5LgrEAiEfwUazrOIBI5nMwVKyNFkeXTZ6b00NbtB/LNc0WEC8WaIYEd
Hh94c+gnegP8GWSefoxPKa4LmOY0lPA7ENoHGHg+ShqSkQhNsEzGj//gJ20rinQ3
bWKSfByjHFhLsUHgXOm9qIVCofMmNIt52Li3JPO2OTsx4TRZ/xgMlBN23P9W2OQO
nNy/zDYEAfkT32puq5VkuHZI/TIgZMhZC7WR956n1MKLQihDnd/0n9WGCHT2H7d1
S5/BeeBjzMgjeLh9px3oNibd0YiFmJqC0zHNa58vjBpZriqgHYqFmogNgQ+4w+Fl
O0GiKWQGUjhP+6hl9vplf7nVGXtjIh4knu8XltmXsMmZOzXNJXsRjQl5IXT5bvWE
dSqAYzRY32romqRXWWBc2o5xdfpa0LcAbalhoT2r4TNDFXijdKazBUkWcFrU0z3F
FGkKJUnIJ0m7xfN0ro8ikxK2txb11vxe+/rUBUrGKER3utg7wNY0M2+3e//UMKEN
qulLbQ9LptMU1NtPc7V26IVMnKYE95apoPJgSO7k7LOnc3LUPOt4LUh5lSYVknLR
i3tYWFMZXido7MchuLt2P1x8dNCX2S8KVycrpWRLWna/S7YUxryXdcQRMQZ33SNV
dVPY6os8ScYdrCdUhBJmfEmNIIGCkL7tMXGMLh7VbXNk5fi8sHddiI+hB0yULki9
HH8qfRulHcWjbtF/TVlHGGV8UBT1m5rTn9ufJ6XTuIDZxnYxRCNomwZDQJIGYjWr
LB5K43EqA3zujNCjt4xK2ZkOVi0LSjURB8vn9PP6CiDTZfGAdyfMZnF1NVGz/Vj6
Q3BnHcLWtvaeAScIISNiOZVDJTAUuYMVvrKzcZDs7/POQl62O7Wr58hAWo1Rgw1V
UhzuGNV5Lsn4YupNhskI5pgO4mVfWdDuNzwH2j+Qd2jRJgxjwYev4Jo5RQQLEWIZ
H8CWHfKNeOfOIIrN1ZxDYIi0ZpTv0VQUvaWqocmjsMkKfxvUiY1wb1bsVN6yHP+0
E6/xy024zvOKMNxVtkYauuIlK1kDhw2WmXJJf1rRRlouND72jvDaik11jmBNCeVy
QP8jjJSf9lCNs4c8ZxB+kUGJBFdG3wKiJQEPxQdDpfHBMkm3VUzi09ktlITwO3pH
r7DMlPmJGx0pzTWKH3QcGRwkCq04X8t3Z8bl+dxzyWjeZZRc34hWI88X//VHNlkp
rlGMqS8idBaTPco9qhZVwMlH0X8d9JcmpxDbPjrstiMjN8hCujioAO/drFUS8nuU
AYNqOZ1wNOPXB9vFSJweX6kCqxubbbuNP+d/j5Y8m/QwFg6JtGRwrp1gof2+nEYB
wLQIOCRTkOBCHWcmxzxTypOcnpI7eS5oQTOcO6sJhp1GWIYf6MubzMzxRGTl4/5f
ACfB8FPy8QHa/L3N6Q/BG2qAJzAKTDi2DW1LFCQUK6B6c0ez84ZS0kqyVsRIUrq7
rjTeu6DIP2hApan6K602FQIRkWSfRkTPvENZ+tyRWIuAzw3G+jKZmYqfLmJRIPg7
Y+Or3TLHjJzQgVcoR4luariHM/5lpcPXLMxQlAg80jhzFHXh7KMdt6CeOkD+2oOk
CSU76OXqyG49fsPPUVkjF3659mdtt3popdWRv0VulBZKQIjtAaeOAwmK5oya9lcy
9XWaKXE7bd1tD3TVerX2RhBkx1uJSj1LM3k5JTD6DOkxsxuPesA9eWlU2J6XVnZW
IW7al+ZHqDfvnBeZMJlF1bg0hc9lFLsDR9eFXiy4Px1rKSXlkboTHzD5ExkkMr3i
/0AWUoLX4iu+4/GkZoX9SZZKaeg3/ieRsWAbQsKz3EAu0gVdXluL91OeiR499+rH
j1Mvh3flUh0ZCoYq+D9WbeUdxxJ/B72bWA5pXD/v6XNFLUF3X6kTYl8jLhRdwId/
lycK6cjXq23IsM8egNp0AdbA+nuU5gAPEeYhxR2YmV3ffdshbGVE8GegFJa5EVa1
qjCtbnysn+5ju1YBAKVNRH+djbF3uKESiBYdzEOEOPp75iFKUUuCAFwh7ivAhPCm
xOkRGvXzmxMHCWxP0ygUiKJRAzJt+0ujsnY12oWYFiJiVWDA5n5HHDqMyF70J3xM
XvqBUEq73c4+IFC0Fdx+UAvJkUZmuFRJFeGTQn5lC2pZ7GR9Xw/14SuxB2cC13SY
jhXzeipT+VboXXzfUOsQ5uoKuLPffhuPOn/EPob3Bht4Ag81SBfBvivGJRkp+3FE
Yj4TpB1QcHE8+030bVORhaMYKHRHsofvyMG1f1UA73eGzfFBtqvL+qHVHsBuj0++
ASUblZa7twnElxhp6mYmp8cJi2AOakzbQJ7uXwa7mh3G3woYGEWNcUO69AX7rCpd
h6vMoXgFs/OS5owLNQ9uaSGRtBso3wZtv0u6atSq7b2ed2JMfULoDm+9R75yy+3f
hbL3bGHWd2IWm0bldV9XGqPWBlonavj+U9AC+4tnMImXuyOETyhRl4Yp7wKSFthC
oAheHcvg+WgdyXXvvmpMhdHx6yCThrCyhklQzNPZrT2eMcNuwZuqxC3wTu0Eb286
c63LOi/WmCjI9yq2Us5UUpIlKcmiydjJflG3bCNzjYrrcwRv6c6VQg0B31amF+kY
aYdunWmMkkYtn+zrXjpax49wzYappaez2KX1K0j2614GUngJnsR+OFGeY52yVLIJ
57djt+GtTeRMuVQ7SRI1nVBBxU91DgM+e44dHjobM4qjsQCIwGh1RBa9DKpV5tOT
ZxQcEJzE8oKL4wpUvSI2Qi3PD3iIWyT2VH2AkW8zKQqMOWOqdt9GOQrrc+ASLWX5
69ebdSpsTB8RARgHp62HPkpzcFjW7fwzO0FD5cHHPXuOjsZH7NEadOW4XxMUohlP
w9p0cmhRvTEvDVble+CgBwTOh95xn6hybJ0LzUFfMQpGHIQn61yUF212bzZjtW6Q
a9hg5tVcTGbpPIzJ5vv9Zc+ZUtxy2t1AlwXN2B7xM/x3/bTijBYasLhlgu7Q7B5s
Vj2UvaVrXr6tjf8oEnfNc8uhURZyQuGHOm55LLB/O/es1q4ePBo7LAE2cQwwPDXR
pQuAqbRc4tJYCr3mwIXTigS7zUYArtfPCj2axNrkDKu9DZ0vtb2iz/L1HlZrU+7a
F4YHKV6zkIC95PN/QiQqxc+ubRoYz6ivjfQxOquw/ThSnuMrXEWdOMbEioxWpck7
sy/WLQt/aXSRMjVI5vSnN41Ch9kf1Lox3SP/UzV3vw9W1X8kd10pDcDvxA9l2QQM
xOScWfucLjhuyRXS9M3N3Wz2XdAOFflCi68Z4NSIpg/SIDMF14SRhf0mtXH2S9Qy
PAZzL8ULQc7x6XQWvAofKkhYwXTN/eHiv0O+dOmwe0pjb+GmV4XuL9iMY3HIK4CH
NBDjN7bOkhE6zJVrGCyLjUz9Nt5yaBxNQN8CIonLKXGneRIifbS/tY4voYLPq9LI
DB0Ns8xk98smeWm5oxU5uACn0oymjWfwDbT0VMKdLSzI7dPz6ZcThA//vSoGdrVQ
0uYllXMWnJA3FL2IrF/ttZyaF1zccvaSzXj/iFTA5Bf2uT7pLaMCz/1ZP36ejhUn
5mACXrj0IYkLpzpP551XCtpr+hsbh1rHDM6wlq+o1hJDfhINBgLN36CavnWYiUZP
HuoPeApvna6NLDPvZURT4hoGYKlWuKl/lPP2DZjt0lkOZoCuRm8f8AhWRPBERpKW
361eoeKJ5GqJr4qTfdaAFiJcv1LD84dSBwuvXXLs5tKOqyUpA7FVfY/MbdJF3TA9
b3+Iww/qEapAcYEznpAEO6nh49wsdhjzxXSIYIM/VjOGvFkdDGU5JFPhfTH8YOPu
xSAOtJb4kX5eG88K+w9XE3ENP5cx/cqr3SpnlRdRehPfGbUXN1GkOKALKZaLS/ei
ZbmSoaK6im3PJHDE9WV0taxYAj3rb2YBNVE1OXQtUyR8qk5ogqGbXJsOF3O5vWYo
L6IVMUgZNbeWBCryox5Oz0pfkL5i+llczz6yQpJtLWqQrg1doqoz82FNBfaJz+M6
e7rL6d0fCv2L9Qgu+B0EmZc3FiyDPxyNRNHALmhk7b/fOj9lgydeUGnqlClyXB3Z
D0hzsl1dt2N4jSxzBl1h6cEPTyJQCa1NqQ1U2O/F7A9zR8lBynBEBPVQxG6wM/o7
Fo1xHJ+ninbX+8cj7VXu3q3Mgjl8krBrcrfO/awI4xaw1mEFq/1Cu/LRn4Y+Y5kZ
i8jfXLM49txhW1OdV8f06IAx1VFtXM5TpeaoQGJX57MrtEQrAANL0BDu+g18omQm
Rb3LkBXbs0YXXj9xvmKwQ46/W/yXyXEXfp62J2Nc6EOv/Hin7DluVHpr482j+E1W
GYPJRHul8sGUXNupzFe8MLT+TWPz5BRLzmNxmFzh2pM2RzuG9Ty4eXBMhs5lUB2E
yjoyR09NvLkGtIAiKiGeq2eOP7bsPhGATVKESldYulC2x5zlKnjSEBBKCep0Uk/i
Ax+CN+vs1RRvaa212fmDdmtL+CFPxsRepZ7tW7qrglAUmLFNsU1pF2NTvfqTn9yq
DgOuQm6e07psRIZK5zEhxL9yk1ZadhN1JsaJj/nvfbnoPj3CC6DYm4A6mv25oQL9
EVHH33VxzeIbD0pZrotkhHzaJGdVZOacWmfzCmXNPhOYPKQTpNAhwSppSrj8QrGZ
6FwFM/Yaxz5pCjj4q8FhiNmN8CRBGet1fj03vjS5eRla7y9K6H/twdCeD1w4EVoM
mR6MwHMbLptIOlVVnv9xd5fQpl1sEScZoJrwAlgLcphViAkA0zzZyWvV7AidwvHq
Mj5v9ZFkp1b2iiVdGfHp1/1ZEKYQ/oTM1wzahbYHj7QVfr5duoz4qYNDQjInWcs7
uTayKOy5xFMipOTlizZsQLvcNhNxLqSuYR8vpx7Io0vhU5oQOJ8N7TsHbJkwOITm
GGPTPnFjlQYPIcRi19HbJ0tcRh5pYxgTBzknC46PrOCjPQgY26bPggskFDYnPt0U
6Wi57os1So9XNPfEp2V1TRVBQrvfNXpHPiI+uFsRgX+iLYlX0dKmlosvbMjz+2E/
PA4qAbFsJwa3wA6tlxZOR7npiUKQuNmXWA4etM46qxTOanMukItejBniG/RbU+ar
Nlg0TZeesvYcMhjECBDVGKjr1FiwZEbOOcK2Qr3uRJE85aeTmqmLRhePj5CdECyA
Qcp+78u7Ek/UCcJs80NeEn0Qxz7s8KG2eHDzdxxeY/aijssQ/0Ezz0Qy1Xl2oj6M
CSL1DZJzzUfHUsF+JZFFtV2geYXjTar9uaB+gWSshCkoHEkRP2gmOgm2ntenW5aF
jxp4hY8+zYOYqJgNVpjmoqMpEGwvtHJii4P4PhAZC3GrmvBYkkwNxBVXPjM2qDj6
lTVCbFWkwt+WKoilSGp6R3uW6ppIg1A5nFXw67R0oF5Y/ljsIkxyDNsCTchvQtOr
goB8Dol4alLhugvhchmVoFf1tGYhqrZUuvy7QV0NTIDExzQVJEllS2SxC8SVtV7T
LM1t6OXBRNvDaGzArPf3VoZCXVSjOdvLZwNxG9zL/vcUM3rHgEWSMHsKMij3Ce2o
ct0zIde51oJ3zZppUXjaiKAhlQe8VgWmkVToHL4gJ054nNl8qeidaNvxWT5slGGk
lIdVPd00/3Z8Mu0RmeZkgx0d0N2A0F6F9dcwXduqnJQQe4ZGLN+mef3HOIMmZxu/
/tX0VYTcRe2wSWXUEgWOisKxDGr6MojMimy+RmQOaDRnTcJOkadSWgFGsMRMi6dY
/U0nwj2L8iGLxSD/mlmsskJGLN27YuIybmilw3HBotootngUivtXKWMHEShbGkOx
Rb6W49UblrFf7kaleYVXeebvwEeBxjpyKUyhMpEcBcSDUM5iURgi0pRhM9Mb33ZL
heW7FnjpY3IiFgKDiRiha4zfpH+vE9v3GPrUd6qJz0KLeymd5t0/XY0/jrggIaY2
bgNbpaOPSSI26WFts0n8S5WIdgLMbiitGrC2NMMJqc3FT9aZewsDlGLteQmBXGjG
oq8KDeOOnDsHgMJKvBarj8ml//OmRBRjzmA5dYxcTsGSxemFe8qojGyO5/uf/Gl8
w4peiy86JVSHW9Awf7IJlc9O2tOA/dq3BvWHGVh14ZwJGShu+Uvhbsck6Js2IIM0
loOulh2rfNzxiUaZl9Rt99gY63kKB1K1RFWCwvq7eaoeHTtd123pVh95fQOx7Mtr
RYZmwkuM3yPqdJg/WUrRwPcwFOPjJPhliTenjgYfT2h4AQPC+kFGeo2hwzW9atZD
Tbj1SnCxNR2VdILvMDYHChVE5fQ5cspy8o0qrXC6/pU3bszFKtXQggDXGrPu9luq
Nnr5j6yEbiyViirmA+giejmow+eXGXNyg9qrjbyjLdoG9WzFV061qFGqwXh4yoCj
zGDyXcSYPaSbhs0T0sQpEDpBpHbqJ7N+lh5h539JBmaLjRJjV+NwT+aNB9MePHSL
S89BA3HfCujwVM8EU8VS3Y5i+PdwjxwA68ACjATX8IDtF4+ic6AafBjk6Io43MQL
fYMwLTbk1K10N4bcSMQ8tF9a+tzlKfgJKuuihuaFHOojQxmvfkfKXl5nUUQIbrMp
cdMSk8X8uauCWg0U1RL5Fb17OyiiNL5MNinZ7EMaHGD2ZSTQ5VHjbrc8aXgtTpFp
aXyy/G3B+/xMvyL7Jovh4nFvu1+w3Moxer/i/Q9qMPBMPr3k85IB1yeqN73dmaz7
0Qu3m8PvIY2FJVJMbLP9Ov6D6tiLhLIUiTz8QzT71kSKGQ42YsGsv2ImXQMPbbk6
azMeN4lRhI//RfQLdyVlPjhe2MW/iftYEBB19zUUVeDTagMqvf2IyiUfk3CZBV72
nZQD/qix3k3LRb6w2YuU21glxSjUqL3lDsHuHDjFkj5GGaluqZrpvHw9G/vxMPnv
dtW7BPu999oa8Z4s1rETWK5Ry2//rravquNf9fN75hQpGy63aihWz2HFihSGvOu+
54AjXdBxVM6WZY6XwxC7MOOap3Mo5LFOrt0SgKMMnyLf93r3X/vRekXVQ6SC/vhh
5hIOqPyD2vzqR+v1sH2wjLSc4NpPbexGB33aHT4ucw7wRbYtpuNyGzUOES7oy/u7
movOY0qir3XoxRnm/H1F3ygwhd0hkL5/xFEfNHsrzoZvBuNKhc1h59lVRJOUvs8z
ttjdOgsyqHqKLRsmLusxhkBOGXEPNPWLHu+jVxxRboc0ytqM443j4sIUCl71NMUI
Mjw3B2B9RYDHG74YwKTyNHvBUqm/eZ5Rl8e/RM+2fDDCz+jpOzYLUrKXyGVp3RAO
ljbfgvd8WO0rknBGR9JP3V9cy7sjKf/b71UoJeZA8IDrE5kJ2qdwEzGp9mZpsTUo
S6EqbU3AUaSgsTh9LvKs7o0JHQgUZOT4O+B8JHqen5LGAXN9CV5j4HCAlHu422uV
ywcf/iFbLY75sc5cB+owEENdQ/pCXhU1zwETqmZC3yuDeAYtuXtYCtM2aHXQJ5k+
IL5VeJWIZZz339sZ5HuBYXl1CrcFsLLd7ngkPzyAKH6gsNxnMokDTPR4bxPzndBc
w180TKKCw3bg4z/lFmLY3ATT0meZ5vp+xMj/3zoJcvOmotly7vvV8G7+vXZcV5s0
9hghKRQrLEPqWtpvb2sEsecM55kX+ubWj8oln8x3/3spa90e+jmuBGsmiVZWqKNf
jnbBqdeNpxVm1tz85U4LkGdbjxLCrPGfVSnKthZZuvfTf/e6pf/tuBNzNHuRAVTe
/XB1vg4k9ZYu/WnTUHNKqckFqVd7VHBJ0LyY6SDePZRD7WCrfeiFIdeDpSXJ5Wwz
h3wPZgVCCftvzpMiuzbooSh+jyLE1Lc3rGWGpPDTbMMXVCtMuEPZGSVAl5XjpOhj
IhRhW49D4a4T5XIOFTc5MgLcdmcRiHCHPOg4iFSo4Ir08x89RFItykIUohHmSrWA
/WdeZMNY1PmEn0oV6pSofOFkH3+yMyXmrwvAswB20KWreYpuOViCDpopbV7mhl+Q
s0y/AFRsE2nAXfhlILO5hJZRUQ35GCU3q1FGNvR7rdfLZcYvLEoD14NVrxdL8Sy7
VyeeGQvbOCSlwUom7R54X3gKQjiqjAvhX+4oIWtCYJ8Q+PfHT/biPpXKgqh1QSBq
HFdHFK3KVDm4PLGAkBIfLFdf7Em6DVj9jCUdbphchcB4L1ogKNxYQqN6Jy5+J3Ie
ND5giWlKM4V7Le/DiGpHRmUli6FuEzjfNrUUNQfJj4qQUdd3DyvnU4CBG8Y1VXUt
nRIEbvAbLk/jlb7VZqzNscm3m0uf/jdwElRhdGzAB3jHyC6Jj1uXiQKD30T/KRe9
Ho0p2E7NB1mIxKFIv3lZFjwpLtp4p9iIWhqic7Lv+RkmvLgFPGqelb7f7N3r0pYJ
C1oyIE+3RZux2+Sm9K3C6hj/zh2oBxChipkojh70cWG+dZ0Fler7xuloMRHd7Tzu
GXYK9AzFGDVP0AsgI8lBbKzBbyNW8TLGWiMi+/4+SZPTJtCoojv7SV/KnnUwPoWI
hnyU2OL3oosBV4L870Uea4lS2iuTL/LY7eroch1JnI6WVp93FD8q02mCh669X5on
nm0nqzE2v5NGvdjuhWjEjFrcHUsUZbcZQk+41Y60RczwZ0OEIi4TY1mN1yrwbUEc
WHfZUpCwc1eq8mz1PVOeu/2sxL7UbCCg9UwgzhUiEbislBTAu3Vm3ArGBCpRU9nM
/855AjTK+X28jlMsBArQXkE3bjhgkjbOvzW3S2+mtrIPwKSDb1ZHzBDc8w9hajAr
CgwLVOBLPlpDYUQykZe+H3yQ262qFLeVE8g7ZfzmJ+7bzMWf/tdjzJYAWZW1ap+K
rwIVC5Auh7vfzASrKDkBoUfzTg2bvN4JtEmN/XfNHaDLwbytDGsCEbcN5gryGdQo
ZpSfmi1dQ6FZk5nENg2cfF1JPM7mq1mXwWRfiNOEIzXuM6UViZx6R2bmEk8dJRrK
t3aStGm3xZOku1bzBmczYQ/rsuJ8qgORdED1fnt25BsJi7s8yfy6ItaCca1V2RLu
vvlFNbw3jA/QTkuQJazHxm+1nrFz3VS5NAGQ3N/RCQtyLhc50BXuJ4UL6lUqXIQV
uPtbuGhcTfRIDI5hxmi5ydRevcvq7dWX9OTm5anXBBCnkk/xg4HkxT8c4SL1MyWo
wCcNwQijcUnb2nTvzbwNyc4xeSAoVgtyHg0GfwaCtorn0aGmBnh6kyO6KlK1aBDz
Gtg60Ta9jL7uFMLg+0DFf/x6pwwMTxpeuK2Wz4+EYdde7xtmx7R65ARwD5HIE4z0
ueGvBevuZ/XME59w3hfS+fKbWKYryML7IAj2X6V2KscRqoGgLC717Hnqh8FCBT/S
6dkNF2dxeA0rwlK/3iJGlNDpY38y/Wok5PrenfBqtaJSNK8F4kQJZYjhGRAZnJQ2
bihJfYiLb9oZpIiXCEGnWq1bJeDNRZ8mLYnoozrY17TOE5gYnZlIexKJQxLH0XHU
BXim5GAjfYX3gPiJ4qGRBtPYoLhs6CC3cWhGv0DNjKrEuu0BRIS67XFS77nBeYYx
7O9z24w9R3JYn0lh+6/9otRRrphlKZNlU6jHrs5VclF6IinTsm4mtRQCg9NJkJ/u
s/zHzkoIV6fsavRu2dCOTmGe0LqA783q85XZZ61jwdDweZ42Yr7kOP/ZWedFj6v7
tuYw+JKhSF322b87HuwKjkjN4H8xNwQQ97rLDLyapOm+baz82WaYlIwRdKtYqu+9
jcC/FawM8xjAQh+xbBAwRJo5WIzU5P2RJC9phCfxv8xd3CNfTKKyHIu1gJKOYwv7
kU9I5xn6g6PoITkbujoZm620SOf5TXR2g1V6JMF0cE9q7g4pooeZ8TKzUoYTnBXR
yc3E4kolZN++r/SPhCBTyRPIY4ZDHRIuhB5x02EJlHYrX6G/KHDTdIVJr4hA/WxP
AtmacUqhPKHYMTAYCDKZpxtARUoy7MRnwVtuupa2s2Pmv+3YO1f60FS1kdpkAJAC
77a1St/Ydzvp/604T/Pb2Cxicf7YNCVRwYRagiT95cZLEkHDv6PY67vBFMN/ebRX
Ern60YS5P7Q9ECEOl2dWpM0Ab1clJC4az20pyJh7Wqy1mpQ60uL2cLnptM6XlI2B
3DbM7qfZkPXuSqhsvNiNCjNpKABT5P0NvsU2Uj/VKVeKCPcq0KRn1W3zgpqAxJ+5
i9Fg8uik94zRLyytWRbkMUsiNeo6hjOCseMx//py0ZWcchBuc8piBLGgbSt2RzO+
naYME3bOD5c8PPsx6lU8CEbpAKOHWDjuv87wNvpHX/kUhPqksPvVzAXWPVrgdDFc
i4UPbmvdejuP6ZaNYaflu/UBDWtHkx/cISl14M3nJmccNeapbD0Y9LaLqdbojlBq
AfAHqN3mJasyDshzFl4mCUIUXrz/pb4fo1F6MSjChkJNFvrTkqtJaN87WCx2yGkM
iEtsBQbksmUuknxuGcCHVkkvh8sIoJB5AKlsHiwj/Tcl3HrjBUJYI6El9TNDg85f
zqNl8s9EpqOCcsbWXVQkCHhxggECVC3SizKniyjaSpH+/OWwD52GTW678bQBKoA3
rgxQ4SBChz6ckI3qLkP413b+sBCmuqoVy/6O6u9WJt0Sb1ZwnVTdgw8VVqxObpFK
CStqxfgCRN0TQ9KGCS5HGdT6cMOpRNAK7tYGGjqfwICPixtgRA3wqjEnjLoGOyeC
jzdhXTBCgcdNpmlI16jn/NVSOZkk8xm7l07n6A4lPtNgsUXzE8ow0As6ZZMFMxEW
i6Vjqg8s57uSfgNyHWAeYJYPIr4rMUtFNpr1cmwujGUmDNkQxvhrkul5zZGd9QOd
jZIKZ7XII1GzLzjSA6XQowrZHb+RL0y7Wyd7+hGbzavFEh+ebL7oli37m8ebLa4m
+FGTOduF+XxMu0EkkT792FJi9vA/rAM69jVzH8Doq+VcihSXvmX3KIaHpARnEgBg
UuO+tNOJ98yIPJ0rwBFQcLk6Amx8+/ADCE9dcuO+IaNfAi92eNWBDVCklfOQh5ua
Zsgt0osW+xaeW4qL/gJDDoCg3dCjZ6EA1gSCCOdttDht5eykrA2eyhwrZuf0yLZS
SXLhGsi8/WtsXfgyf6/JrzhdvZiz9I/eFwYNxpzwhVUt++VdrCQ50FG1zqxNOAK0
7AtwImDmuw2UFzeqVAgFBeIq4KEaqn4np2Rbw6wJeFfSfMHV+c1/83WLI6HvbfcS
OMV/6UBBVAgYN0V6UfxixBHwEZ4lGS1Zk/KjDPRPRB8E1dBSGUrmM2k3ikNWWo0u
Gq2zPdgBLM3rDI34/9A+u431xCedfenXx7y0IBAb1ChK3RUO/8uJ1nY6JPLRSZME
gpUeWYYj8mf6PQ+uAftlNGxMAPkMJQZRR2q6HsIPngKd8gBoHbUHLrGkTjIdozZi
8CM4fsfXhjVPKiTXPXPeEFxzFNw/pIdh1M4FqvGfNiuPsqAh7UGSK0RYczBDamfs
02QVmOtVbz9OBY1IuLtQzKmWmIIRrRYMPl+mx/V2I/dLnitmIcJ4r9IlXapQIWXl
svLrXb5TkCJeeqBQdPikT2apgzQVI0V6NWQb4Oz6/AevyDy72cv7QzBx0InHjjPI
Rryii9zIxruuaSjfIXCUo4cKWjQxopGBDFA0z0Hd+OPc6FDxgrbZi9xM0ufhqsVa
VJdzZim1e347JXUvHbZiu0fmXUgNP/pxQD6fm5Y4371GMChW2uhw6ly+qy4Zjl01
VEWqMOEApVT7xXhn6YlXzAzUOQ/DfKEFyqHgBr0Mh0d8JBVpIIE/3dtZONAFLs3Y
xDWO82JENqyxl5nyzoTfdTlcfsyy3i6b+r2R676srpRYXcBqWD+jfcD3JahXUQNp
4spE3UvKdQ2rdMiEEyLogWDuZdC9041SO5ExkreXYbZOfiNX/qR0jfnQC8QMOlRt
QprGwWS2HT4KcJHCBKJYfc9eEO1DE22Ww8XoDJKxD8T7MA9DEgKtTBE7t00g/rIb
LxgVMBNJHOihB3qC1EraF6eZEPHHdfrBcv7ii1NaV5/QjzaQ++UH9qMePRf/ZFpr
8H6mqkSZMCZTiXF5Bfl0X2ioXP5nTvI23u3CPvc5OQsQnYQWzJRWOySmN/HEl8E2
SdeSMczuulmnx6k1EhHurUkDoLz+ysV8+Bet6L7WaC4caXXSCxFgum64AP6hvqkj
O//d9AU5if5ieUbxo+HJDnof1jwp4t0nZn+cg4ceC+m4VIeHzSUkbkLpKu1NQgR5
vgXzXg3rBq1MJktw9eJ/2gS6kQboFv8zLKUui7XBXSy/XxDOJ52PlM9mZPeCUzu9
+nAy0UDUOei4Fhyd+rgRnHopdpNHn2wYkJsZFEnqoiW/ND7+7BHaSRRlQpSDkwbg
1h4cYpU2hgb7Oebj+0cGxn/or4fM/xuPt7/9DuzaR64FwgRkPQrFdrnX+4+DpfWU
nLx6IDzqSbVtxo6sITIEGqXXA+I/k8aY6ZsPEHvBkIqEKZfBvCkH5i25WtNpNGz4
ITndI3Pz+ggHQIiGoImNA887b54m/dbDn93VZaKP98DxPxJsrF8xUhdrr4xE4SoF
eourjBcDTQfwsD7H43TeUHdpAHx/gLJ6GXAQQJ0tAn1gzKG7KfCo591lfyg4GOIr
TFucwkpFPp7/ynfKmlMdwofFPY4NrGd1OuqyfX70uFyEvCvrpixtWQDX+F76259t
X54+gKR0cFjaQbrKkArovgNapesn2y+PAIcwkCKcOLjPw9NTgu4aVmI1GmPikmhM
/smG7UcFNDhjLIPgIeB5S3tYEQ/ngi4gb49wxhh6muSYehzW3tlsU2CuiPMWq7Qg
hWI+HLfeoEFjOgkvxEI0xfw1oV7SVh9bgC3w0cGwM38YUzSY6ovuwjZk2HC9tmYP
TvjkAmnXl+KOjZ1hVBBsm3Aqo79/gqkx63+OauWoohN1I5eBuHzwf0niZQbvh8w5
K3krHOy/esZoIADVxUfWbJ9UlwPpRTD9Z6xrPWFaHCh46TZkd4cEwDWpbXRDtEHO
xQFHakjjNl5oE3ujh8NrtK8Tgf0rRKgF1HODtbFKl27L+9Bh4FNBvEnPpbpgbCcV
kxq63SH/Wz7nSvjUqyl4XeeXjMqQsvqFslWnwWnusE4R5XHsiVzNyYEOzyG1YKPz
XYTOt+940P65GKe6yZu+KCSKAwGZLG1c6eFel8VzhGWWyrLwURAA9bE7+CckYifi
PlsOIhsk0dk9JK2g932Z6zBaiYEvar6OxXMiUxzu1Zijy76ndBDmUGKSdcmLnEXM
J+eG3MkABUVQJGPD4R6SKrMn905NMZbO3a5s9fYgGmSwPnxJF80bJgN7FeVhk383
Cp/XKtFKSAIkW3sMnM5h7LHZf7qDIu9cQk4T1cDDHcPvPxeQW6bkq7X141WhxS2X
4Lil9xej1HptJEsOwmukaZJR5H5/do25OiHdwEdI3WVUD8ihtcdDfbPrcZe+fJtm
tLyFy9+nQXRbtzOjzfbsTsazVOn3gj2ZC5wpMz3FEMDFs+Fid/TPpJbeF0hrvrxV
z+481aWALPJCC47QCUart6s3PQ9vbo38ABDOXzYmoXNVw0u1bEtrKudmgsT8AkCr
N2NVb+i6LqgrkG1Zq49M5kQ/zzlfhidA6Ai5+4kIS8Y1HOTiWwpbH92Vuysd02lY
LQrorKOOMgSG0qmEGYsbTSgkUNnN0VUMBFYykHOpqcis4f+iECApS5HshjvtP94v
OOPIyze3w2SY6B22IepBLxMgEB5OdGGKKsTPe/x4DiJmCM2CB4Xl6KOEStWcKJHK
do1MkI2A3NVIoJzlPWOk4DBQgVTcnR075hUXcZKvzJbygo0gRXsH2hraZSoZELxu
09JZVz1GBHQ5dH7R3U7jG96U2bozcSxCgDb5HQgW0eoZQf3Rd/qvOMtCHdDhPu7b
U+5y7VWZk0KWRKSQC3sN6Ugk7q1znhAMlUzn/eqrIkCIrbB044BLBOYAb5+WWbal
uZ/d0ngmdpJd42NQoauhKEUKoKoMLYO3WnMp2c54EiI+XNVu3KJQAz0hjE/r8ntl
fjUQ7CmYywcvPcFWccqXJbnULZOl97Y2cGgjzBAFa4IA413kM5BygE65zr/YAKgs
osLVCSfjMdS5NlU8uPdKWu1w1bSsifC+He4IdROhJFwMdSJiuk1knMp+AUdcnpbV
5nAHXX/1HfTGy7sqxsrINbrOn7K7XpNtob58OchSmpS9KPad3aYosVyWXuWeNyA9
z4tkMcHZyLFEaRFCjhxTBKKbHzzvBI1/FCY1Sr5b/wdASNKS6RIb/gfH1LGVSQDc
DunR9NnX2d9Pg4EbIWBLemrAmu1x1Q/Jdl/67ihOBmSawAva29feopGK43OWpvAz
Qbh9ZO2WFHSLSba+F83SCmZpNH9z0+AEfXPr5YhU5NjG1K28BtIZrBgsI/KL2/6C
zCzEPgWrBOF/ZN3FtpnGednD5pQoujN7Leso6cF3zYGvuJpYgtxUdps4JEeYalQk
MhsAlEtsJcfPhaxfvm67uy3hFAvVzEw9Bypq/GOL6YJDhT4cT+N4nizpnNxh+nKP
WI18qCTZ4b9YMp3OoEmhsICW6iGwlBzZAw2BHNKm9BOSspc+czvQnzdigrVHEHsT
y3uilKQlvnvVGyB4itYghPAtXdkY1eOklWS1dIhiv62ZkpCRgdNKtBTJlYBI0cHs
rfVQl0wLtfiSIFyMDxBgCOXfqqlEHoSG4MMcA3w0WsDY1b/92ZvwoqflWDne9H4R
MbecF9jeMslFQs1KkXajzbmgyShbzz00S1TL1T8LcA3G/EC1XMpbZUNQmnX/u34D
EMRJ2uRNOsHTe7CEumVxhtlhEJ+8W1MKvFrSTZYFaR/M6wakaAa3JTWO45BL7L4p
SHJbBC1ao4Got9yiGrTGPTmjD3Y8ePNXXrDestoRxq3a73bu8BS3iVcYTmlvXxI6
BWoy1RHPE0n36ml875IL5Wk4CUkdFOAqdiQ2HHKP+42AEuNzUt5SYqvb+o+BElBr
BBpw7USRvMX/NRwRrzTYX5KmFXEdjR2itPXSuoXMWLLv7J2STCxiohrp9wX4wAMP
vlVqqIU7J1JyaIGKdB7Nbgy2slVE5TeS2NLrnEg46tXL4Nn1j3dEsV4ZL84L9FFi
U83C15cUG6hCtPQ6bSxLHIY0pj4VPeK/2VugEljsJ7e8Zj0UaP7+f4AvEhujF+Ls
43ru7k+/h9oUGZrX7wSAJqjQdPBMQFX2VcAmhtATLMJ5qFmoWePiqUfxDOF6+w2O
Fj1j8GLO5rajp4omsTPXQWJId+hUby1A0V9mdcaDZuMj7zhoeCUtMXD+Bf4oJUdn
FWoEcDqvjsgzNkIW8sx5y8ybTw4lgJfVymouas7ErNCLmHFGIhMbWHKi0IFiGLps
i+9ZzexLnRBdgS76B01J6tiEET6AIKzbYoy+FUd9Ab1kKw3IaX5s+t4p6LcCevRP
vqxXbtgr6CbEhH/3pRivREwOcEHqtWiOgXYYUL4LdAsjHrxfotE9AOjDjLlbnevQ
6WieWDMWmYbiD2jVktqu0+WWckFm/tRS6WYTaJV0YKP5zUcBS11czQDFuQOdmKUD
UKvkNN5D6ZZ6UVDBKokj9m2Dri2qr52vK/Bsnyj6FSH3MKYf9u8DQU+Y8liJwEc8
xsVszfTQeF7Xh9JurylHTqKg6CLS2zTzEC3Fc2FpdomuL/7Cc+Zjc2/JtomrfFod
+PcjrnEFCJT9kW9RfUol9yiBEwH2VEa+nLYmIs9o6HuKREaKWsw5mVBhYmC+qy0s
isQdyLc8ZL3PzwB87ydAhVfKYBBrZUwkRRPgDuDBS2Rs+5wMPXJltGgU3ZaaX8Hr
aA0UzwJCJ0J/xY+O8QkjIrJg+yKF7cv2DcFFT8+lzljIcGjDDJ7EOt9wYSHKEHab
0tXPYZfQaXaHunvu/CiM/U48EQwB3LqurdIxMYfq4WFwxm+CKtaeBhmmHk5BmDoh
wKf2kh6hPdtc9YA58eq4vNeyPYRcgyr4dT93slxILrP3CyWhwfsM4ZpAsvHyymUT
J35bezonFd3cEenOl1QOloQYMiPRoG5irmBBG8gj5FglkXDl/FiECffQV/jEgYsc
CMR6qOEUSxQxo4vONiCZ+4cF+4ykQQKyhXUFh97Hj0T8+vQ3lCmefSv6hAbnF7Iv
RRfaUxZTj4hGna8U7vLMW7quf+mx0H3gx6oXFErd6TzjKM7C56hlFnKOZlcz/ny0
Cp+287r34TPyRUqcknt69xUlHLY6oNwXPyKMXHDL+Hf8rOlNlUTe+cKcSUatfAyU
Gq4GhwpdDqnM+DhNy1kzbJ2EusfODy7WdvY1N7KeJctB7ROO9DLXc4VlvWPtEmyt
78YCEeQYIJn6ww+NqmU2SO9s2ZyaYWRavYArWBjmKLOhb0W4aYc7hDpOKFJEqiva
1CdssEyLGKjvrcpOG8hWCjqf98kqgEEQ3uPloL8mCtrZeT6QzIsD7RYG+Qyatap5
//mqqldj+1P9LQXnvUIbo+ZKQxJXMOmozLgpFX47sig7iTxQ0eQ+qGoJFDeBPjX5
7gbWxSjTbi3V0IydsriQL6NyxP6kbCxpB1PISUArrb6JErYrQAL/4tFhkTryROIG
gYOI+LG5g+edB1EvbWWnNb3OgQehZ2oAJl1AJXmEyVqxrUCa3rRiUh5HRW1nNdKI
4EgQee31CNE8Ml8lLcBQBKswpoHXkG2Avv0JxPnaltZsUdm+kuSHrw3XmcTpVWDl
02FiXMxL6So/zlhsYxGD2pNR10QaeW5u+8PbC4XXLZvBu8CGyIEHjkBRuX8xQabU
tsy0e3L+J1A9AFANrAN2Fn7IMS2pKirlMs4Onw74UfblEEG29zXCDozGlGrJ8XJU
9jrXgMGbp//fWo87DvHyZCrkkgS605AYEG57rXO/U7YQay37p2I8XJelOo1Bh/jj
IjeHgaP9vxZFPVKSaz2vVxO6rKntq1ayspf76uNzmlA1IguXuFtUie4S/L/V4HSf
ezH5XE+Ct1Dc6YyojxS/FzIi4dqCu1NtM5Fk1Fzq1claHjBUn+nTHnfLlPQqDs35
Bvp9CP5fO0a4WwVpq2+L6LdCAvuupIQPKH16ct4wVal3rysjObLH0akr3+FGIthu
4QJ4AwBB2ZedF8WiYMvK9EbchzhmAAD84Xaevhn8MpOm8r3bEl66xqDluu/jltio
AVCOdBakqMFHQDyN39ljmsYcIKjJFNB5wpW79WNM67vbYkVIsqLjxG241PGD47yV
TPFKlJ1yadHH3Q9UimAiU/aX1p6yDXudUw6M76HT7Bip6GKMoiTu6EvEsGj/mdkJ
X9T0aXH1/xkk/7JbrgWO6UQuBKO2V9XSvRX+D2Bvl7Bb0QEzbezFL5KyND4fgC4Q
Xkt0IBgjEZMcTpyxQSf2Ux2IfDZIYBQDtAMiw2JDHNHeioyT49ZwAr4vYoYzz/0Y
hQlIbdAVasHUpU9iMD1A+fj34vtdA7FEGr+soRjsfjk+D7j7JfY4AdJsbvG75Kff
YmHhGIFZVYKHhXuvfVjm00vhFmIbsryo1O1BCM5rIk9CzPxVpV/CEiz4TE4LeDG3
gnRJjOT69BNSmOZrXi3VnvgjtTD4A2WU0qgYObtiabome25YsRDOWZPRylY61kG9
Kaj9WosC5VXwrr4y7tBRxqQxP1Z5hEVKC9f3uL7bIjBXfjgIAu5xuIvh7I2QuTR/
WpEe2xM2qMpKPzE5Kbdch4xzWVDhHifzHgdHMCkXbJlda2YzP8S/h7h9S48lc+bK
Hl+tQBELiXDK5CyFgprXu8kSHuZzKkdUbPWOAt0zHde0MzrQmXYvFy6RfTOI5iG3
Vz+sETqdZyrx5iyT6ELWdYYn2IYefoxN289dbCCu8sxJ5OcsEvc1gQX2Brwy2gER
KcoVvg3n1IiRlPqoJz5pWSc3l4sVAiMjDH7v/9L0bxUlWnapFdLt/8mvF9h0c1Tu
u4SOa/aWQFVG0YDubpb9jeuxNQ/YDhlZM2bGHwv1U+Es1vWW5YZdivpUxTMUmnD2
URs5iebPIJRQsS91Z9ddkuN7TzTFG89L7beFiXwWqJAoUDcjEj1PDX+2xX39qjB9
lbI8+LQZ7hUWzwGdaSzQwhqWPpo4bono3dP9YlPMKC0189o5Bl8GZU7jHBHn5gjt
E5jnCaLaNV5L09yBi+7PUciLkap1LvDbtwQZ2+amTtuwKWPC1VXmO7WPPMoEfgoX
wjNhK58KGFrPCpFYoPEnOmstQWTFAMlh3tax62Nj+frEqb4rY2asBo/Yf38xPvDU
USRUwHvi9VgR+4hS+UehHQbQ2ioenwhNxmaD5FJBF+VzS2VHz0dYh51i4W2Y7ExP
oixEH7KGEvgg1SegUTQJwxlWuhnj2YWF5kpTD5WspyQ6Tvnz1VNiDWQLHE9jB2sz
2fTp/wyPo8ca5KIRuHkWEohCLFBOGA64Hqjhst68Sacfq5FmmWU63fiXPMCcPesz
PylKG3685N9qQF4EbUWpExaYjCr0npQ1/U2KZ4hl0vlrwbyGwgGUWz/CQvVirKXV
kmnuqS8FXTOVp9KZ3u0FRofyHA5NyyhWsuqkKg8ttmh95TeUN7t0KxdasPvNTSks
ePxZNVChv4lkg4fRVUoK6icvFSbZGRBFfttqblZ6enTq+Qw7eAMcY3Dmacg/Qq9u
0exFH22zQlAPMRWn8kv0zHVnN79RH0miGv7jYnU1b/nGJKHu+Cxwba6oH/XzI4UU
NIjQkWjylLd6FcyjA1EHku3JomCPKgRgySNRueFk+hyU7YTP7TKqm3NlVIKVXP1n
rt0wAHIgzOMOD056DX2WSOcNdkSSTezIzE3hw9tjhYjdvks6aexINwBkVrAJpegG
6LI3SvZSNQ/JOhtrd2hbn8QwlDKDSe/TCOZ0oR2GlwgXRWC5A63l91TyahaUnvPm
lmoxj9GbWs+9zgDiwGO2gYP/tCalmK6VouKDfV+alZ5OEYkm11KjMlLyltulp6A4
XeqDXymoVpuYTqMAVRczH4CNWTZKnZDAQBBLPzet+JLlDoHzYHeaZGCCVlCEjGb9
mRh+vlHjh7AZfi5Hzz+S9ff1mlc3nXKvqatM6d4i6sBdERWBI77kwlzipTqezNs+
ZJHjK0PbN7kozD1uhvRyrTQQGSOlUq+v431soAOgIu85rlKEx44qeIvV6EqzcBsg
O0bSknHqOeZwItV5JrXIEaSmEEcfq6McDNDu3PyGErBE/FZnPseS0OJoqym8vz0s
BafUg+k0VTcyQ2p9xJzHUSHh3VvaSab6VbEBalNdrogHwxDXnrtKK1HAZUGhiIif
FbejzAHbaDFvoEkD8ZyiPwWfO8wa6aS2u0FhujFzf08HRo588CI3Sm7yaFtl5SXF
Sgf71yNLl8sqzEzJEnKErYubKSADKu08Isa2Bz1a4mK1v7ZIbThgrmHC/72tUOeQ
tio2XpGqJtzxMchJUlbnAJ9C5pF2tBrvPo+I2i4cnUrQNLw4oGcij7Fm7atHfP6P
CjiuRLwwPij8Zqdt4rTsjXphzKym74YTMMu3mWoWTNewKFM2QUyePMv0b6wm403E
tbR8ERt2+b5lcYQjJBKjiJ6ceZiXbiyqJBM3BfnPnfSm4PZ+bOjdESPNNEOpOsV8
x3JsBHtDSxMBILLllTrW6PLoByAqrRVkdX5GWEqd20cIh4+qCA7uyEvYylbMtPig
uRkQJ57RbkOv6Tf2g6Y2Ufis9GRwf0cqrDdl1ZAY5Kv1YB2Ss+TNApYGTa8bPEYD
RW6YW56gLN30uPSZDLhy14cgERXxudnvKIGNmw/G14HHCEFTl6ZBXHANsop/wPD9
gHwg6Rkco76zwd+ffsHiRxsdXCJwufaXEiQW3RjzfQiwNhAQWve4AuWj6sLfv3N5
KkvE7dc4FOwpYbfCNpmRonRzOF9Vb4F0Yo+eucRRJ4+/FNwgOUfzVAAK2kdZGkC1
lfuK+mrFG1Rj/QAubIzcQX3iK9c3nytqWKDZmn85AkOvTsbbPElGQRk7YJtwOh4A
A4JPulwyrQbfSLgNonhQwuFUcqQKUwYAUTB6/9LO4BU45hVa6lFpfzqyXOOKis2a
DP4yJVaCm7pm3Jhhqu8rLRhajiaPCCA6vGQOs/UU0l0B8KlyBpKh2zsuup25hSi8
C2vCf5h0QsV94w0plQ1b53ql0MTiEGbZmy8/9DNs+nDsJiDSq5xfmzpPXmrSPGOy
FeJFK1iNr5Pi1VdGMhtgTdDvs2dyMEeN1Ns0AhU5nEu1+HvKrEQEd9dc+zz9dlRw
pc3nfDMDrjw6xTfLccr3QSRztxQRMgwGpk0OSXYLptWWCBENnwpPRn27nuqPMBBR
2kAa/aw5z7DXYgIekOkXQd69tQpCNRKqNO7M0YM3qbv4AMYHuYQij6XpeQ10ZRYb
+J7LCaa9y0+xAWqcLfposY9q387bsNZr/2Ra//VNa7SsDQ3U+YEi9Zil8k8gQd4X
/WFX2tXalNhTthIto0CQiywKWoQanA6+CDHJ+3ZUOhFkJiDxjRLxXMQ04iZ/bOcr
ltYPS0oBnuf0XyKqRO0oR7UAdm8N9gNXLmZtZ5N+fV20o4+Gy/L8n7o+20jgmJS6
/NjUaAHeiQ1JGUWTj5lRdkTP7Gn/rvQw/VnHlzYH6l7MgqVPUFTa0Sjm1HJ3VUIO
vR781kf2plqWlYK/13jv1aK1IFRuE9qFzcB5LT41NCSwG2GfMovPV2SPEK8xwbSe
aOhj3IS8esBmmly3SI8wnhQex1YVhByrLrOVPdtMVboKnmqHvBjzIAnVX++Ty8yK
9czYKB+1ZqEOb1Yjh4no++vvne6TFnX1z7klmFiFWfXUEQtl52bN7U6QJO7JLMu+
4wtVNY6NcDLZaGNA5hHlupwTMkHL/LMKk7HfVoKX8zii4s0hNePMxgySftKyRlbs
CV6lOac+no29vr0hAbGJHujZ5OFUVoLQSPLCO/MlEiygiwiZe00Z2lxAvkh8pxQQ
4QovpY3B9vQ01qMduazgJ4vemxglPoq2XhEYnUlHkSCYDYRQeOkHN4gGE0Z/v1km
d4TSkYPbqjkwA181KTtiRFPhUddMg/MWJDRFRljWYavEJTjMaLIK/QWRG/vX5Gd0
MENb+WEp6haG8yt9qE+UETPSHbhN5MiAnYoItZ4XbmI8TjxFF2pXZRVop6/kv9/E
nWji4+ROiUZq4d3VQMgoqUr3AdTW6ZAxNyZFipJCs8pn2t827qEYI7HmkPJIhKOq
Ct+QBDbOtHf0epBttJcd4E7y3MfrxUNT1RQyEeNLK5zsMPtkUtbhA/v6PsLu0OkQ
NHJwpF7niCBptSWhkvz8SCpBlufqXhqZjTBkyNqP5NKQbKHKqQ5AiK82KhmBEdzw
PhDRgWiSAKQTlcgtpLGACdbWwi7bc7Z7Jfq8RSSCleNXamhd1zrOspEhfOR8PrQH
LvCCn41apPKkrn34Cz3C0HMPdLeVkbFFhYANjLBc5+ZyuoHPoIa6kB+EWfBRDPQ3
5Z/jJlUi/01Tm3SK1u74wySTI8az8AG5gaNJPVXmPMiHUIkETUHj+TESSdM5FOS7
p7m3Lh+kE0EnE6PlM3ihINRaOZ/uN11Grgbnks/sSsPuEcUjrBqtbaEOUFeu4d1g
X8CQ6DoCAsm6CRK4gyti7q7jPrHcczSgKFIgu38o2tbpD1+a5PNwOWir86cZpVxL
zurE5ZaEeHGjqnaOuQbD4UpIlQHh7IJJ883f365V4bpfm4MeTJvk0BZBX60EAiSv
7UTWqXRW0Zc5rBncIfsddBMnxa43VxJPHJ4OajannotbrEJmrIL5qinjZFBQRQOx
4O0AXU6iIQ8lKyA6+zf9Ukkoys8unky8FTpl0VGFN4nXcvZXO0M1WhbQ+ZG3eY5a
mgRuT4mvc9wuI3Hp47ntDTSf3lo4KM0FLhjHmpWVRx6xR0rzbRTMUhZdk0ZDhBk7
V0T4pzcavfF41VpxMbj9iE5FigOuLslPtJKWyVx/EVUJdZS6ML9mjz/Yz6DEIr+7
1M4OvhtZigkxDsSm3YMv56iCp8Gj1jKpQDKx51Mnmoshb5nAJ5/8SOM5WVzkHXqc
1KCqDc7a5wxngf24QY0nuV8zbG+vESnd0MOw96lpm6zaq+d2gu+VAThmHD+B4peL
RHI7swNblk3E1yMjaPkTHtE4l7XKe6POn3Zd4rBVjbg8RO4Ff4LEnjzzVu450EIS
OQ+kj5YyGS0bHHFzcDHeoclfzdox4R5b2MxW/XJ3OOw2/XJh/QxX4++r3JxB5JeB
318FTtmm3ysBp26VUAw5fffdLlbIHeimzLqAVdlvklr6MiZicYUaRMT3HfJyD2IJ
Vxc9L1z43gE0foLddZKRf1IOuWlSSPB4toetUxlUzMVSmh0yzmeQYuDqJewOuJWo
mDGShC+8M4AKndS3fmw2U9cmJSckiUnFu+jFw9b4CMCo2uvGG3KgyoSPULBe/wmp
Z2ZhriWOXGNxShu+yLCGrzef75u1MKVVIWJ50tHwBPTG4JxM7lT0urkoa76VE3K5
5826jddsbR2oBEdebG6kcDYr4amUXXGSW0v4UijVSK8qIuEYo3gyKNm9lang0ETd
uBVvV2a4GdxSZNbVqiu1+tk15Ff/l7zWNm6QtbqpyJi4NYAHgjwPbccVru3nLP25
4TiRVNBNFkbpBV3aIo4wmRhdtqs/tk2FmyifYWWshhDePZX1QBzWMDOes+aZ75PX
6pPm5H9QQtu6Ufpfew6H1ICFnpI4RI5WSbN7CXK3Q6wxeExpU4nHnueIg7Ukok1k
yNwE5ZY60AttfgIKEvHqAzAEPMcCJ2QjIFrfuPcHKZyBCjzNwM12dQa+WZQPH5lW
D6ZH2XrKeNlYfZ3t4LlBf0M5f5wn/TDCdXkwNemy7nNb8YoW2K8tH7WfIyIYY+Lw
U5cVcHUXiLjdB9rB9+/C/rpgXuUeOfHnJ5HkRQwmBH9Rp7XIKCCI6+NvB+WEIIyO
DTiw6sIXpRlWEl85h0MqIQpPiiu3VL3QMhMySdfqXsq2/H5klQAyPUOS9XgicAHq
ahjZWNMvTY7uUAqTWFtbg2/T6vbHNlTRh1w4JWrZLuj3/UhxP3cXvFKel826ie8H
UHbKOEbh+nGuZNbu+sPlD0Mp2eo3eaQTU6/2B08GagxQkacBSTLEmQqRsphg1b32
yF8Fy25NL9T95PibucOI4tT61FrHvNjjrqXYAPKL1Wf+8Wj/wo932tDAHGK/gOlV
wlQp8aARfjnkpw9y7ywgMXFPoOsTsUZkL++uNw8+UR19NesgedbETU9l+/pbiufG
ZCNTN58yeS4XyCWtmpqNH46jgRuxyndsM8LQqSlBAMhTBxf484lAxyHH8iZXfyBW
g9CK1SsBIJ8LwzOmG0IZB9dAPIIzCnXI59lUlNO8ahXFrYzW9uE/kyaLwvSQPYpq
NuwgnjC8PTpTmN1rFzthfICe5u8kbzAemAos30q4POzsjmoGDSDyjpE5ZlrqGEUU
daigG0ndgEScGYehO3gROMwfekwCMGXAhrYRN/XIL9Aaa8Zbp7V+iK5Q/UYMv9J2
gm+OL6T1HZQsyIA32O/slHgjgOk3Yr5CXmP5XPStcBHemTZiWAyX7pmNptZbpW+0
WZVDnbtvqELvKYlPbwr66leFlJRhwbAeVinzmZ3biN8yvfTxqdkHMDbq446wFmez
gA6OKRk0HrO+rtOT3Z7sfPWQjPn2h1LAPvhyCBzVZ94AkqQgZbZ9KBqK9w6/bYPs
8Bbrd8ZTbvKFO9l8E+7tJ7k7feluhIJaSpwWl0Ei4nczCxEcznmDVl02F2CiKy2H
BTlmXqroObVFsw1JOMoEs+9OC6VjC3SifHGuqRnvUP0MMAgjNsQI+kpalZg9zic/
OfeVUdHNWNSM/hYazdJzfWmVYdUufi3rzIQ14dv3cqtiGAyv0Ksx+8pNiED0dOQu
35SxjQ1ukj49ITmE/E1XqWxCbnnEx/FrOu/6kmoIW8fD+ayMKlnarD9BZrFJK56z
crkE5yACbUcIN2dr99ZBpGAug63P6qg6wHVABSl703IkwMTj8e/0A0FaxI4Yd9pa
0bXS2FVKeLpUCEnyiqqBbfPUfG5WeomAdcpEsRHpfGfVG8ndO7QB5dITYnI4MvAu
EjG8m91ST0DhDnspUEWzSLhi2U7QeFDGjsTXFpBUHj2KmzbQRCmqAFTE4rT89wPC
On1jltwvb9F4bnxy1kAXRfR04PZ7JdNTmN16LUYX90Qxe4CZetnwopCRjeiad7PM
6KirGZRDotFVyS8TZN5ej8RSpckICnGqtmUZTCSXoGKo15cLSqh7h9/JBF4yjPJc
Q+zCJLQIRI8ZH41Q8lqdsneAirRVvjrg6VHvFe6rDJkhMgX5JjjLFgCNygw8Jwz4
fVMeqdSGVn4HkXLCCDer4icgbgHVPd9Fqopa/SLZc1R4CI7Y+tMsukONz3vpOeWM
EodvN+lOo0YqxAn2l9ExLI3+jG/kpA5TK8sZ5iP88VEUqtiISU4MY+Lit1nPsAdp
Og+nmCxUeW9hcgAADll6zv/Ht3FehP45L75sM/kKD4D3vP66b5fxZD1nDZi9zhVc
AqeAvmm/MTgW8BTJwsxar/6ctPWaXgJA/aIliQtqUjeGzY19zaoDNeo2q8BrS50z
Qs9C4EIE90q/BOI2geBds0/OKSGszw9Jrsli3qdANKTKtx5XFEsaYZDmysz5FBeM
GWw9STl04NO2yL43PZE+uO12qbRhnM7Jyt2Cn7qQR0jIdMKgf0XLgymrDWSVphNM
PqIP/2GnQX0RkqS+sftVlpQPiyn7jP7OOeYaT3T/alDxo4iGpawzAvHEvVo5S1Kr
YQSEAebHDROBiPNHKqxnZKeD96ztX8YllwlTNjpIpoRqE8fuqBuFelu5RFXexwQb
eCQyzbuM7tKJWvVi20ZJmBxZgmhkMEQrgmxqN38VzN1IMSCiez4j7QrjKVDned8R
cjuPzLCP9eRjlvbG85sxt5PbBFUWIN4YXM7NC4roJRmLPSDJD1GBAJBZTSXd2QbY
CcMziJyIrj4r0W+d0ui8QbnNFsleXjUBPYi+Q2Tt4V6erdd+LBSOoQM0zvycHU6t
wZfnJzVtCXBUh+d45bxktlkacJTcU3esiWKMdyAxgmKwbUuUaFi4WxHSle024XRB
kjAODm4blvXY9p0nck9CposKQnFNiPJJKJpAq7jUiDRAUSMWPARgbsgU6avx04sT
PMEkFHFXbVMopou8ZSFu85U+1d2FbtDP5adwNEaln1WWDTWcestCT3zMIe58xxfF
SwKq6hEkK9JsiQ9LeaULrfmfM4h0GrSx94XfQG9yenkreSIPAOkfJCHpGFJugKKq
359ExWHU4+zTxFEuu01VQl6uFNqbQV0KU2wOjfrAlzioMOhRVaU3PGZydrCZRPMS
ubejDzMG67PVj0zcuD62RxHZ1/kRN8qHHTTBMUSI9GCysAqacQRdU+MZ8l1DkUZD
ONFotCEb+N2qt8MwElLHql2YztFL+LqzmykemMg8DG588I6SRAWSmDGfJ9Lq7iiJ
Il4rFJ1GNBil+21y7VzfwgDdcN1H74MQvmDtk3k4Sd7v7/dPrH3DcCI/zwcPIpu8
e1bwL445SkU1XofeSGkSHa8vGGaeTQKkYq3cladJHYXg/E4wiJcQ4gQrXFfG7tP2
+yk/se1EsPiKuZ+VUrV1e7XI2YYg6hLN6gFY3qz8tjMdKz2jv7YwD7dpjcZr1j8e
L58kvXYCoc2KSGdUb0kK5D9kkTw3BmycasJqg7zQ372DuMX26pF7AAwpq9YjSiRd
WMAheMcsfgA0CgRzKHF72X9vmNUBbtQNzp3WeRzmff+LWW98CbG5ZQoHmWoH2v+u
O1QslG22L7jNtrhdfxmGfpdR+0QJXjD6dntS4o2JA4WIoVsK5ofdLNDwwjir/T92
bX09i4HY06sr9OIRXkfr/Xb583Vel/OV0o//UgmlPrN18hS8nQalxcMd6Rzt5XoA
VqvzhPo1sL2McMHqUqSCiQpN0LZUgsz5u6ps1i+dLYHWc5mNGvSPIbJHi7syFDGb
1Xh67CtWx+E35g9TWj6w7vAkNt4D7z58T2E7pdZepKzfETAaYUptlCzPDq46WIxW
vC83PGJD/cKKFPVbENzl/Wb7TSJo9wx3rSJ82gJOMFsom3UEzLDCaiGCiIz1q88e
99YO3V68ccX0cPknQV8n3pMfe/RRBw7ZWtxuOgxyWY4kk4lvWfsTOY4XIqnxNWB+
sXyEWwQybQ4BxLWVmr+JU4WroRtz7nrGLX6yZSrUkmodgKzWiwhso81XPw4ivr6O
urYTh8z1uPHexCmepDUriJ/7MYOjSkr+IxvzEdhpcqOBciYDjWyCy5l8HSKDx8lw
nZpIegDnuWi8FmZd2F6pFQ/eSgv0i0Y1A43vBDyBZe01OUoTZg26btvqDdMNztjw
sOWOdzLFBlT9TMDIgekVTZWf8RbtQOtlzZfAXoIiS529X+t1kMKd2O8PvauLjqYy
GA/uC2Q8lt3BQMcncqi9DKd5ryCTcXQBiZA26A5JsOvhxJR6ih+aY55IwzvgbdRp
2/f3iueWw5cfw0Hxxhw6+0ArTT8K6+wMUu1jUR5no2nRJ9uyauN2Y+kKaJ87Pjh/
2igV3DUKwfcnz1x9LhnKJJYN+jkcR+4re9K9QzNg3fRcyKseiEsQ9slCZIA8hvn6
aNoLVCcLLUWx42CQdR014aJGwIl1VrJexWPG95DJENFNfbsvT1b/E6zJAs5uaKNt
omUGq+Dpj/EieYYkDZ4jUaVj/3ROvONSwqJAZqyeU5T08aK8YO8lFcUxFHYyyhwX
33v8PbZAFc4jLfGmdSzX5QJGiiW4iSGl+IRppeDn498C7aJKaMAxM1RSnw9bugy+
201cXO+2iMJjo0SxFXB8Q3RqHzQN6MqMhtUu+KeOH6yCDTl8ov7w/VFzk6FsMBJh
tC3fp3xZZElqW7pqiouCPGwqsxjvbIPa8F13a95Qd+3wxrZS1eiQkCz9Q6f4Z7lE
GR6+SdQN/qs/mQEtDkN+rvS+V9H0nuZ3LALSEcrqD2eTNVyWzQt7zsfwd0d93dXw
v1Z2FnSRtGLprMjnAeAZJT7CEQJmimjepgU9xkyeyI3dHd0WZo9TsrPj5gGg8roW
WUt1I2I0da4FuV+Abb/wkmJH5poBKWHgr3mZ0n17BuGp1m5mDlR9/D4ZHbhGDv96
vo9sxX2pdlQ7/UuT+kQOrsftM8ctPt8FI+pR+kGK9KRM+GiZfywyMRtByBTOCDsA
2jAf53m+ZqfPBL6d4Jcw4xiNmQQQne2wiqxMfF+JbcIMBPKEsnhzj3N4KKnerBfZ
R547XUT0lYlhRmR4EBqSyUxplgHEkNHCdQLunqpnPvpKoRkUE5itIXBX+Ci2y+M4
cEU4/VnjpHjfWPbZkM+9DLDXXr8ZGCPJsFMTuuVBD3zkFqcP8oBkMW0QCAj4mnoo
TJV4/57DSYhliWrPJpVhTP+wsZneWBpYn+o1b/CUXDTKDdeh02xmOjQEEETXTn0F
K3cSAbkuyCVyJWoYCeLCdcfJ3dJGmjokuivpX9+jrtNQWuUGJXMt9RMPSJCa7Y06
ZadN2a3No3Llzt4cS1YN3Vzoze/ZM4EWI7svceJhDeqbIM0vXT/V+2wQGKkIeMV/
NKTbtu5WHArCNrhdsuZjbAAV5gad0kq/ZSMYguJPu7aeJXK5npU/AP8RaTWkU9Bg
ttSsYgf174QMVP6IqSbcXcZohPWSTWHk4/vF12/gItm4nefO4GG0Fw7OHLU59jyX
HN6JNg+3WcnElPCynlVYz45PKyahSlkA1xUCaTuMZQbGE3gZfyExPOoNsDpyYe3y
fcHUS+Rp+SUCOCMi1N46W0BP69YfNeMU4CbdASGPopbcff6U4V6P37i+SWB+HJ/m
PXbzbqvQ2V7S0EeBS7oTLR8nYx1nhtTARYH7XF5HcJ1GJoUJdtGYhnhacbfsNzbQ
U7tbSd5rRHCLsDfa2/wLNQiB1FshOXDadynwfvkS0sIsho8KbaRK0DqqBsHFr+JZ
++hojEbUzS55JRXKAYZjS+wXgNqRU3ZPEs7yt4iqe2AZA7Hys8GhuuV5NFWqup7J
vZyI0xdkc51DItA9g/P4RAVBJPvZSsnGxw8SboiIVrckgkl/WMUFtAAOMPnNjbpl
xom9J6FZ/j+Y9EPGLM5564p1mwGU7fa8zfx4DaPgN7MGiVK3IYC5gByt+CZ48PJF
5vFTNNn5gfE9mYSfDoGJn5+TzhBZjpFgPBcppp1TqplA63Xmfy/xHp0SQxrHuC5a
Cy3RJ0/QdSnlkWJU7d7OW82w+kIBxy09yfL5O75ggucDIWtGBVaypjwYAEASmTIR
yySv799yJvKT/f8+3rD1FwR1u5Tw0Or1ZiAMPW3w7LWJKnlhTcyovEiolLnWYtRW
9fd3NIb5vDOoUqMZYQvio6KtN5A+8vmdO7P7laJqj7z2LGBEk0WFhHLyxZG6+VvD
9rx4UI17P0/iYUwqtEFGXzkoOnssw6xA5bZ3A8uoQ2GhNSVfwJ+K2720ztqJRx2D
EiTj8/R8zlW+NmPGLgUU9jhIexnJHajEHAtgzKdnfTa0nPJY6WTKcYelfV4QyT1U
OksSHnSeA/rIRwOWqMcqjG51PcWoKSFM5tb6ljCzbxHU02XiBPgsNRhc5BKgoMCH
I68w/5UZyqnjFFgzDAN0fskVYf6n8TH1ucMksUOrFBBu00NZMUbqFBchXJ9FpU/p
mMAXCQisX1X4usUN60TNM17ocLHm8NuvW1unFhxvCk6CoDFU4bCp/Dd3dh76I2yq
QPQINfa2+tO/eJUXqK6zGnLrTVwByNTNsKRg8M8NVBIem1EaDjZzQ6F3COp2euwJ
shbJwxx9EXEkuK2r9j22QaOjdl0AsFigboYEujehW8kDLxN7xWHiX2vfcmRGCjSX
wdAhmX4+/AC6H+ICBvFW+tbdr6U8Yc30WHPfJTt4dRzXg+aDq5BDxo5L5Gk8rxZk
Kpfo6Iei4JUNc1yk5unvAAOrCQ6nzloVS5Y/x89lK7Q3I2cYV6my+m7cYpOE+xk9
I+yII42ehQ3EafU73Qhg2NNIT9EGkS3T0w5dTKCbob7ZnVYs8Fut9vTTpVEuhkza
zgTzH4Wv+6bSzWIceelcLpipntOrAEgDGlXIHXexxpYruP1B9qc4j0pz90FjtzaW
9sCox4Qkk8vPZqrfC6iR1iY4U+ijiJoBDtxSX4xR084MzvsTw1N8hioowhg7KZuM
dBsQb8q/tKTCbCqO2vCpYh8HYKq9bYCajW/x99W0nkuGPqE494SLBJh6pt34TckC
rJ9u3MCb1yvakO39NQyYTeNPXiZYRG21Q3KZ9qMl6DC3dU/dXxY2eHcoRhgxZXnV
arh19GE3S+8QBKlWGENVZQsqhXCgFswfEHs2C4VUWFiI2bYsuoQWTCFqSnxzhEfV
WIACaaN22W3WdnOATswMgS3UnLGvGNQVnT0Jw4r0z2iJX5hkmionm1uh4RN92Qf9
jJifuYsGEGIVniKZcv++0Ru3hwKgnhcQLhLY0Vso3c7Ses5ZRhluUpOt95cWiWx+
+ki+iw2YJwAeqXjDDfZ+mUWLqNAGL6uA5ZfWKhcPQ+EqXPg2sWiYtOqn8QrSa8nx
Rsel8YRvWPEEtS4fglbR2A==
`protect end_protected