`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2320 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
XVHVS6SW8Hb+XzH/poMIoE+OaGYBc5u2Vk4E/WRKpQnpl8WTv+KLULq+sJkjEQWP
IcUrCW/bU3CFMKIjgi0F6D2OweMJ9NHAGxnaMUTJvahND5P/PGtAXq3SXhIlWs/0
nDWiOYntU8Zlv/474MjVI9U5WLqHGJsKhgLhTx7z6YoQrYJvcBKw8JWMcTxsFJdp
1GUZiC2/P79xc/Ie5BfXzDlUk53A97KLLk2aVegNvaVFAoJ9OOl/JBQLbq/QkdaP
v6VCLjc14tIatR5sIGBtIICSptgJeVn5ZRAa5P7nyFeeGEEjMva9OyLOEy8wlTkX
hiuVmPg4Z+spmTCUJJXlWw73OVrn30jLTgfwwtr0JwDshunaMaJdKi6ZdpYPDlH4
YppPwuej176e/nSTDB2CJ/eCIrPEDYXguTYuxPqZ/C8y2J6w8RSciwVptENK7+VW
BfRJ0092wj6ceMbSqbcOsB4LgQ7Hz6Yk/kZHV8PucSlWEH7Cr7+Q/09mRqzMRRT+
uRrNo+SToDUH2A5xN505WK+wsuXyUPp5QFmIekIqlZ4e4vpVmjpw1v2F/PD9mwFc
czXTUFaOrrl7RrFKk4oFQDRdd3Jvi/XbNUa/u2KImPyN9VVRmXk8lxFcp5/8gxeG
4joCOAm4WjEvnyqJ83NXjBjs/sleOJIXbRaEAarpII65LZQV2JOQanEVD6yyqvdr
qWBNSUENJ6bjqZVD/95QbAM882OxctK+unsQ/Zb6QGYXwi6oYLi2wt7pECEp7w1e
I6d8WmK+D1fzjoyF08rotPgT7YXY2oV0wHAWCE6/3XqVMhHkQcM39iSIIYO4oXP2
n9wEAoGqOkyo9PmJghQE55j53VlaMYuJgj27u8KWfKhFV81i40FHnKKaMxQt6tq1
d7+ItwsO2AQ+6r2htN9MHUl7uVvt23LseVZtR/Xvuq+kTyWTyCO3ci3l65tvKDF9
w0JO5ePgy4H99+hLaQbxECnWili4731Hh6bNfSmUTHeT7uClW70cTOnDJFur3NL3
jnq4MH8jpgjGBdPCdfeyDW8pdr3bFvVOhxL46ED6Go5U2BnnOqk6Okxj3cPbmPEw
aXYTY1b0jjCtZG+kg9gUm+f9El/7C8K3G4tCdwGGGOnUUCAITLY6qqpStjfazSiR
1PNN6/qKqKeLHmeRvn8K3v6Qj+JG575WAaoQRNMbqFaqsSBYXR4LcnwJstDgAqQh
nqh/VVAqavBEzzTeq38bNtotu30JUlAbJiLCuaUWZ0/sXf9SEIODXJLeRdaoLPms
faT+DtPfJxW0JnC9s3QtrGYzJ1EJ71mbbim8M8rPAD99/h8UdfondsKk7lJMGP9k
rESlQN9E9uTNikChd1ZxZRWZUoOygCOwfRijdAHKkENhWLF0sT1AioO5GDqE67PD
iS8DwHgbNV702/dDsnYfsTgW+8sM3a3wqCzaWOwr/+4005MY2qmiKP9RZaYhNIN5
OJgDIrK6+v0sp9nG45ndb4PAaWZ5eC7ygvd/6a8IQGcCwwUSSS2aFrLK0A2pwnL2
CgsHUD/JxcHMuI+eapF+prRKGLIZgex8D7DVr6QXLnpITBBYm/UzYiM5ey9ws35I
UXcLRbavUhSyWC5By8De5aWVAGF1wWzAVw9VAVm6gDNKAU35YkTb9VyxWEphE/5k
Sw7emapaVbFDYoIMdWB5yNRHSQD11uthXsNdqu5L4Bx0mkkQsUhie66uZbFsbqgE
m3zeKFc0UKObxAGkOvaSNUj5PRW8CkZCeKzQPCa+JC992NNLq/0XhWNuPOe3WnNz
7eBJHdWk6hpcAWnPM8a3iHmzhHi1XasARayHDYPZfYzukXGnrjzpfvJJMvy3JwjN
YwCMMcrUarg/8AZHBw2FdTWUKVi7xynWqxT48Ohakh1suKKOXq36eSNttBfSfBPp
UdvYmZpZS1iIemRLg0zzaDylP5B4xc1rPJ877O4FxtlCdH/sS1eAeOLyNXXFxF8/
D10QXOeQCdBkQmaY34WH24dYJJ15bf7x6ngH2hDvzc49s+72iU6ByFi3DKxcGs7R
g6WEzyRegqFgZO0Kmjrm+FqVz7a01yNQsufag5Xvo0PY2ptHOWvcO2HvbMQeMAlx
rTP9JFrZQVbokGmp6wjLh5UyXwDfKQV9VEr6naoSEdNmTzvErGStkxjy8goAEd1U
T099aebGyGIp1EkNEp5Z+/mN2eZPVEgIVID7PBkw8vcxffn97K9waGpScOgeHshh
szCfBtwMcwomYVW1Y5a5FpOl4lyABvn3nJXWW5VVP3MPltH0w6HMqFBJ88y8C4U4
ilGNIySoRgmSHGtCc+OgMDC3pQsoOXCH/2+ylDiedLXzn9HLl+2cQCTvJIlrsqts
uz0K9OP3D/IplmQ27QJ+1OXwPmhbiX+oSTOt0M/+/NLkbeWw5keaXGuWiJ+bdYBi
Ikw0fnESkieyLtq2rX78qVE62gw/JfOh9UDQg2vRc+xc6opkElwm6EvRqJ7gre/k
9XCx/DuyRzLcjCeBsREKODbUOletVH8Dsyjl8OKItSxVvK7cq41aplJTE7hVF4OO
pS4aor4Car/4tHG1c/ESXbUkPqOXm0hWfqdYk0WeQib+BNaVlyZPhTnnjOvDwatP
brMs2NzvnsRkHpuN8mcv6JJlpqZ48AMy0deTQIT5uNAbGD4ZY7egwwLmIg6sQOip
s0VSqaTNiAIFu6kEME8GRyi/5dGCPctkNhF+E1vuHPM/HCMHkKyCfAIphyjlfqab
kGU0mKVJ8eiZBeApb5NsEQ89H770FPpYAYvOdMp7tQqElWYKMfvHrNo6Y2zfhND8
wiXbp721GGVQZ3rCy7/FVtyS8J7XBgb2V80WrWwKea+9Y20o/0dkxB3h5kTLPMEa
uLaWavyvw+rR86rWL//rbNZF6LLGRxH1JbjMt4SJXn7pOrIiRfqetFjaPh6zVBDS
YjG/q7MBmwuBOnYTIw8MrA==
`protect end_protected