`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7EpPiMK+Qq1h7p6l90CUpAjN
g0iC6fuMZ5J8rgquZavA9P+HxYrPQ1PvXp00D2el5eG8+xbP9hxsyY8LH+tVrnCt
XVMZSfm/5bOvsaapYhQuit9qRZ59O0DdFAm3LB8bVG7tFe2frg5oe4fuy7NCMtsV
nO58f6vQN8oX5oavuypVFrZhhlVYWPql4sVmryeDQayK9sHJpRx0ixfNobiMteTi
nIeaQYcCAnWV/xCU9sdB8xzBkFAKmamH3sriujIJTRNjt1hnJSTZpJZtLgkdO/+g
l78q7EV0QJjVO+lyhLM+yvzHIkiXIW+Qw1xHaql53gBy6rdIb03CHVpyMRuyL8s/
Ys1H2AGG18dmk2x6k9VhN3IJ7iXG5ZtSMsbP4/9qxi/Yf0QqGNooEv/a8LBhVwbL
5n29NY9Y7SXAlZFV7pqfTV5n5ObR6J/dKMp9ecgnZpJKftKl8V46GTjSQfpOE4/q
1LdYUg1EyoOW5EVZB2a+3inpTJl/3+WCAfclLZexIlJ/bSaqxmnOppmxC6UCBwIy
h0Rin3chC8sUQ9yw3sCj3OWUeWTKwfnv0O4KSepitbxrrwPIOZHw5ozNylHDGoHK
puhwZ43V7hq66GuSKi5serfh5d0iKr9Wv9esB8JMduWe52IhRCnalZJwk5XF1ZG/
b5mX4++zbARsZOUULvy86uC3EgKMlI1PXvcBSfknex4vu0ufzfuaq5RoCOF4jij3
SKHfYrNuf9/vTASKCKmIXQksYl4yNd8/4VLgNT4wKSdJUVCXnji+7HMZHefgHlCP
lepP+MkwkqymwmhuFpzzOzdb+zpmUzM1jvAhqxY6iKMn2WaKWKz7AnkYtfXHQCU2
EVbHlby0t9FMBMVV3620M7PslOrfC2bjEm79BYTy1O95s5GkFgqfIMIEfu88YlFw
I7mOZQyW3MutsfEBDgrguuf3rUJ+oJZaEwaXlyRDOVbjKXoO6IBpJWSr2Mjgj1bX
sJdfNAMQ0B3QILzGB8IHJNXK9r/5pY94ZnD6sj3345mfB/O4CS+Y7woEzpbPkaDz
noZ8MulHWZWF7qRfOVoz+Y5cxrzYY/KxLba94h1CtTag2JHOHmq/NucCHOLc7zS9
J1LGGC8lXf5cbMJtlUQXxoutamMedJFSGbIIVc39gHUqG0su836of2mIIv2Ysg+r
ZQ5qylnBj8wofa/ebq+yhsRhZm/FUggq4rxZ4yYqHiqVQ0k5wN6cVFhiWCOdkilE
PGmpOayHrYET2CuAx6taKWrnYY7HdgkqjHEsuXvS2pLDgOV178kidbeyrwZlP2eN
FVvA26sVKe2AFe2aWQ9imybVPDVoGxVGEaiBVjzjgARqvspXNQ7wnh1MVhXaFGmo
o4k+Z3Em2O7Rl89vHbrPWvVXvoOyz/8baPwifN21sFEMGqybUJpxlUfPRdjr9IAQ
+b2s8qsr94fpHufMIdVRCpKILcwOWm9BMikVP6sAjkRn+wPIfO/Y16I4qhEC2SQ2
vEdyA53b7HWA/F1qgmzMI/zQeF6pJ+wKzLiZOLclRkMBZ6TZwBwIrIDFoUzW9R3D
SCztO3OMyJOoT/oR/JWuobhKfKEmND0F74RtAni2fnWg+Wafc8rPCVQ9dgzJfD98
TmC3NeGUCAbARC5ha/EC40QYxLYWYPVIEI5bPJ15bCoVNloMGvkqT9xX81MMVJLk
OJM1rWwr4vRLDWGheKMX55BL9J0zme5W+BpbD88uPjqK6ItDdOC5qn5NCtABrwUc
shUZYXcak/t0RxCgJ5iCgdWRowl7XTja5HYoVawYZsUD9k9QZ4hZiOUaq6KJ73Nf
2uDy4KyGzWr3Ck86k24OYraS0oFpXpS8NopGthcjvUB9/ZR6UBx35S/Bp7Ommzgy
W1vLi3DcFVTAkOcj3XISVosvrO414M/umwf+BM8iiVHn7rglD/DJd774wVM5GaFY
rV6qD33oxt3SjTkZTpeJcG5VwwihIjmI59OjGeyCSV76GbZz2Cn58gid0+cjL1nV
jzZksnz9qgJsa1V7SSFLR7QkYyGMCi2wbG4qxoOk81QMQNpt6toz9iT/hkVgUKuD
X49wT3SgevTy2F8PWBtUGAyZfa8jHHJ2qy5vrnnI+SIX/X8EnOBhh728Aaqrwlgt
Hh8ml+52ql3zmfvkUyhfLXLFhkmtfvuDx5I9bcFL9UxIgAOQcVuXGWYKOFJbAk0G
v1mls0a/Nr7WMn2YvCSfsipcKWN4t/pedz9z25IsIDkg3r1x+8ks8gevFjOPg88U
dUpgOJZNKlRPZOennngX+3d61odNG/zDQgzVWKaBXsZ2/TsHQY9Dk1I3AxCNShY8
zd8Oh4XWkxPlp9jPEqYfwA4zDPWQKEwuGxFnSCcIJIDRNrUGb8DRAtMUGc27wROE
sqr6IMMnq9BUYxmoHw/KL4Xat/JPIJRm+qq1ZALDxkaQH+yQDLZLtBiRvCnirB9c
A+BhjyHv+k9B7cI/qNb3fibVdyurRZDaai2Thn9fbfOobmLl3zNSb7ywdIBalhXI
T0NsfNbo+15Zj7KJOXRUM4BcjRMPZISPI23vea79aif5FBPQyda6DpZm8QkXpnn+
OugM9B2LmYCo5lCVe6ejJhbQl/FEIjT4DvSybcQnAPmdlfUd10n5179VDIALr5fw
FXP87txbe0vslWxCY57r0WbKpMDhnVeEf+vAZOh4yuCJQqJnQ3SywTcMrQnOlvuT
wlW4mkL9BsHQTflLmNBs3DGERsUTdUJfPdHGzSJh9vTSyKhgN0t+hKBVXK//yehN
K1EfG7A+05rdHIjBy/2hfCxBBmUslh+KayLJxFFFzo086K+FkbJ28zr4+C3+iTAg
uJ/5J2Ha25hkjEtkMv41WdbuVljt7EJKUeXEMmIh0+p57bErD395OVIgfWp0T4qJ
Tre3nYRVdlfODdSYVPhgbJ/lWMADn3f9Vce/5nUZML/egohiOKP9GM2gGtP34jaR
XefM2wwngnXYJdtSGy4Pyb+VGJ7hcP/4nuXbKqxa9ZnzMFq9kJ6IGRmukqTp+HRF
iXxHKHIfhMFZyRtAgrJVJha/NoWTwCqe7ve+hexrYD2elFMqAGRx2RjmVU5SeN6Z
qj6b4Wy7adlo7sFsm0l8ndEWW/R7JIi7LNt3TFUAuPM7OBdutjnd1HKw4hQOZ081
vj5JO2fj9unLqhwK9/FqpqUwl25LD7i7Meqdx0EsBvLBfTb59PbwdJFFuJdzs639
4WNzpk/ed9/BgPWrStPQTCh9azQ+fAHqEiJjAip7y+YbsFiGBPwUL55xxTWaI8dI
t0rNGG2IPUJt0OW3vS4eikI1swMpYZ/xKs1t8U7Hy8jD2qx/VtOYT4qf4sGUb4Ke
1V9M1Y4btc1omEuJxweavLBZ6D3PNkzX0IHZVgNX2q3QdXGi8IU61zKMSH7zYxvM
XXl60+A3WIS5dCSKFMY3fbO2qlrJKR/WKc2yGK0nRqSHm6KjBGU+3vja3Mr9kTor
ck4CZph0iq+0dzrJayVp+dCgpShsau8tAT3usQhZ1MiAwuIIzKCiqeUl3sQXv9zo
CfIQC2NLYkVrrcsfhdvb2X9PWYjZ5NQG/3l6eIfOawqIMClGw8EpjnPJUsei0wYC
xfpL7hiOxd0le19MwSVI7IQ77Lw05Y0Id/BYhPxNvnmW3gEoRkzZgMLKVgZPWihI
hV1MacKERGzz2qY5YIi5gV36JHDUsHW2wWqEv1r7YVuAvKwddclm+AUaxgW0BKNN
ZSTmd6+JqwOEf4F6evHlD8j8qgtDl+O7VQlQ4PguiGWYLQ4IPgHOixCaLiTX7wls
wI1sUz0c8po8fnLlk4+GwEgzxpz7eHcRxdP3otDgK1cXgVol+M7asOr7oKqQTbY1
LrneNTroudHFrQC/fr1bpm/+//uG6ZgFuKKmUMs6rYZ9sdbXQ8jdVyHsPySvrc5Q
hZdRT5FHQF76D811C4zcxgu8qH7LF09HyeEBue5B7+/IV7l2jwKvAhyMrIH90mPO
qSOSffd/B48BkfTNIzoDOIOuaNYSqDCpCgwjjtaapNoR1TbcZWjsDwsl4dAwQ29/
H6T/lMMmKJF6VG/SOqrbo9BbVSWMyAcTBsXV6X1a0V4xDK3BqyrdpwKeZNYULwnf
a5mzOYZIJ+mpr99nUdTNLYC1KDoUuo+v3ZFUz/ykiFEhQYLV4FOE3PuR5j+IgkgB
+DZ5QigfzVIUpLMkVBLt5y1x1HRc0qU53YZHEewIP2uG7hRB9Sst0IH160qmekis
XaF6vSOgvhPUeq4v1Ik/i0aYssuu3A+j8W3LTuVo9hr7yxYAiYlnMJHV4VN3gRNt
efh2m2tlTyT9xTDv4xO/8ZH8cPlADbBhiVOh05eCfR0lUspunleLLjDcDqIvXWho
JLW4DrX0OoWpKbesseumbqkMVGdC3TY0T4WJfzi407ddU4TZHgsOlwvhOrjU9RIb
tGrtVivZbm7aOwrD9l6R+fnxAws2HoJE03XE/UtKrtuCzaDeZfq4vKS1lE8IaVqO
4W3SU5UhgO894fKth+RnLkF5NSy3zDB1W9QNpxrUkMBLztxPOtxSmHqIQQBFvb2V
cHcBuxtPprg5EN5FmCcq0soKDQEJCBqeftPTdNVOpM+Pjasq2NsEIBcjlA3WW8a8
C7i5ieteXrs3IYjL2sfgwFaqqNSruTzueZoe+kQHxcHpQFpFQFgpBWL9YzoS8ECy
eUwUBoeCYXVV4DTJ2h1IexmR2Hbi18o+hbeFsRYZlOCZJKxG9ypWw69IrY1BQIC3
PYyr6xvjHeTHPAVq4B+agHSoZ5IcbQajX9Xa5IXbyKWkTsS2hYH2Nuhwq97Rv/nb
yJTr8SyHvHTaynA4KElJZU/d+OoAAbtHQFVJVYLGCs5zuhBsLhmEo1BfWcbBIOwo
rOe98pTqxbIk+Z2O1pFpUguY6LzyRitxqKqMHlJvjsJoIIQ+rPRChou00DaDfVHF
C2Yj6j8sJEAYQ8o4nH22X1tLDwOig8CYKNodfGIZPqP0IIsF5IjOzPRJTUF/XrE4
2cAKidP6HNSNXrwGbR0RXXOvZ8HGHizLEVB+34oZ/FZTSJ4IFSP/ooKmtCFp7RVm
asWGj46RG4bki7bRoSRuhs4POi/4i3loi94glEWPyLCqogJPiK05nXQadGuce5iv
VqQzuGEbQtiFeRmtSL9ZSwentx0eD82tEV1xelehOZDxgH0F6UAtehEnL0s0MJBn
zFUK6JvYFEd978z0fJgrrNlv/KOKzfl8uM0A9eeNNoitlfxPJ447WMB2IrPToMpW
FN06R51kK8rKRRACEqlHYaaKLQdKCkttR5GLoutjXaCALOJIl433qlOR0/oKF88t
RGD6f4Xd0oeChNe5wA5Fo516wsNJnw9UlasnTeEMdYk/kUsXcG3hrdWW4IqHzWfh
b9ks1hfXaV4h/5f/dxEqf00OK+QRlTJRkLU6NnnyWSqAbST7gP6gWyRSOpzm1V0T
h+EvZ1FUMFyLHCsYdchU55N0er0fkyEAb+gLIbIBsvKpggFk6FkM+bSOJcC0cCrH
G0JdcjiVhWkGTdWMNUcouW5n2iOfZAnMOE68FdcMmMwYnzaZ2P+A5Hrf6MdAWyE7
diio3UUqSAo2XTBS99c9Ky6M3rkrlD+AGljTxjGe246CiDBQ85c4lgzXRK94RIKI
pPJaW7W2N/0ih9M5UYy9O0FZUSy2E3f9/2LA0HkyY6tuXTG8V6wKW5A6Qz2daFH8
IQz1Pbytt85vpnesIIDm8zjCRaU+hV9yBc0tMBMRr4TZ536Q10+P7C6XtCNIKgEO
32I2mIWelCR7j5mNedbeW4BqpTstjYxmwnMIzt6+wcxGLTZHPp/ma5ltGJGqIvGt
dJjBcy1sYO/9OyvbyrTaSPvINa96Kis6JExl4TZ6xnXCSoA8PuhK4gLdFf/kq8lo
xSTE0r+qyqRsMqEiUYFvF/ln+S9daT+1Tq61v7UkDMHaOIm8y1iE/khVvNWrIpKb
lVpivI9B/Zd+Agn5ID3jpb6lxHit+TpZNbsns0m6wzk6KKDHXUeq7079g/IJCqyn
vX3b47g8qvBhg4tnjXjd6IzItHgZpshUFNIQq11y+FVIuMHmcueFflwwicgooG5h
2/p8fNcKeFFZIkptYImin3O8+5UtYgLwSJJ8k/zEMbH6IoQX9rHM7NkX/IEimCcG
w8I7/QaZa9YEdaEqVxYutwqZAF6FWl9m9g8j8RE9l+rBwu4N1ULfPX2QS/eB2gUl
2WlunZwFLTWixGrLecen1fRSvNqtIl8n45Fh/s4dEhsSQhmRtzuSv7W/Zv0dy+Q6
vAjZieMXFLZ+HBDdL743uXGIQuu+MTfSnZxbZ74btzUwjRUWi9SxlVGTszMmau2f
4AjmsWLgZgbnpUsNPgPe4a4HqdL5bKiMEgOGpAFjMaQw5SyRQ92IxZHwTWCLfu3V
WriuQhWtZ6x5/GDXmIQdz2XMbdIODIYmYZYBrqC1LK2tz49ZzpEvVMsySSAiIq/2
HMV7OTqusN9k+NWhbqe/JbkaKt2LXu5sGhdDnYd8tySLRVByGWrZucimJldijlGT
TN506bPEJMWgu3xIjrUWLUw8PVsq2jvbXabSxqAHQ8k9WUVJfKAu0TaqiZeycyt1
DYERZ2D9nVCDeW2ZnGmcpPLfv+eRd2b2BhDWTUg8eIB98yVmumP0hdmoYx6+R8xn
PDyAVGdwkiYjVTyoBihX1h6TS+GSPFWuUcu2RWAVFt756GgvkYlAF2ut/3imLn1G
gWXBGfkqvlsbuuNwqkoIbj2hOLWCrBLkSPnQRou3K5Z0vhWK2sqSpopo/a/2ouy7
1U0lITzIRpZlVSjjCsF5xGSgTTL5go82I9gTnWn2z11VaLH6/bNz+N01g773H6hq
GjTJlmM5hGIFynPrXCa90w6V/8q0CS5Bekdkj+nJVdxr6cxVh/bwSXBT+QQf6v8R
yCnnEI4zJbHNbPPf6TrSQ1Mj0g/SdlTV0U9ubghu0qPcBthQm4TDSCI+cdqHccEw
vrhUQtydf+ujTOANroxsLR+hcyGgcu6mdhhPFMEGq6Y5fn02Zo8ifEmolJorSfZH
Idda20OXiDvhu/P0Y0mRF8Fi7FYyV1SoJ9l4T5MZDgV72jaGwmvPJjFYgdH6fArS
PYr+myYSyZD3uE1jtVucfhIJx/DIQRSOZzripIQ1czJ5hwvIoW+AoR1Vy+Lw5aVF
59fecfh+i4nolyCzSZhhAVdxAh76aDEaAWggqG4uf+1jhmrwSqE0CMQ9SJZnT3jx
RWIogznkhqEm9obWvjuGjC7vwvSOgiPzDozAkNv3Fvbpr1YMB3x1yw5PgssJSKxv
pcEV6i0DFsiRHKaGMBv3OIVJ7lwgq3vfxmdku0m1DY7Sb0tbhzMMOkBA0lwIaQRa
0zzlfyuO6PP3wNaBgKkAnQCBBvTMW8rncH8pul28sEo0h3aHFEjeBNBE3i8LBuLZ
R+f+SfPgGZro89ZeRt+ztorZWj6Mct7QkzrzbSysiKRhMHWNzIut/4uQvGldtNLj
YfCfT0LhDGwh1lEb4NlqEaeHt2qw2IGfA/7g0C19Ps+lARGnLawEwieOtNT8CZAD
mjWpZHO5VUDybDyYUn/gnjaDgGInYqtAxO2lwMfzCfSIBt0gFWgjRVEvjW0vURte
iZnZL3EiUScKh3IFXlbOCSq2EFSH6nJxgx/zbYhMiAbioG9ye0JTNk8nt/Dp7AoN
ntMmFrAIumT6PwwZXfEqA7gwWhdGIvp6PjcQiabAeICQoHBZl0OD2L99CVUV3PFW
yp0z7cxKcIIOcNeobaqx28e0ZcZXiTUXh/bJsJ/qbX7kZbu8FWQVyBdRR+25PXOM
+eJWqk+Jf5Mq04MyBsy2Zi1Gn9bf/0X6HotMGHJkq3gDLCDUFF22HKtr7hoy6tpr
8uU27ZV/KXN3LQpusyHJpg52iDVARWRgclRExSkGt0JaH7Ne2IYVJXB9ct+oXFDe
SPlZJRfLwQicr37f18W4nKrqwjNkqnmpEdDNIEu/qwSxuKpWolgXRPBsvdLJhDSa
j87HhJEjOFSlzcxlz20362qP69iY99NjKrRuhKkLU0c6chM+5r2lpL3HBtJscqxi
6gowHuebF5IA/59eYsFsAgwTD13biSVkdkrWiwrrnmB2V8bSSRcS9OUymPJlB7/S
Iu6acxysFo0bo9IhCX1I9+LTqNRcNYzgusdEmOdM6H2W1tPHi6dT7CJvhYeGI03c
Vswk01YVUxWwpeWgrg2kLBvmZjd9TK1G26TB1uZYF0D6L46Uh2u+d1liubQuGItI
mx0IoLbMtnCYaeECAGizo2A543c9jI/9IAhpfQwtfZfBJ+QuR6vFfZvgko8QyzHz
FYxtfNUzx5AtW/9KrQ4BqKNEolMyCcVCEzhcBoSC0XQV8GnCotoEB7lyvxfoKMza
nclz2m8zkZKiJ1L8gw5Id2A1Z1J18oZeb/qfKn/yfhetI2X56Rkl/5SsG521Z+OQ
p58LqJlO4hgrNMNk9NongKfBkFCWGjelhd1dtXTmCAwGGY2Dx5nhZf8yaT7kP+FI
I5wmo2vSrNjwgzsZ+A6/IqxobeesFp26I0c1b/WQC0r7KpvSAo+2z3qKP+iBY7Oc
Y/cWY/vQVv0z8lAbWNVgD6IMuvLRtal1BjjwetbapiENbFkk+SUEatRDCNNaXe1h
tIZJkHeYukcGcKX3IxKtwmLH73iQuL75ncLjtiFNLcEwcdcnGKvFRoHB7dQ7Oz78
YzFPDa3QQRn5QpE9OILoBlRn3LyfwhowcqPkhyqgLzgI+wE6grdB/MneM9+E9ZgT
i6Zsz9kLWCyhkkrbGMxfzw16N2TSyp+4m5dLoPnUj5RYqdE9Eb6UF1r3u03Lc11C
LNik7m0re4YoYvgLzY5yevTCDdGHkVOSU3qv77EW3vsb3Ph7i3Omk9pdDl3n7OTr
ruaJs8LqkxixXGfqJhRPwlv6uHzGKRKijPpnANbRDTz9mfnEM+h7wut90zvtx2HT
S9p9entiOddfEVhD0Obm3oEEkdQdPtp4F4+HObxkq7Xlqy+pTtr/tkjZ6N/VV0Q/
ZAGczt0hVJ/z5VymH0ZcaN/omcILzVCOcW7ALebpn17KwW19819BRf2ChOd7a5d3
myFwkG0rnJn5TMcKxCu0hMoIl44GksUAsxx0lB5m8mq5XNoL65mOV+sbVEk9SEFa
SNk3yAi+kU61fQMEOjcnWdVviIaLgTI9eO50s42HYlrbF3RRCeY5/h4hemcGVx4l
Zq//hQiEi5ExEEiSv9WiFqELK8RHvgXHbJ2Cob2hj8DFas13+8vtxMbYWpcUJIJI
FcQ2HQYE/ASH4TeRvy25ZrLADCEIlq9U+3G7O0nkpiI1obrjInBcfVHJLLkjDkms
m9AEsE0UPTLF+sfZg5bkt2vES6ofAWytYCK0GlUXXCE/MOTOznQluy74CtA7Lvt3
UnHMvV1t13ePo0XmpfJh5K8nfOamr1E05eyIR7eOpNLXWwGRado3G6/mFWzhRs+E
+eqAYed2RCUt2ydwRjatJMETzJTVUpRLEYxlOLrtevUaEcrLuMMjxpX9dT2Y/nl0
ZkeFiCMVDO+ANRIWKlXxNr5YtBJX+U6uxF5uNwb3iXUBIFJredlVc4MEFoptZDnX
Tpmtiu4lszL5ooisLIw9gC2UwdJNMO0LL009kY6v8rQ8l12gx9fklfWR9Hc+yMXg
2TTGlezukdjgUr2rTZdlz99odDNsDfdQAZPk9dGVLaTU0p5Mk7RlZqSdfQ1K9hOr
g11cxKXf21jCFVmhcByr6QhKhB2ilkqKC7aqgoV56w3YnYdQ64DQOAgGR5+0BF4w
Lmfpi8wTDqDnBpqtjKqlNXxYyVaXqUseKWWDOG8DJx+0dr9XZstFtBEqXGDGokVA
0rhfjVcgpB41NYCRviKOpb1qrqXg+A89pXwcw+ZdoicpYjV2IfPAEaeLSodr3lQd
22QC2sSbZzbPAYQPJ+EOX4AHRU9GqVSRnACGSWMFNZXvEBvjDc5C5aIFgEUZevYj
KyvoCu2MjfJgMEMuBNSH/YVvJsdn5T3YMC9qdl7Q4HHc2Mw4z+F5OGPmbQ8qslXu
omGNEVVpb8ZiE2Kt1gp3R1KiVDhIIzo7cOYwO5vZ04OlTxK03Ap9Zhga5LNLjFPy
IV1pBuyfyIPK+Wi3bihgHeuHbBwh335ci8VIYWSaKhND/yrfYnNVMN840kAcd48S
0bovywUU2HIBCuui7Y/uB/uF0dZBWrK8LAR3asnVjS+0rPldkAkL2923sPgRwuYv
VhR23he4CVX7FH0ICVMUbjKfKxpDUxgJ776lhDPtb2C0vUnqJdyCY84i4hADvYiE
bDwYfZ2qfSEj/jql2ltM8NX/uFNNws1GgVw95kOlidXmhXT6xWrVVrFvVmlPLGKB
sPjetUUY+ugEuiHMojA27+WcVbEIClCEbL1ug0B1KqY8IkBlNQLfaBGXV7aqa9kU
3HXWfuVCwgVdveLu2lHPuJrv/q0wM4wUyHOWrcKlM2ykiKP552M22k4GglBW+IRT
txprnp4FJaPjP3q8cFxTiwBCz/ASvzae8i64lttwdB8cRcCU3YwKoFL+f6J+wz+c
HL51dymJeqp6k2bPrfVdvRPcvJD1meSNJcQDLiqPpbR/9uvkvxPswqorVwLCGeeK
GHYqCAVL8jnmrSf2KVaOTcnBKY4+Fljb+4nprh8d7Jm68yvpBYWsJP1mXz2v7qqk
YxRFKMCri/uo4cofm5SKFdGn864Xf22kFXVrRHIAk+R/PmeGlL5Y/wp/1lFhby8i
ugzm5wweUDKuzwhfIwusqNq5n9ZwdQJeqYaAtXX9n8VExDgVbS/yPJLo0g4L+8CT
j8wrJZLGNpFTk2ABXSZAZeMwoPD1YpXUvvVxrTuHchKH3KadwhkrVtCHlA09/XDP
IzGf4JkL6OKis09KqiqaDlO8yazx9zdYZP5LI1nMEg9NMzt2ypngEkkG/MYrcNJC
sdCdfCH5+HEnuKYIv4275pfnfXlPM0dai03S5LBywEVukhnsplorEnfTLYhoqA3k
pYwLJepXsKz/u/ZpKzq3aNbJTIFICUatjtZiLgG/azwsUFsAHvSEHsYLM8cu6OlF
/nFCn7oFJKd4n61dMNO2mYh1r40HWlKurEb+fCpwvpKUvYnWJxcUkfYGxVXzk3Nf
tUQVzD9QLquNN13FwmdWDingjW1Wi1GZoTV8kxq7Xb66faHEGVDUCuZS8nqzCeHY
IChXqor6GgSp0KohZmxmOIOapktrjwnRPezdxbWpSsUjqn20Eq5H8TcRDBBg9e05
r+0n1kKMVydl6YeXlaAi+bgKe8sI2fzENHJwEO6LibyWADUkhfGYxB0iKQnriOJQ
/iIbk9qLYM+5B/47r58seppYFcJkVogGHly+BHzxF1fIPOWkdC7JhDzpy9KGPVuP
gxMw7H3YmYhunolibX9LWmcTvLV/kINBiDPHXOcgK/1ou+C/MTZbdXpWKqN0Pko4
sNBPDurjrSjPGM1Sa8zSnRjHce4bg9ESNJ0INAd1vtHBrGxvNKmD7uieGrqBocKb
wZ6eeDx9Xc82s+bnop+Qs+HfU7dLVqG4Oa3fD51VPYIESw1t45YrvZvsO49Eo2Sc
ESeKqmZmNYG9RC6wzvWdhe7JT18znk6WhgsZ3SG4kEiWi2NoEhJL40xYnZbSL37u
7X5dI35r1maJBCH7oxmzfWIDmrdylCMJT/AyDYx698ovWn1iSbvpDzeO+UK7zGal
v8wK/39L6vb82P8LwtFHCh/l/nXMBDPz/22kCa5JfQiC2Q+vQ9WAmkP9iuvEfq20
sBDQNHu+CiQaIIy4NGz7OXUVn/eisWLsqWi3W4veejP9GD1ieCPOAnC03dCffMBF
VTKdsj9KHS+PdaOv2r2xN33qQ5XKnZJu5k/XVPpSjEqRUCiK0KtsPac2kWLdUrCB
6qbUdPOtoad1XLPaWoBEkshHXGA560dL+0gyhkawMJRGG9BEXCrr8eqFUi+KiLHJ
VTdLdY9+lbRJA+uaKRhzNBbEfOQVPxE33LkJwL23teJa03tx8WbZYTOPAP3Bn+Nu
VFVzp2VcycjWfHNE/61N/pIbhbGhi/Kb29BKOWSJQhE7p8iLhXk1UgEk+NzOgeom
ZtjA01h3V61/dQkzNXikv6CNW0j3wcjLaU36XhXFP3b1uD8z3DxfNJm71ND9f7fl
0c243hyZcy8B5V2AXJm8cTa+lWI+G426Syj7dK9s46yjbFgEEAubeM4TUmn9xE6I
iX4znsJ83TGAhJylkA5EC+tmCQtCQpAOgPutSFCF5WQ6kAn+aQW7VIs9AvO8I/tW
mmFZq9qZW8DK/2bjA4uHt6wZJxc3UBppN5E8wTHN4WrKAkIBNIlhwssMDzY/QY0R
w1erfIb3sX3C9t01FjrEZofSK8PizcRATC/GveyGzN4tSecsnFZqBTmNeUBj4Jr3
3cPNHoNSsGKfnjjlenncPADCCUfwyFFvZYnUNnTP/CrvLzOk6Ssjwp3GeGew1SEj
BzhgtctdmXlxNqhWJNqDSHeQuekShcVAgwq01Q18w/+f/wApEgopAhe+JAPPLbHc
O7a9j8iJnhBP5FX6SxR/AB19IyjiLExQeiBaj+kcKx3jzuTizgEJ6VM7pcs/HTtI
F99oGosvIurzyBOHUJeVrYpOno0clxWEbfimzY36izN/9KZvd5MjE6oxlqC+sklh
TofHMoWH8Tjq1a71pLBYj2pHtCIByujkYAzaiTM/a+5TI+VT0HudydlnCq9h28N5
Xg9sSRXagX6m8uc4k8+N1sa0aC+p/n+xV46xc7Hfv+t5IqT0atRRz3GR81QlHpbg
e915NtnK4o27ruh5H/vRGtmtRTnHYnZVm/dJvcPfBg3XNfkiLRCJuD5W8tPm5ASf
QBGg+9vcQp0F7KAH84QFiwgwTS47YNwiiZgthSo2Q6L6nXPe3YY8fnqyvjhAVmhr
ZT46wA+eIeJFUtKvueqX6/WiDo3rblFFArna7xik7l87XJC1Lycb7zvKvoJZ97o4
E4+sjmc9BPmn6dzRh47Gzr+nMvgsr0Z/xMZWg8Cr0G4YPydILVBJDiRbIvenrtqW
BDvwIZrIearmlrqL2UJ8zyuD7ropgRuwl5/CLnH2DQs3kdahwPeuMvn1LrE2Hxqi
9H5njHpX1BZ95owd7X8f0u7Y+yGIeTiu17XjYpWZDCxUzkbLw8wLq4woQE78brWt
5ZhHlbdv/+OCi5EHqIzGEKj0R+F6EOJdvhHWX3/Pi9oJjQuQhGZWP/EKvCIQSuPy
Ud+Q9Ov4INm1VM1wGvgZORxr3Pite5I2tR3lNFBzhrrkizMxzH06QwUn3MjbFY71
LzSaw3IQZsjUr14YMqg/6M1DlOFwaE5GwecV3G7X6IYPKZn3wO3C0IIs9syw6qE0
6Wi4nZz1z3GP6uDuKmTq2283Tc1o7guycRY5qtLCISY3n6EGm3DsMmjaJE6x6KB4
qnCTWxP4HZ+g6Fl7EwYPMo6y3yuBnAsg3F/JpT+HGbi/2V03o4uWxNmbJEGN1Uyq
iEm0L2Sdtir9qXR4Azgm9MOuKR/UQW+0PLHdvZhA0Xtshr5m751zJDaAa+BCoHRE
hCgoFjigmOeOAjaKpqQfsE6XbaNRiL27AFLb02YRedd4+IfCNY0ock8qGwaPj85c
S9ldnzk/uNoQLTN8UCK5bN9Y/mswONu67CmyqMhjBFjjVpYcPEYrU7hA30O7blAf
yozCykTo1mk3pKHeYriMSv5CiqmLGOe8U3gUCUgREiwHm5ZvISkay100yQJt1xJ2
43ei73BQk8DJbqCJ4KXcZdlfqo+hd1vOcCGPv/QO6wqQ7vS+lnoO0g8zOhO0TGuV
rllv1vhDPbh3yPlh+Wb8Dxp8XgVvDWuR7bWGXoFzJwd2GEff2sw0uUcaLHAfNPN4
nZFmx+iCK//8QAF3a0ZQkFDjTPo5H4UW+a16BgKKNiJaydyqo0tTppC8f38jCTG9
Qg7edKy8USuUhlBr2K47LuiDO46CzNdL3eV+86xbCOogCDyyyjNKTb7iLRO13gKK
Ex4iUSwUHYw3xeY4zl0Yh0qG2I4IagktDrsBIs33ZleRydwxrhgEESAXxjc28xrX
S26IfZJLeQfDg6CRzb3rOaMfvcIsmXh5LeTwjEOgPVGyqzXS4ddmcOik+0MGltfZ
DuzW82zRA8FN/aopG6LpiMTTp1MSIjbEmLZVQHsI3A5N4XT2//kWTCfExaA5uxQN
1BVhHSNFSayvx0IEc9tA20USapX6csefjIIcMVfWR3J5JXhR8OqFpGAMlJtj97yb
nqQXSwfx+e/vwOj95axyxohH+a1UySxONLyI7heggqrwxxA+oC/fDVTbjiFhSvxy
GRMwoOd8PaXciy/Sp6lk1OKxOFD00ntMioXrD22r011K52bJ+4BEiaEI/jCvB1Or
LvAQEO6QtmnPsWlvF/0eTXqSIIBXPYqRhaY2dR9Bt+zGGhF561J6rjYogOAo07C1
lMgmSL5KZFkyejVWDqe+FaOA802lt+KPA1+VYjzNlgPOus/UZO8a1oQqaLHqWC4M
qxKI3+DdXnO7FBQf0RaeHsbIOQtX9iTWU4RskRPQ0TSlSCDK5e8ekDLIIcI3e4kq
f7KLyMn9Vm4Wdx3sDlhWolc3dBXkykeEwjOEn4WiZP91pCv8z3XA1TwvveRiCrG+
ELWMf8AKYYmFoXhGXKSONSWJrUTFKeMot5wiu3/qE8JTs2BjJwfISZ33SXHyoqol
TUh2ZGPNoZxMxla3+XtFlJ+qtSbxajtKjE+XCXgSKuus72UmriB02lOi/JpTdFmv
SfIfnP17lruuDGcJjONQfOfIbZeJbJxKQHaxIS97QANFY//yXDmWe7luLkDVM7qT
3OCdrnifTUbW8eiW7NHnbwZuKEs6xp86wA/l/n4x7z2b1/EGNMNcWdF2iq6Sn9QZ
w9rH8+VZLZ7reryDfIrATTwTdQUBNNViASXD4dYMMHR6bf7aIi8E3igKezwar5hx
mzeuxizo0DeY3QIshA1tLzOeGH9E20An10nFlhZH717DrMO6aJsqjfKcWJDlk9Kj
ZSE/ZgTuaC/4YQvbGG/SH1PFhzQv+8fMw0LaOaez7k2VgXccK47xfi/mO/jQImqv
WLETeOQzVgqqnrKWJ8+ahaWLZKXKp8x32BaSAcNB2KCMGC9RCLJ0w90XlnzBllJV
30OFrNqzKxs3oFkO0l5JfvjwkWCS1TOFSMnK0qeQvKhoXBde6BzybcRuyBwwecSy
BdRKQsxPkhQT5By5F/1ZQHTNeirnnHFLc3qfypWHhrnN0svGcvIvY0+KFeDntYS6
WxkF9ru5V30mfLJ7FctFcqPIrnZCsu2I5BfgT7hUyvtUA1kRbgPJJhyYvZP1TobH
bpSCj32+pyJrIrh+MLaew0Mm9hZfZJmPj+z3bp3FivPZ9OTGsGFDirpvizskpYyy
IcU2fjP1t7CpW8fXA820GWidNjcb7CzN6dyaTKqGhUbMnzYYoxEgk8xrfaS8gQDU
aegvuX3cNjnQ/bnJ5w0WvehipA12bJ7IpV+qiA7we6CNSi9vayeu9G9IN40EDsmn
K7hW3uljQRBkyxECJlhIip/Ta6o3FrL6RQgCrIK2MIXDDVXUYaxIhxemD6N2LdUS
vjsDNIzwO7LHFDaCX9bzVRJU1kuKHcsFy2CcmagUcOljQZSxauzS7CbBRO0RmUYc
1wLCUl618LHFAhi0Cq1WPcOUikhuf+7as8WFaePbFzJVz9li5U8gHNJzD5LdtIFG
5UsTOX522JGxOi50UH7ay8+JOlYYoXZzNJkFoVOREdydNZ8AZRLb44d4o7//1vUY
E6m1EEUqtEx/1u/FXyb5RFml5mwW+Ip9eaCsfnDkibhJzpqh/NKoGaX59yVSdWk+
z2E2/X+cdZ4ywZ3bPJxMvy6aAGjACpZMQAlPzRdTp8L6hJt8QwGpbwV14yK5TgEG
9vSsmz3JZ9RN7UD8Xhpigjd3GVAwQxn/LnbBE7LyF+Y9yKGO3+/DiE+9Yxk5bLJ1
DaFizj32lR1eDqS9OvZyotGHrAr8UOCKFfd8lCzCWBlInmSq56N+aSSIGJaNayx9
XLg0WdBb1sTG5Vn1S7Xq4b5+VfmlR+YPvPJc6V7ObkUVvUMp4401/4Nr4phB7q90
Q4SIIW5N4R5gwFiNJW3b5n3FVuhQY9pQLySccgDEs0oTbVMS62D5wke2PUz3pvn4
BhFERoj/0URhgmRScDd3claduDKPdouBU1t31n7l+v/rI/dNEtVUIQbNEnPgEUr0
LG1XcKqjCUIhhEDjCGabtwpgMjbY57X8KFlqpwB3br+7x67LZZqjoprfl80LKSCH
JgxKvY5wrJzvmHoe4byqng7K7FZzeV2cAkHWFhyIxbRJnKGxSqBlpE4x6XKKGkWT
EWtHkCEy/OYpYA4x472fG0HBi9e8iRlu6D2jtf3/9+1st0QXg0Hn7oTDh4Nn0Q+H
PhP+9ZUjo2cBnyIhyvYYylrKpsLGGIN6TuuHJezo7agciuZZpmdSKONspXyyk6Oc
irKuklt5z+2b082N7Q8oTRE70r1OllvI6iELgTmjpVw4EyA4M8fWpM/UCwomjmCP
pInTNYr/ycc4rSde/deLhTNmWboriBJ+fo5pvSRh6wKUXUlChn/7qYKFIGINfqyJ
5Ia8dihjfM9Zmu3SBqz79AhS4NubGrTuK+yaPfbiTwqvlqwaUUmqj6bP8jDsDNSz
aJJfcnwRBjzikqG22JyuUFxnoYFCkw0hhhziz70qU3Jq2lHYmtFLcphksZfDOEPj
NwxiUIU/wAcUtaMgMAN+Gz5cD74qFku4j17p+68TMKReTY8jA73p1ZzE2ybSVQQM
8kzYC+spsPp2dTxVZSbHC3BC+KNAgu4jASPRo565HcAiIDARwdlEJmNWxYWMv//Z
Pwk0IGYHZqu0MfLW7GKojNgbCUBYOjcEQHniJFFJd7lJUqJow81nT8h7amX1GzGU
Cq0M+uFCqmNblpd287Qltgeqo2hgfTTp1G+nCkCnIk1UdAPd7Z32BeF5RwCb5yG0
o/Kd2fBiNb10JKGlNXl6NT7Vg3amprddD+8vLQwwaUZ7pZOrNezEVdlSN6Ic45pa
c1ZWl9MatoKvuLWLqa68GKcjIA4CaJtbh9gowNtxwlwF82/809nyqklBIZLKuFY0
gFZYafCPykJWT8HihAlK3gVlppXp6/K/oo988FG8SQDm/kFBKL7hDv1TZHedasdn
Al+UJBLsPQXWpnmR5OKk/iIjlAi05QDIpnXLk1Xszej2At+eEa5PdtyhtV2LXcg+
w861EnHNBEU8rCHHBvxH4wvIvA2F5JzR+1ks37tn8WH66z9Rm9WO3EAupVILO2vi
0btLTwzBZJGBM8fFXRWUOooLPCxJIm6pg1v9p40wXgFjeHR/qt4I1qCCUi+vKPV4
6zjttCo4XT6YA5gKgDguGplFNwmrdjtJv8zCGqSZSZ2gw2ujgZsdzcR6HL3fid5A
Xk5JXBg3AApMqGbsSYLEcxo77BG2zR3t3hW6KnwFuh4NvLYb4PJd7LyJRJTo1P2Y
eUm02jKCQdooYJJ55Q5a+Ri0l/33aBwTByDat+qVz0U4jWRu1henKZrDOcclWfEM
nh12wjPozJVPn7fwTvif2GHx/Tujh9OFzTuWii16AsbV83qQcY6YpgL1LTxETTbo
Qes9YxEjOrfSqG3KK46nH3ERiU4Ka970wlJERW2BepYON8T3EvjEJgMcI/j9UnDD
w6xkdtX0cI1tTaKxeuamUbCGuVEY60JAkkpIQKcnqXUFixM0HenrEOKzdZDpQI6y
1KdhjsKf3q1Y/CF0LIo8TXPYER2zKnEoVi5AtUmxHUyxTzpryHW2j25Peds48lQw
CLR1nf6xAXZrUtPDieu7jgmjnSMqZK8KnalpHtrMKKAf0Il7vedy26toBdrxhVz6
ICMgOaybmGBNued+z3US+xWU/jl3ydVhZ5G+DOVefUgu70d7pkHiU5T2H/tyfJE1
5ykayp4QDDcNbWi0s5Up3k3fsi5/N+hqe51Ud+XVdSZ5jG7AocqTTdjnzE+x6DlK
W3+SSLJIwV9k7xokggi90vAL1Q1bJJ75SPPlPxQjN9m+pAN+b1UkQ2594p9aKWmu
xGcS9RHfdDrw+SVhOIPaHZxUm1tqV4djD2Y+Yj148DLoyaT9Qgj0XkM2yU6mCE5Q
NF071NNyLBxf8WQF4bqw3Ymqd2TMs7YpvL5Rt7Q9guK2NfLx46akTe3jfV7lceNk
05ga7FBvBf1/Akr9CD5U858kMpySgFRV+jSBCf1K01vbmPUieF99G2fiWChSlJ77
oyi6Bn02Z38qx+6sBVR6QPsPR0uoyNnhtZ/19VvKa8ihd7Z8v0KMBXHJTM8j4n8H
m/OQQaLAdgXicvPHs+44KebJkkOVY3x5p4oibusQZuyk8SPl7DlbWdU7nB5GJZRL
qZRxIK5j31YxRqAK2ifY9SHbqtuZhldX9FMB3/RkeQPzxY+v1D+/o27yVXyCM71r
UXSfKmmuil4+1COZCM2J+/n2XZV1f48MFolez2cYBW+Cnqqxtl4WFrrMwDgOsGCs
1gqTujJBIn2eECoItqBI7+S8wtaZxFeYDCv4bRTEVymjsLNS6cnaYWVdLBZid1Kl
Be749+xOHBvLIpuolgmjUxUc9lrYz5Jwa/qi2G7qyjb7gP2n5Vme9rHKAxBnLDVr
EYP2JZc7mjp8FDl5XuGCgHWG3fC8hZM9nFFCycUaKAaRWqZP9bxweNCakfWaXc1Z
5qB/jbjrrpHPlkNkkOB/H88MnBgdLuxEAmDNqx1sPb2cpJmIdQUakhWfIt0Ti2I5
DrhJgW1HAC0tLvHLlUUomDCwzD3GFQnPilLMflmyuBQFUl/MIYrr9idSoEXGgLnT
eWUOXp/vnrA9D78fpYZ0VrEcW8RJoViY7cr8jNz5hYxxYcfLeDo+lgju3+bpnLBf
VKtNSKUG5lmq2HejjDDapmsG1ytiFruMqpypzb1d9WlyNKtWB+RzwxZr9Sr47tU/
Nb6ug5UqSq7JoNMXRkKIbNFrA7B4+Qqpcpq5Y6O1nl7lPjZq5loP81YzswfdtEVX
XO1uSd7/CioQlNbSYBGIEYHWvxdNgWje+TVcIh1WPY1ILQVJ2bSdesfZPWw201tS
PceGhQy3cb4DlxH+RiHuV1c9TU6bb0CQYgWAxBm/H+RkZx/7HUv0/yesmsxRucKC
8grUpG2WY5/JxhByNrRSZM/OppGyULEayScomi+SVVIMuspddy+vgZv9B7bOsYYf
F3ORamAlREWDCNsAV3w2Iuw1w0EWGnpwC+etrXvRmb9FFzixCCU7WW3FtM2qm3m2
SdM88Yh8uacgssEIFv/p6/zsCbwooqq6GGXskVDhzcvSVRPoUjUZ/Vx+rtzVitmB
Kb2Jzf7CnWRoANsfbUWjcpr5F99Xn1XAjkeIXpSx1slOI+45e67XpG/P7bPL/bgi
wahkWser7VV0JD+VqBogHFdrzHEnSEgYr601gwgRaJseCJmOL35qGTzMEulPlzS/
WiB/rlGxaucGqDm1wN4iNs7+khNHaO6MSuLowEr6ssYsF456wdjYPO7v/NtVhST0
7ozIB8K7G6VPWzuNinyCspwc77w111tmudG0XDNepUNhhxEALPhigZXo+uBGI+rn
/0ivcjpN8g8E0jbrMswzvUdp9QKqp7O+ClFAEv/Cxu39yRzn/llIwbaEUHrUCONK
p2ZYRZMTWrD04kb08SNQRgz6OSAuCGEZRrauYjh6NX8QwnYwxezfycXrwFaADy6B
xRvVzDTA8/oxwIjk6GqGVFBcJAnN0AM2GEWS5mcIJyl4C/LPsBYQzOu+L7DZeErS
2nT6lv3BKEz6JeezEqqK4BkMJx9K5wT3f+urpngS6RHjug2NAJAXCpwS3hqF1y5U
i3q2nJRrO3R4L1CLj7f+eJV0xORBfFCstNdPl5W7jWInhjTa77Sr3C0bc1vv+ZMR
mjif1mEoU2ZtL0+ZsbTu5+YeyYUlHZANs6qxXpmVSKJFXswqztxnDSmVKuTmc+BV
LjfArjE3UhTBXjBgw48RkZGvZOQhJODqr7qUfDXFve9CiMGRqyJO5pgHuSlzs/u8
JqRCyYlVqbyGzPSEJdMPBxwbLxcoN7Jm/xMxnJrK+Kc43PIl6VleUbTviS2U18lt
POjQiJ9NutXd7s4N04w9JAsJx/PJTyjoUnwk5Du/fsrEBXgd5UBzdpcA2P5AxQC9
5N6YSLPqj8XIFBrYcC6eIGeaJaVnB5BSVmLlkNfWbv2LK/W2IMz7Qzk2HRqUL2UG
WjLv8EcOS9iW2OU9BIf2yJaV8DtQJc3mlC4y8bHyg7Li0rx3IeQWE/bZ8kADtgTX
7P01fohI9P4o6+W5CF2bsdB0YUkM6PUQ82ysc8TzBCbLJIpQ/tO+1Dr34h1DTH8z
YMGCVnTDmoF4miyYkZ+kyZfNqXO+cpAd1YUreiTHnjpToew6qmPKu/ILjpfBm2GU
bK7hpvwWQdZCNb0j4dCazddBjf9ui1h1jdmkhxLNplK2bjOJfVaE2cX5gdfjiZYr
n/OZiGKEoCOq0tWJFc0NtaUJX29f9UmDQs3g0USvcrnipsDEQ5iuA/WS7xbhXaZU
gcl/CJUCi6UDq7tNahlzIIphWqDCAa8Yn9kT1S7GJ89jdRLrwhuTRSDhGO5FbpO7
t8oerlyjAhBXobo13wxw3/D1hO8HREJevNH2nfjxASW7AbtjT4Sk/sdISjtboJ2D
bHJeKoSE0sD192XYTo8VAio/eelSAAW3ga73R0Ou2Xn4BnxGqTJ622+genSbR9zs
BONtydhjsIPI782nXnu8fmmkgACXUszSP/HPPqTWXyj34Zhm65DpMIrN8WnVN9hZ
mSDpNUV0i5YTYPq0Y6AlmADH3OtLuCKUr3uW24GTbJYMOCLsdAL9kJx41Sk3Dq/A
phFtoFx/lBaYzXQf9BK43z+dc6nWcXztMAK/L/lJDkdU4EKDILPnmch7sp+2A3l0
buE2DyrN6wUHXOEPqanyfv6CFaDY8M9x65JP6k+GcKIHzUCTIfqV5co479QtrLZR
wVs34v1x9yXZ00WxDq3+msY4pI8mcvZcDMyzmMTP/5mKwrzQc4+c43ViwTtWTSFV
A78ZGWDD5bOMM2jkMfYwGnSGnYHZaK25MRP4Gnh9WpzStyr3cBMjQowaWroCXHuS
8TLVn86uYEbyRkzU/apvTZDNOK2DlaYnx5gSh3gmLyQ/pJh4mfq/ntGFnclD56Hd
a3D3HEwBghtTSJagqKFvOrF0SyS7r4TK5eaHqItWA3pFWZnDTpw/FoRaf22InTrx
ZECjI204OggngLMAS/iqx8hOYD3kh3tLS6CPcq/Ui0kzQCQaD4EKtCzZYRYeny0r
qWCCcxC2l7QaYvAZJPzBC9TtmvjbrNaXJIgsQG4ZsBAqUTZUUGAxHUBRABicDX6l
9Rgw+WqbGLqczBx6qwmjCAm+evZrGbwBJQFQ9ncsDfkv7iEyj7kFRJYHXqUA/QiC
u13XX1nTFjvL5eKTQYDIx8vuQaVgA6/xeK+37jpjL+zs/MKyBAOeIyP36BFd23el
QNokOMhOHGMcLaJh5OPb6dNOzEGKXqxUklxywk7cyKOspHC2tHry7Nxa+nQtgJR7
icnlIC8D2NHKdtb53GqJkncrBwYMRtUrim3E0Gbx4d/rAEsfIekunjLC9gStPyQ7
OmKbMgky6SafHpoRo34wyIlSYwQpRjIlmjXbhi2h0lsjpmvT2FFzkrga92hTGOCc
CdtvoxG53J+pW3K7BAaeXH0Ezm2hB62MnAxA25oUlxND2c8/NjS0JkaL8ZRLCP+F
opuo9VPnJ3M1nxB3W1UrRPx7yLYP/MnBpnyKkssSwnRhEH4+g1yNLPcVYUkkmuBv
qUZ9RiaMZM4yWQ2e8B6/oCHA7u2CPqD+VuGkAqAFupJsJTZUk1QyRi0TWaHbfSqD
Us1Wuc0ZNvnEGGRjrLuEGD79zBr6zQm0b3fM+GKIP3T8daOZuju8+ID4YsoHj/JW
YLnvw91yIXjwFOwjiXiQ5PPtZ4GTa/za5qzVfLs9/tR3sR+j1b+KPHC3P6Kino9y
xdl4KbSmod6EP/7uE0KZQDg3jkPef6J75tlaikn9QqXAcXimUBuFAmBR0FQkRmR/
wjvLXJEEdo/lToMCNiygl9KGjo51c19tuQ2Ek4i428hFxPNJrl0tHJGreHF9rTbK
t4NHY0ymTMRzLdYC4vRSnjlXLK+qoTdeGpKVdGQQn6KJjFTs7b1KSq6F2Oh+U3dl
7EdBUN9hTVOzMYOlv6sWx+SNYR6Qus16WJK5kqboMbI9V747Y6r1ZJ8hXSzOoFjo
pEVL558Y+dvxpMHnwVhBS8kL/6Qqe43zZuKPWdBkOgYA37I/yx7o3NBoYaO7JY36
vTChWvidT7RyuYyZv/LIJtMn+LlP4S9ulDIu03WQVJUFJ9aSPJmExS9yIy1dj0ZF
MDeWd/De8daiHiZn5LP/4YF0/Ah5xB1Pe7Oh+zcgV+8vxE5um6LNthAhgvuBHqai
zn6qB+8d4+qk3CdtFmeJznANrCBl94pZBI0fWMW0OHPOOdr8hDl4CfsmbsszVHXB
uw4MpaMi1KnFoBRjGRyL1dNIbaI9zWpZMpL6aHmHdsRGgjYXaZ2QVLHbCPOL9x6k
AvQUQ38tfcTlmW/WFyZ/wPlWujSpgYcMCkPsdbzd9/9NnnGbvNMzAcMvdnO+BvPD
HfjmYTsGeVnWZ4RKLF7kTS01WB8ioVZmcIQFxsvZzPBg8noGysId81mdtzdilyod
XN3HAIqflQ/5abIEgb4LTBI6Aq2sor3aDIlKN2Rs4di02LxQZpaXPdaLeB7m8yMF
qg2uAXqtUcEAlyNtu/bBI3Yzr84kUI+s4PxUZgTGoiaFFKlfbBEcO+v1VANKwdJ9
hWVjVcFyRxsfzRdSbCIvnb03q/N4TJ+ryQqOttfhANC1IczZQqGghhD50OyDURVe
wJFKqldnKa514lrO4kjqWzPK5FuSHUL2KmDKPXz/tQkehmFfXqG04YG87nfjyf5n
U6nWVJzKcRhEFhCQY7+2ilrPLZRlkFhNzTEfUscn76GUOh37zspvkNdbnsLH4M/x
4PvTCaV2a/6uxe37eedBQFSa3ELADv2Ln5a/WTEbPAkYpx1CI5WnspNp6EPYdzet
jShzGfAPNccGww1fviWuiuLsMBRA3AN89knK+ymRADMZR3s0Vqs5nJLudP1ZbPjG
8ruDC48sjHK1YtHKeT3yXVCGAAVN8oZqP5rWg5fYQsZ/m40EKnbvEBCnzz2IlLyy
sm7xd/H8ckj5WOH8dixJT0DZFRGVmEb/we+mciWBolteTbUTfJub9tvgHXxU9Si5
UUjty4gxDKAG4cl/RwCCtzd0h0eEr/y1eUHPkL0UiunbkiKQYFwq7W5Qqj0Wbh9K
CPOwWb7C+sTmkmhFYMfLRnd0w/kf9pUOQvtQTDUbqlI1HJbJPmz9j4MGDvTlgcrd
KeWVC38/EN1WvHROFCD2encdmEfJtXLqCKOITsuGFDVEFgiJgbu31z0W3Ue9ZbAb
X5blEK06KJ4VFhEYlgjlmaqlzgZju1deaCjRQM5ZxX0jLWmNzH/pKcpDjT/ZurqB
6M0/rdAFPe7erdfgR6fJC2TrElWTywA60TazvLBoTPJYHwLVoUgP5EnHQo/TdZ7t
fCq/kM9In2ShZ/wXn0h6Xrb7zGkxX9LqmrGIeiwS+IF7kobWoqba294z6eNpcC5t
UWWSpJZftEN15JgTdsugqcG8NwQgT3FetNrKvC7aLhNya9DbHO+lcD+d1+cYRcIB
wfEMIO3L9KGQh8nTATe2J9mNuFzJKqwa11c2RBG+Fool9eK0nFM5+dR6mO+9LZF8
0BZQjSVvDi/oVTWa1pmgfhI9ON30eI7ivQVEXd/6nzNexXaTHCpCWOnXW+lZCRxl
8fq+oKYDyr50v/CGFBtXCBTw1xnhhVxK74PwSo4bWlaLGaNKUzAmGhBb5lCExbXl
q52WC1Wtla1ml+xDDs7FHRC41AeJflkRKutbHM0+Ye1n7QnsnZZGKUuUAzfGJcDp
4YjVOVGDtzzgDW6WY9ozCl3bS3hTqU7ySi/5ZjgRHbvK7Bjfhieu3j1rwGAZjC6D
ui2E5dao6p3V5TTpb2nxRogdeZIkZIt9DKttU/2qDKw3jGG1UrscmRAI8AO3tq4W
YlS8yJy61cBFgSV5FurpOxZSw191TrH6y/6CLdAeoVpeiz9WyoVXMzOVD6ZTYkad
a7p7uz1VH3y7xi+T2Pg1yugWu0y0a31ZHYUcwgTrbXnOS88dUBAYrzqTdS6550wp
WWxHiUWIYoCIsToK6lJ5gi5kI4i1JxiT6poOdfIpOW7VEijY3qpNe0F4jrRWlCvf
7dLSKLUcHkyuYcF6Ilv6kzomiUnBM/7e1v/1+7p0nj1yInlNxHJTZb36WDc/urNh
atowNgogfJWiYhkgZEyvJ/milK7ra2kT+jHSTky+c7cooodGkWpanjMIeT/HYw5s
p2pURrbF82B8y8Q53YxpO4aSbddOHiUYp9J4YlTEynF1Y2ZnDLhrzpSX33EHNhZP
CgWZ+3PjF3Ag/dVwJkmkBRlF4J/va7mYFU0a0ZoHbcSrIYF1WgCetq7og1/SeXf7
BfWrx+i8491RryXWcvaQpqB8NwrZd6IqZ4LKLn4n7LOlBosd4U+jfvjlkR2ns+FA
zsZvzelPxurdPCBioo2M9YHiHgZXzsnDOBNVDzg81xvrUcLIzAb+JmMzSElaQFjj
8wHQ+apJpyTNCG/VVBOs2LZhlmbfWj6kuF3y+QXsb2rii3qp7L/m48qnCLcqOorx
EfIf5A4frO4AgNdCYq667AZhqc/wyY6KZQ1TiJ3bK1ZfvbLgvOTCn4dKxhlI1jSy
0WDRoXRLsEtjaTh/GBMmXhrsRMkuPVCzuJjLuL0RXyHJvD649Z1vROg7uqNl7E18
XAlYe1A9AUBgTDRJ+8fX7IBr09372jGCA2MSIe4FmXsbVwAGs6saQDwvgWOB1X9N
w4W+hN6lj9JyClAw2VRhqqWAtvyjRUh4uC6Rbis+M7c722KSe2gFRMlMM92bZoXO
aLoMFPPc1u0aCAuwGpyreb2pUZfaK5/1QbaZiAH8pOGAC6qhmbqAX3KNY6GrgRkK
RU064h242Gz85N+TeOFI5syLPk+/gAoaIMZ6lIpepR6zwzgaGcT7zC2/Eep4hrml
MFvaj/06SZgZBmaZAzYDZac9kNKoKd4rklndOKCkz3Z2AOgJPWRX9ByB7C5TZICl
l9kxGph5np8P3AlOXhcuCo+pQynlrST18bkAu5YxfnDBLhH36g1sPnB61lgAaSvb
zR5Enh3+xjbHGQQaHl8iHRMmmt9NPxJrMcDcmMFBWlY8JL7Gtf5hFSZikYAsrVrC
rBXzsMR7W0UiR9p/kGfRmQtUJSRCyXGY4Dmd1U5hD1P7QiYik4h0VEwtFFC1Tg+G
PUk/pqGj5Gs+iQZcwpB4FW2iwJOyuQxyw8PzcD2mWgfb2Znz/+D7me8leazjkVl6
P9PKmQG+wNIvlj1PJOvGc68PTrU09SDppWFp0IPrnwVcVNBykMyF6ubZvXt66Iun
hzAXt386Wkp1cOWZdQrcm4X6et4c4ZKhgLvbWqDD5WK+eqA1Pb8UWXMlC5zd9MNZ
NwPnjI7BGBCa6kJyKHJW9/5U2nkWosyhgnPx3CFlGfe9U0X/dxRzzJu3+OOIZGg0
3qXxPzm0KaxuMv6ycCaG1TgLgx3xQCSk+c78vxVBNM1DbeD5otT5E7M5DilL+iUG
kosLqAFkxK4qx7ioYS3Njh7E0jNzDzjKNseELJxG2NxpG6xhaFilCTXZ7hUkBxyh
aU2hG9aXabtN5SqwjxM+Yc8IijSSB5oHEUaR27TGExt1eP4hVTxoN1ICMQK+MQwj
Bgp+Yd1eU+B3pitpZFCUn/kvVKsw81RabLSTMJeqYaKJpuDSJ9UW1bxyIMOr3FAA
Yy1LX7ifgX0aFlGorW8fKEQ1kaPtpXOIBGHYxq/b6kQdK9P8i+/q0sOcfIwVamvE
LfwySSLlyNM32/B3CdgaUNuhIRTkXru0H+RTHNdYwefS/MPNWkjEKSj2kh6YWFSX
C5iRIZvjsqCJe+m3RMvUDX4dGbVQCSSTjaFVMV0GIk2GEOaJ26DW9fHSQ4PK4iJT
kgMnCdn2lY0C50ogX/VYm2y7jK9dkzF4IJDzZ3OuB3ofx8Ka1IFNjGmF8SJTSL1/
bhoAut3P4UgVIB/xBggpLGqlWjDjCoGnyuskpxDLDsep785uVpnVMmQ1OyrGyBYo
XG53Q9X8RIzdWF6P5fEQEQfIn0ZFeVJkvrbxem/TdA4N8rstsg7kpuyISD4OQf7V
piWz388A8gF9Bwz+mnkVT4fLkFGifh2uGzyU+9HI7sDdt01jDdgYAoswME8OHX0z
pQg0e/NONki3WTVmbK5WPUSTx38bQfnZNShpZ2C5vq1+gwfExMKNqNw455A6jUVW
rh0xkfMJSj1Jm3JUfYCKO3IpA9Cb/CPTvBXIPe2Vd4g0YNWiuiZSrz3pKImFLo97
u5GtF7C385hZnyVB1Uo14+qUtO576uUhNJ2BNfX+k29F3XqajY0Tt38flapagqYk
C4rkICxN7xUKu+EU83knlCJJNwwE5n3KKDsgP7ZHCyxGO9HW4ForYvQer4vfZPCe
PgPkepXC4GOKzDX9hg48HxhqAm6Di5HPaOWNWDiC8rZL1HtYkgjCJSK61VMDLFQQ
uV3PG5tSZRj/AXCfr1waNGOKus5vS9SXkYN/OVBg5t022ZRkJ8TImDLSo+dC1dNj
byOjveizJNcCiO/T2IzPXbRKfadWQA5bv6ANCUdHGSLN+7lFO2JEI46rgcslmxuB
OhLBCjMH2h9483VXUwZHw4Z9vPO19Nexm4gfXLPEjsQrssq6mvBarrnJ1uBdJ+E/
uz8aegSL92n/AvW19xAJzOyUdNqhxPi2qXT5z+T7a7vvyKqbyA5EBH5XnTsJoWbo
6gEQo4z/8eE/RzhX2tKNnXoE6rDrwKl9tliz4hEJUtE4lmCXbfPxbF3HGE/gEibf
aWZ4mv/2EPbS1eyrSypipPcXEUXp69003zXut4XSrawpgK3ZlisScMS+iyktFTGp
t87Wu+Ktl/GWGCvZlZ0Fp5IbfDiu5lefkJPYg6OZmxyEMetRvfxeUrGD+lA2aU4e
XnQvo3cC5PUBD9vVSTqnzVj5eblSC6E5keSnT94POzjJFE9h1oVUVDbC3JVq4q1/
/fuqY2lWSbHkKVg/pUgQ8+P88QLebPzPMYXwOIIiJtS6BC3ZCS2rGzYaUI1BL/Ev
6fdP5ZjWRqThqzuPW7q1lXRHCX423u2ekS+tpFCwB0OtZMLpOKt61M6FtenhQ81k
9MxPIq57qPcqBBb/IMFz75dyK6CLa3b3RiTfgHt5CUVdLYik1cLO5UYpnGocel1U
g37d/cO6o2b5ksNCYp3EG9BfEiDZx3SHCYbw4WiujZyZtZUXbRfH/9zcZERdC2VC
JMsBVC7lP3pXfOLwqNzhcuKo91K2tCLHN1A9sFz7RwDzG2nq5TrxmQhiCEJ6OMjd
47VFUnvKD86cRKoL4evUSPS3j6X/nO2wzFIV/WySTg9+UEoB91jQ6qlPPHDURrUk
ER26PZN2IRRsJC1DyIfc3tsoRjN5IM3By8kwCdYuVLL8YlBnSdA+SOy8YsPV54ka
OsGPqepWSC7ydyZRAkv4v+l5niBlPGw/ia4NB6xTpiMhmzmRRKwFjWvYERbpK62I
6+ambxIO8Xyq4hUi7xhE6c65rxQpCQrqt/prYU9fuadTyEw+L3YsrLl4Fo7XiT0s
iW4H4W9noU+dD5Fq8bwhY1b7gTnQXcZrj43DSKAgI+MR2ZkS7bUYY9vV6hwqFDpq
QLLIEbTwEVmfHYQV7W8RjP66aKKeijKXYRty+JDmXrVG0dZIm0heWqQ3Rtm2xPgY
3F21qyxk+QD5Af6c5svaQyoadudXMLRDfpVlspYbJ5W7YTF1Y1ro4shRjOJf7tet
Tx9pNytIRbjjGV0HXh+OO+IhksFRZdigXvqfXmnaQ25N39irsb+PlDA/XJY88s/8
CdgDxowK/VJZFLmvXkzOtQvbdiuC8ysYKRi1SX3lsZNZjYQBixi+1cxRyJiAJimd
cJKVYfR/spejfXWA9c/8lnE5Ia6Aen3BXmteTJTGb4lCkOUWplfMs3K4eYuxQVBI
pRyIfzwVEHP2E2Oh/A2Gfe6MBtJxdmySOTyr2ZFUck65DcnEtpBvR2qmxnCUBRWm
hts2ROik3yKvurRzDNTOTvStmD3DBu9z/5HVuLIlYrXezGPdP+gJnZ8vLRpIIofy
x1kLp1Gkm5Jg5ex3JYI5znBWMQehSfEcO/WuWA17bWty8Z5ZGl4bvrmDlbCEARiz
aaYUGtYy1jZVGxppLftnl5lVTC5uOtOo5L8fY1t+qn14e5GwWiCpQakmPTby0veG
Z0dHToC9w6hkFvLLTZ+4DDd/1Bco0X+06xdpgTWTIW98cGszC6Vu/TA3ntooYA0t
mVKCK+m4WX/M3GgRDGaAT62ksl7Md5AssKklj24ZYPNAOzCoa+2HdIrJTuy7fXOK
b1sPB7cn3bI+VzISSwmAm0eSW0c3FCe8uXJjho0BMfMC+gSjViLBXRwrX5Jjj0TS
KihiYpfYRSvg5jQUA7kH8WwLKZwaovL0rrpC18DN8M0lf/XCaMeD1RQmmU4f4oJH
7eKKDsvL0/gx3XN9qT52pysZAUkTjNGtZYVlVU5qcpRKp1XbUXH+uJtfboUoh+CY
9lrEzveMqLjzTzxPDtcx49jNF5LgVminKVsz05jrw9R0SvfBRKmFK6V6z9xMdeGI
uh+/pQSpLbp3ZKDsvcpxL37ozftz22PkeOVpXxPjErmoBQ7+i8xTQ9k1hTsYO9RL
3J5/pvcgisk5V74hYuyKCioM1LbWNXgqNla/Gojz3ZGUM8WLUqxAlSD4J1zuzLpw
DuRCrM6nW4uO8h3u++3cGnKhhHgVoHJGxo5A79K2Gjc2MHkTUmxrEZf6MNduXioY
8u0degSXd9Ozm7FTxaL0NRaUo5prgy3va5QOOp0EEghZERNG60txNOSmNpB25TdJ
1CvLh68pL0I2ZNa+h6lqR6GpFCHl0+c8yErmpok4y+J5Y+sD0HUDiEsPxNA8Qe96
8+kgXp418nCiC9sRVVcegWvPJWkhOuVRAu3KUIaDhAQ6gGyToCCKfH+hG5KFpq5Y
DEGPGNdFxieraG7Um/NvE0giIAwLVem9JsuZx3uqnbOK+70loT2RnlWone8519OY
Jz8nSKuXwsBRaKUjC7/lZaTNFFLG2fXUghfAQRrXBjYoOiD9RLiWUrfz7Jq13VY/
k6eFy10Lhwy29GNwTuKFYKF8phCMmRS3Kew5pV+f3i64J7KVwva9i/XPVT5jdlwh
MaL6DTKed6slS1ehrQAJS3YSEFwIMu4MAeBlLs8R+1ANE9CWsxSFoakpTS9lMCuo
VEBWZQZzn0xx8d2OYsW/Hi9B5nIgltrPTBgSQ6/KaCiuqZgBS4n2YVFqyuXzhgCE
tDm4r0n7fJc9zEcwcWYBQWrg4FblvVIR94WZ5+cNfDhnPKRHkYy5NFGbrEDkTerM
2mzpUXoksJ05/1cJMI8gADgbcQQIRHViB7N02Y5oufN1az7Jio5SgzMPvKTQ9teD
Vh9Vhc2WcPP47fEzp8x2xcR0CsF99Q0smSrQIp6+EBS4K1dCcrmnJlH6hhqUa8AG
0gNAzviKr97ezCNe5KNF0hBN/9DZlGgwE7zDX/WvuolK3fx+TN65Gw/oVl6eNS95
JnIOJHS25OFj/iTQvORUhHJws9lDGCNYYVTbGLAmZWwqO8wFRJZR5nZPfmMEcuVh
fkhvrjJCbDRemrjb1yJnVnV5ZEHsqXKR/IN9lW843GEiOELyLwA3CwEqSyfMJOBP
qDyEC9eJI7ad90vm0MZS3xCA1OOG8HgTTw29/j69zMSeM7xt25WYu348yrOcU/AC
N9MONSuIKsqAZJjK4bCx4hvxQe78dIzOwALNkxS1xM8EkJrJJRP4oY3f0tnE4anO
yYse2sK+ytJCMOKaXgJfV0uNlvILRgUhUK3lV8FwLPqF6XqRyt6ZlnAzr3Nsuu5r
GAx5m0TU/DUJHlijwdANCNImw00dnSabonb5fOXes7NDwOOFkd+2qR7DvlN1RFhN
7C/ENneP8EbkEWOPhIxiqVB6rMmTk5T7yh3hnGKQaLLFOKzo4TTAmp5uBLCbFJju
2uFcckz8TC2gWKz6BsB5AZervLy+i/TZTlRWcbbOoUmJGfF+nGTDLpZAjMiZ+7+Q
OFXcb37Sxw3Ra1BnQaApLjyW/NFi4yXkkuIW0XBdLoj8wYTgD61eL2jQ3z/mnDLa
MdpqrfT62gSKZ97ORT5Yox4+7qB6IzeTDnXPc9FbXhXzKn03u3mI35R78Wsqaw1o
wz0VUyzcy7OGkM7YsnbpNirl8JX+Ct3tEleTabesz5AY8uNTwZ6x1vtoJ9or008b
X+ePRIaQbYmdykjhQAAfhwwYC4s2QVI8DZDwvcmJmcOHj1vJZaZgQZfNuNy2F4Iu
qDjaNbkWFZY9ziVBACu+d3Aby5EA6C01MG1cLrZcam2GTAF1LbEUI5mRV6ELrxBx
90N/GlGuSmEhSKgqHHwx8dgRHVQRpgv1w1ePyYLtU5jYKNxcs/OIMqEhaHnr9w2Y
da/xdyYRPA+uPRwUdsiGMmqluEd9DCrnf+bQ97qD7bLdW4qd+X8ccbcOKsCDZ/l8
mszEbjGXUN5EbdTmkuNHuBPh/Az5sF5veGRIDyolhtIeEaW2rHmF5dvXcc6zqCQk
UcS0N/MFOXS+a4DYWezUtXqQZ9RNr+Su/OtmJITvIHqVZJDOvGCA69pkvJED8vQo
9LNN2yTiJ7TBWtSDc9q3jAu7uuuf60odYlkv6HFQ8H8PdvHun6LIzWqSZgsvpuZR
UtpE3O7fXNlJSa67hxMp/XFrgG7uOfpOKEgCOzMdhpdWnpEkAZ41e9vUbpV9TDin
u+aqJUuzpgKzrC57FVcrxlAB/vDyyLLg+drAW2mzkV/5AP03Q8zqBBQ3Dtfcjf7d
0o5bBS4FHdyOdiPeb+gdnTyNjRXcIGuh8sDl36BXS2JqCmpkcy9XG64ko38sFv/b
TpDbpcJ0N9OUDhScaDsTrMKL3QPSMzW2487AWEt2OsbW7NsPpV4O5U2SgDAVIO3r
O6Km6bdftrkKn9/CWxQiEtA53WR6SEQRYAwij8mmhOra4iyFxy2mayb7oZaRPMTM
c6Oorc9/zvLD+tUjx1JddNCp17zQsiVGw6lji/T0wIzg57ZnctPAmtopdPws30Le
U8GX3ViGIt0MuEUUWq6LSj9l0IF7Ci4UOuRb/O928bcCH5QHMXAuzWoLU8RE+inD
fuXOvARI+HMP5YGb+GJtHsFCJFEzB9h2bhRS9VVdXmVr5ig52aEZwzB+rQjH1dpj
mkiFLvYGh20SsMw21YcDtyVfv9oKJdehVZOnc+XiLLfQMsooSAWIYb9NMCkxFRBQ
yX6Y4fmZfRZcLz5hUTsPWxoexYEQSuc3LU5bIrkz1ZW+ihZqSWhPPigVwmrpfT4T
uvvKGahi/5SW/mNl4lKuJIJPoS0xCD4kQm1pPiSO23cEDOWWByrBGfvYLhVOCyYI
I7qffM6w51SiKc3Vkvtfe+9GgyqtkrXmHy5pYFezW05sCVLB2C8aPi6OoM6Sq3Vh
AC/VgmADgv0CTeCzBkZrReRndGB9ZtGbnWur0BkBhQV5iH5tEpiafFwRvHju8uZd
dSoZeH8MBsG8/kMmoffrSf2cyXOyQKUpWrjNznrshMMIKexl5VXXE6AMheFIyN6d
6+Pq8wze7QVPgPJP9wpxspifyPeEgdHO/SIaiod59jqxzbEoeNQPEb+IPhj/I0/m
KbZ2GtCfRAvBCkSzqi3VpgiD27COZCYwsMPxzYinRQT617fuq0kNkvhKIW6unz4q
fzmV8sgQLOBkA3Swl20n1VzoAlpm51K3jjUAMcg+c2I/a4/Wq4kRM6EVP33Z3xh9
oMn3qR891ciUcajPCLTdc8m6nH+az3hEAKmQTL5Awws/uehdm28h0jSb0mmFxtxR
bSdKfdSeTwnikz9642d+TgP42PMfkQKmt83r/euLZndBhwHWM65wQo3bZupxVmFT
+FoTVTC4cl9RvdkJstDM/Pa1HkLdCwOwWTFAdHMtISJPFu+7K+8T8l0f3+jlho9w
CRI06EZ+XKkS2JrZrKHVBn/z8DMeEi6A99Y0ecua+s+yvY2q0drVCyY+O033Fofb
z7VvYJRV7bJoHLr8FXoT+6dB7JKclRswpPUls/xkzxYm0F1TRNVvnuVxTT+pBSaI
RjWcZ/Q85NH+miCGCwhGrgqaLYVbVXYdjp270GrF0GbPDwaMQsnRfZU1s8X8Jfbo
hZaOFVINftX/O9y+5TiL/8efoEzQ9VVFQAaBXKrsNskCUjSEmE75FvEkS+8+07Fk
hRIadnntURnOIsXsZtpr8sJQlzEmCwDoAKttsoieDahECdDhZr/tJWJlH1S1tups
MZUqVv5jYF+pRieL0DhQNEypKDPm2I0Hb/YX7Rao5q+y2cIgLug16F6dhkMBEmXj
9zWqObFexC8Ok1BOwqYAkAGi9NzIOQ2ZsaYNwpbmNrBCtXUb2+J9VK+8uBtRuimB
7aF1kPE+vJ4dncIUn4r15KGw4Bt4cbGCRJHnZpASvlSF7KaSSCrFDmj/lIRF5rJl
fHbqp2BGgnnVVE3q+3o3lxBtJEPbRoi9vqD+gpXYds54+w///VbN/xw+6m7CIHzt
IyUCJNAbZzAwCTJntFZxWbV2fjsTjQBrc7YUofdUMlVPa3miYMxVZgUKaXoazPo3
mHWCamRBjSEcCJW4qnBKVWGGoTi0h2Z+6GQdJ78f/c0EjbgJhYC2Pb/nQS5do8Mu
FrHtcFkyT3zaveArZKsjL2GAngsmTW2bG1joSwHG6R4fgq/USh1l5u9+WmI6V0Lo
oUd1vu+YqjzAZPfqPAWbtNKGvnrnc0AOdjcCrFuYcO/Ut2cE841sbkB6dZwjiL5S
vTfNoLTXdkY+faBQnlm12NqvO+wFr+ENSzNNn+rvSI5rUNSdCvDDZoqIixWrDInZ
RjNmpyn7cSk7LGEc955LIKeYPb3mb2BQFA/WDs+YXpbDdw/ZtMVUz/ezPS+zciSa
3jx9LeUKrGeb2wyrpjm+iFh6AHkTnWMMsGqIKz8bUOk7VsgJjUV/XpzO/Pg7Dr4c
RhqsVsW2uxdiOAnBhrAgbc2Lphc+XP1KxaBZw+pWZNRU6I023Vqsw6hTeg9g9VEs
zRaAyHZ5xk2aR4asx5N42pRbttC16LOG5bK88OTdNKTroDStV8w9BISZmT5nQb8D
Y2gjDOy78ZpCA52PZj31tw60y7Vd+RL7YDL8kNj3EtQ8JQ48+9Ha8EMM4Nw211S+
r21AV+KH+LrzgAL1CQtR6QOetYvD9SvQzXqg0KhRsR6h6qCFLsZ5SsUGMG4M73M3
rD4G6rsXYnThV9iizzbySnzj2BP4uKDKeW1WvN9wXZER73ww8s/XZMuH3kOOyc5o
WZCuFTazfXVT3DGeZ3a7A+7MqX/883X/g3ef6eWsTtCZIvAGYsn9tSjZB0qdeWZ1
o5Jaz2YS5DvSUzvcG7ghCKdOnc2DO3xBG2F7chxPKE334BsXnyH4SkWSTpxRC+2e
YVG2hVcOlGyIFxCbnRnz+ewLgk+gC/gX+ISzgIBo648FrSHlVrbEgCfqE5Lmxnjs
0GbNzfKQXuAAYttEPXCca+jvl7ySyWFkvHUKvQFK1XB69JqKlhUko9O1H+BZRj0E
o275tmsnMdOgk+9taA+ZjUUJS48cDk/04V2A6xJiRBdWVGmnpewfrFkEhW8e0qVx
bRoY+LGgFh7s2dvgQfU6kT4hMMiTr0Tf1HJM7vpqS4sO++xPYkvaklxZRpKAwIkC
mjwo6R/sr5/xROGiNviG1gK+dY89Waz2qOhGZkuIMdY0Yl8N+2wueg7ZAyevmHC7
h5+JLyaRx0a4eC8lzOExq+rRDhHq0tmrbbFwiq6IRpdAPxyi6B4vWzxHe/gZY8vx
SRjCoTMnxse9JOSXwhBo5NkJZqX71Sv74JREZMMuX4tXvGlCyKdchTxbzMZRmhHE
DsJUJCDLljUOFxA7YH9BZZkx8gl/TWvqjGI5Ctp0/s/vV7/p8EbTsG3cYK4pLtu1
whQnOS2wYUnCd4AOWj4wtiv9ZU07a8esofQP3SIGT6zaPN05N+GXe0UH1SHASduw
5pm+yZjI1Nxes8KngThqDzG+kd51QsowQkminOUgGByTM9RyIRD6YJhzVkPgx4BD
t15ciKMiGctbqhfUK/Pua6jPu/NDL2pu4BTS045J49+znHfnbKuctdR6KbbeofZQ
D8/GvNyOYgAW7cdP/KVGSdsXvxnLobyDTEJtsxotCOsjCYJi72QFQRjjh1mDRq6B
1usdnhSM4yqewDClBvuM6TlgZOBaUyjy4K1Mz6uyDYtLQySUclFdrdYKgjcPTE/d
OtmhKu7Pvn7kxailadeeXeDwh9GLOzrrUFD0nIxc8mH3v2o55n9yKKIvuLpdwSDz
y1//VERHYmh5i7GF91rEKTA9cGwBQvjXOeeHxCMwgYpiHy31fxe8qjS7fqIy+dV1
Sj3loNFRRbsoeSNnLO3/Z7IuP3janLcGPT0ld6v/RP1H88N8vpwd/KJiWO094J7o
d7nPPjIQTwEpk9cT3BSSaIZnkFXZor3lRkWIM/2n/KNM7fZwE13exUtjuCdGoSJs
JCFDcgBJXpvv0vw50Y+2gfhIxuYfYM8Q3DUesmEzDpo85bI0dmI+v7i6TBrJ6U9g
rdUA8JS9c+8WZJIC5NT7IhbJ/1xzfsDn+2e/t0XAd7CBoL6jgMh9iWFUUSPm4tsR
Nlh2+fVAw/JR+JCZh8PauNpcq5bGEQIUAnoZLvFUVoB5aVFcG5jo3UsvOW4tqTWU
oclBfyk7TqJ/zDVmVmfGe2XHwf0/qBEidSJMCRXeTjks/n9370f8gfQXJvxk07WB
E56skoYSDh96oS8VLSEyrADsw8/uJMtOiPwWJtqzJzXhiQI6+015BowfXsnji76h
ubOlaBTYb3+Fr4rY5q3L1LxZwIGhqIGqBHwSzi3HDv2t3sHtz/OaiJ8em7pDPY38
X4g+kmC4wAP3g3CTdiEq9bQ0gR4NqiQ+zmYhdeP6SomAINkAtd9eCfbXeBh79VGm
xAS0jUN63MDDwP/diTyQpFGWCfL01thkuM8pfbwfyDyJuNr0aqbzw2IA0xrI4sDQ
6EIOXYNSYkTUmpcjBJJHnUq8DXhBt5S1fYW/evCXvgUa1RVP7QtzhsDJjwAbyPld
my80APHr7gaUobKESNF7CFy765qLTLqrDp6jPVoZXrlYihWktXhLv/e67wQI05hL
5IlJAV22jdTQLc/eXIu9JuYgo8WEunNzweK8t4BgvlPfOu/3YpYtr3XE+zMkHaAQ
8m3TjaIa8W9dlCWa8WSlR3Sn9xiRA0nKZI+fUtX7YGvr23FeLqa6dPiWNew2oH7u
nHPfdUdHJxWZaRiCyLBkF1N/hOsZqHkYwTWPTGiL6M8=
`protect end_protected