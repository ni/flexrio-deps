`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOefPfq6U1Z3z6JZJo3IxjM5vOICIlc22FGjNzIak88gV
OG+Sy3ERAuncDp+oXU41W829IS7Ua3Qee0fK8K2XRVmpcJyW0Tv4gGO94GvcoPwv
/TlFVEhm85ky8c/B3R/8ah9ulYBiZhOuThIRW+7p5W02Q8OfMS70JmE73pV2fzIT
T2PNg4eTldD/7WZuycGbOwp3w/22Ps28rrIS560OqjncVRqlO6JuRdE52ih4zhDX
+ActX8XTaPre30xxD5XrQKDD6EJAgJqbBgtG5KYHGA/HeC/O9JsEGMELuA6Df48B
fqbx9XF+Oq+tZeqdbltqqg9g2uBM8O8xpZeOdlbkSyGX0t9xLqo+5VaLMc9r2ryZ
fdfP6C9eusrZh71UI2iEZ8bQW5aLbv6BZM3+d45kpf62+by5/K3K5A/05TedorLb
lIzOx2BzIuKPpqoEe808mABXLtrfMvHr1IIuvS1gaAeqPiLxcMB+WgWJ1WbLRcEw
gEdIJXqSvXlkMCFgT2sXljUtAh9JF7c5/+oHB3WajkbL2QrARLwBZ9QJ6rUZBKAi
OxRK+A1X66fIFGd4d4w0G62Ix6GIGiBZpTeZ99HQowhYsu+kOIWCYK4KkZeWsMRU
zEUda0mnRyV8wEcu2jZ0sYZODsupJvppoUH/zodsEy6+XjNSj0uMFumiU8EpruZx
rsYW/SxifWLd+s7m+C3gdj/VtJEL0Uuc+kKRPS9BTjeQcVrFTx7A74OBfTaGqVJV
U3jHvFrx0BXslVqSLh9WEPzb1gCtVHpumwId4D3o82G03DZ4VChYiOefHdzslwpF
/1MgJBnwskzzuwbG/cL0C1kS6QCqwszxOkC2mhyklPFEYYeJtwj7FK4w0wBVNZay
P8s5/TlTgUJZWXc/8kJ6eJbhpVKElYaTiLayXeBi+RbvXaP2K+KLxKGDp1SiYy2+
aHt+ik9BCfWa1nAJE4zar6+pkj4pwvyRj18aSNPtTBh0NRzP3uhpjXQUo0KRg/I2
MBDDkmZ3u/ATEPpSrtH0zHZ1RiMsCGJ/G2CcsMvCpTAJsDf6HlnJgVMApk58MGXL
QTTer9Q0DrU6SDE89av6PovSk9G7aIQ7HXGKIG4Qk6eocwvTIyy86EvaaTuncuaT
b2KARGos7A40MbEGPWYiH+ioxbPhy2itKL38CV5Vgbh6b8RlPW7TirUGY6Ss4I+O
nOWa+gP6C3QKggJU2I8vZq1vU1cRfyWPotTf2kZJxoWOpZyz5BZ2RbjPMB5i3rEJ
fc9LmV8a0/J3mRGZCmQtkWWlr8WC3COpmPPnYj2dLBLOq9OPM1YBFUczivOENdUt
aPXmTajxNvWGWaenxRot4A+RlUqC5pJeUSx5W9fi0dsVjUED6Cr6MQwpDtc/aroM
tskd68c9paP8XVNv4gAQpaUr2sz9ODLI/Vk1/E3reRbqomL/hFntQsEDxMcXseqx
f1vD4hFyW+MTLnZwBU6j2NDqpuH3v8OKKwbhFrEYSyqW1xypgH/BCN+t1rt2TZ05
BwWScac0fEBOyWMN9a2q8Pi7v0naiEC8jkuH2PumzfgInWarR/B9kTE8hAs8CBwl
F7HApSsdQgXJ6xqcGv+1PpBbnUASaeDiZLevcDjMg8CWo/JFUHtf67YiG9qhlT1p
TSgJygcvDtlzK/iSMgZW5vnv1x13TWzBwQG64hNKeECwnLjGDgIW3X640UzydqN/
v/fCZupRIzKr91WrP1wJ1OGTPnGS4kf7PFcKfJbuSOUphSbdt6p0SKyu22rNSoxg
T6djQkJqp102XPScuFyTVsSwRGrZzbRfpJjjoeD/ZOtEvH2VCvP1Py43Puc5mCa8
0+GavIUPFWppr/L0eRoQT3bdRvrM5T5PLmlc3ufA3pmsGN92hgZwTOtF3cLfKLmJ
+tnsFdFHRMYxet0hAU1LGdTlRgbOdowDVIzdvimcfm3DWUjIbEhJxwvuHkNR4TXw
MtgtjjPxSPp4fcrvlj3vEdejBj0jC+1FLeXOqcnbIkJO+R35yL25Ob3VgYE089t9
Keaa1N+DUtHyF86sV8F2tTb1Xg8x8vWqkrSWW5sEhZX8ab7NAywX9R7ueVhY34Fu
G8gGaYHIpeKIyPPc1WmJEw1kzPGC8UyIWsSCQTTLOavFnoaGMLUrzJUwnUt7bAYu
oJTUz/FB0cJObA6F0PVtU0/JY0cdQokTZfju54RMlLqYV+hm3yI2LUjIHg9ClMyA
zShtwtvdeTMRojso4MAhtYJnQjrKCkZots1dnWUDoX/TXORWYtMBrltmCB7evHfu
7Hi4IXtdmrB219kPwIj9KDadQJa9TMedEqC5ns1r1cC7gowm0tQxI4E4NY3H27LJ
FBHQ/VwpWCbUxgjnh5Sg7b5dVexxIyc+Gs9UIJ5dvk9rX7tjbNvFjDHAJo4h0IdY
Btmsb6aotkv2WElFXAgzDzP3hzEgoWcrjkJpn5DAB9O9izOLNYOC7JYo2Wb/kxP5
F6rQNG0KmtKNq7z0W6108CnFnbS6d114JYfay4hwAZRKBl5DF5YOstllj7EPTC13
HtZlN7GNmGE+pKZ6KmUbVyKMCwRDYDs5hHOynU1e8Xforkruwhv0G4MSnBfb6isk
0KsQsUX6EAG1g4YnjQngfhhKK1GAD9kvYnF9vQqe/PHJ31MeZq1TQe7hUoLWZuMv
K6tDZwBoOv9j9NcReyA76XsYF1t38hLb8nB/FDg1X5v+AVJT3sSWNqQbp/i1PZcx
xYJRv5Llny2NXbj0Tm35Oxa+3gZqO07z5qPsEuEct9muKk5ZM3wYcXeRFA7ozpdU
U6Q+JMUghV2lADVxZhoTKojm2fcHTLM7sTOTcw/UQDDKJARaQzEoxM8bXwoq2LlE
GsbCHPxyu4ze/XsIHHHTRIVXxXF2nnXydrp0/GZb/Wb1iGQjEKa1Dxd9MsSUqX8J
yGZjvusjUdH8bCI2RYjz9GuwGcFpYwcX415V4t+firPxn1oX/O1VXooZ32nG1lTe
7wmFMg+Koq+a59AB65ucRFLi+c25XWw08UmOJxY44JT88rQeHHny9vFeP6kML/wu
dcKRh2KKVUK94wvExGuFRGHPr55yCXG3dQuDMsyUkR3FDLBO6hSZJDHH7wJkhuMj
CbGus4e8D6s/vIeC1/3qgVXiAxRWJbjtlrqwFcdcULqRvGGtH0oHpf6n8jg0uEpV
Bon1a7S0nUkJtHJYN27ePLtgDRBGaBGqFEKouy19vNd3avCcVmYTWzlS1TE2DTFc
yei4+LVGANG0ssxTqr2H0ZdIUsuSl260UkH1sKetuw52M3lvqadmbJNK/OSgXZzU
cOktG895Xug4nbb4qh/g9gW0OoqQjrL+v2athzY/2eXMZWgMHRyW4EwcAvqfhvjC
rrVzjd4C1EnVobRFvD3Ck/yvuCjceVg6oTu2oIoeA5eDLlYnp/I0qRMt6Dj95k3r
nnIq7WY1weiydhHuByb/9hWzTz0BTN3FbGNHZ/dwvOzCrx3KJjT37bAnwBDRRpoi
ig3rhyRKY7c2QmtsvxZzFywHZs1gKGWvdTy25FSKBUDQmxXCB//1d4swFlQ0h+lT
flMKJ/ak0EXtQfTLuqwm3YhjH7Ifa14oE8AA44W4hlOOmTG0pkt1z8NuZ5egt3Iq
882FSoKY77oSnmFQejMGjbpix0agm6x3jF1+9JH6UD+RMnf4nAcA5Q1h2ooBPXwA
USRY5WDcqRleQ7L9lqCUwL/o8uVJSjCWpqK6rLK6LI4ymUtV8xIeeRc8m66SJcqU
4aPL+YfD5mho4UZOnUX3gDTxki0orS+dhFGo7LEiu7F3hk7dG+kUD5RPxMkU6rHf
rshR7d9pMdtWzgdLclFgt83wLCv7EjuyY7YYlgNtAO/X17GkUfgTI+gFArAeU51c
f7tEmi9pjl74JQp6yUpqFdxGOTkwq5h3fXlBpzizgmzwbwyviyhtdB3FGi+QE3Jd
r2f3+wpyBXDqNtHx0uZLr2M+Q13iTBlQV4fWjmuKDEC+oKdVpz4IYwfu+69HXwH/
gZLKCCM6V4lJdP+pWU3sxCSBGw8Pc6it7Kd3A0S52yrEK9UDOHN89TJeqRiImPyh
gsB3y1yesOxBIXElh8zsNxYEQz3mhkFJIkFlKveJKlcS/A4vLpvLj2/O+rCHgw44
KowD8kQfyd6L2kGhQGnSzmKyN69arhGIq/Z2dk7Omw8uDYOzGZscv0BmQ0C5FKfW
ED++gMY7gx1+wZt4+nfAU4gKoYDHBHS6XY7MXF32u6hm5ovbJS7O5ZhfM6fHzoT9
FteR5r53x83QE0mPkK6RFsEXy0wLvszY3V6QoWjoF/b5DKduk0p0i9731mRVxH8I
lgIXqXuAB5QjKyQDEPVafYePXt5nBluMwT3fWmyr3VM+xMXn/Jb/QKUQeoEJfyVD
dBnTtWL5U3w48nh/z6wpC/FcW8jFslE5RWDxgLhD7vB8iqyb7qsN2b38P+TGUsrC
9mQrVAggP/i3SZ9HMLfwN4biWwOuFsHFY+yUu/boBGxF+FqVCCBghr96F8rAfC8L
2YkrAmvqqHQGzTYdTaajbEq3nIQXCmFTJikD52Hto74i0XPe3XXjN6Z8/WrbH+YM
PzuYz5tH8G8ovuKm9J32N3Apjk7q7UQa4Ws5Z8XTptj8SNOoT7AMpRGvf2ZXURlY
Mv24rghEXPuejYpj+b6xrjFocQgnsiaUyxFj93F5HU35zoYbkl1TtQrDMUyFQ6/w
n/kZJo/faSv0em1K2ZNuV47l29PSunH6WtlmpkbtzYABKGOzPSi0oUfM6CY0w9N+
uFaz6EIoLbm1QevDLLD7QwlB4SC5k9+6XV/JAEx6HjwXd/5ptvWGcCFpcEYvuZh/
psIf/Qm+o9z939AwRm93mmy19x4bIQ8PUqqtkDtkOXbqZDALLKUVe7Z6mLfL7n2Q
t2acyaUh42rcJdnGQSDm/E4qVh5I0d/a9n6eZTCCo7dZ6C2Jdt7D9yporwaNB8x6
rquzM77wtdbCHDvtS69O6jNO9bvW8NqlzjF/RmnyE17sHMQqkwIrX284yxft8voF
HmoaJokvUHtl6A3LH/MBap9fZobgKhp9A6UMSjvNibvsdqPM6Wk2/o3ezmJ2xo7J
Rx+3nTazFGhSUM434iWJc1/482QIzryuG+6TsBPqXOOnWdLBLJmVvvpyrm6GKOj2
CA03T6o2tCA9ieshHW59IWOqVA4XZ7GEP4/jpb+GUhs3SKn8zejpEQr2iswSpMX0
kdoKyl+9B2HqdWUb/w18vMrRwXEPwkKSY316j77qQsUGMP9w0GAh3qMD19gIAOC1
57gMtSSWHyC8WcCu+BHuiuAnq6Ucz765vaZrVZ5vothmQ0rH2xCirZACM0rT8ibF
s4P2l7IAHG99O80Rur21I9byAu3b2FiIrP/x6849B2f2P3r0vktwr3upfku+VlG+
aAKRY2c9yjXkpEHfcC2mBqu8B0Lp4FWfQRxLgoSz0lenymFcGXVZv9qp0A3vnOSa
D7FeanH6r94naIaWf9vAywdA1P9glmKssfHbNzzKHqEYE42esfDLtt9mg8P9FsFt
S+KFfKwT2x7emgMsPv1CdYYdUkwatdA+lVmE96tJWKCiL+oswV6pp1YBpXfhSQcv
fSs4YaEcuZA0hFlByGrktax0INmGQnYuKCm1VHd8yc0pOQyC5eoXfigc3J8RNGxZ
i2HxOLAcN7gmuDuISh/JQn6fML6kI5mSyCIDxnwSM/bX4ytDDnFnIRZ77zsa+LSb
4MQTcgCKkDX6p0rR4iW5MiLHrTyuRxn9d54QPSha3vbSPa3M5oLuUKVl27TS0RNZ
UKPrBHPUBk0k391xsV9/zgnn0a848qlAx9T3DHTs8W6vjwyTXT8szsL1vTKeSlqV
pYI4L6rO506pWa2Wc4Nvvyt/K2TWrfGAxPXPvhM9VR2U2/kPitdfXq0v6OmplzCj
IQ11m6hB3TBIkCD05y/qChaiUrYsyH5ZcwL6I151YHMkX0q/fe2///quja6PxV5w
/9OnYcqecwH3du2fd9/eeIjjrjUkF5blleW784rKyc8xI9uLLAWoIT9RZRg2Txr6
gA3M05yIUvzREkZjLt9lvw/UXzIlPTVeZknAtpFu43QD0IqG9DmRYvVxpoHClIbE
Pzd+D+nS39xwUXvPHiZ42t6HYS1eD9l3gvzpAWe2Pg5/1n2csiVs1G5SH4OEhEfJ
vlGYEDU8cM/oEUkScUAginVCz7URUNSxTqaY1bfeSp/lpi0B5U6iP0R9odzmF119
KnG9C+JItnnjmE0GlAR0nfMMZ5ZHLqXNn57iQG2Tl49ugi7R5WBWdQsScW/fn37Z
2dfFrN1zW3Y/RnJsxmxRmehgEckk+uwDtYN7HqHkImGFcgugbjdyo7n9J5xJDTtv
kkVhJEyBttx92IK38MfQmAaSucK2qwn4CeeB0sx8O4tjIMvMVWxX9X8WWieLVxBH
VDhY45eqU+GunNqzveJe6oPgebECNVLR8VjrtmCFXEcb3tMK1270tHW8XvdBXmvE
gGX0ih/pc64xFJyi996Xrciw/6vnqUXbzPOyu5tzo5CJD471G3PiseRJQK6vCCVm
9GlSApWPyXmjZdhROfaNs6SRtErn8vKMNp2i3fylJvMXnU7Kzuw+4qp7t1TafWe+
2cjYex+q2gPmY18JgfBrMvjS/ZO0R7TJPLgwIKmbJGbY/72qggmWFSzwDLCA+JQD
7lAOCRKVlXtDMFTb/alttA/IC1b3VpAhSpZW27pz01s7oTZSyKTCjex2XadDirNL
4pTQrbW8Pkq7tnpyeiGqQ5tpx9hw8t9xrPUGEMxrhlq6igRnr01jyuWtuw1Ppuxy
CIbF4JR7CSwcSPGzaw+KsDz6BoDi8uYE9DHEAaw6U6LRevSuhbwTDJ5nWpsvjn/W
EWPaGdAywX+bSDxdQUeRRRlj0Z/6iX3zKS2I8B25E2gvhtkB9LAYFTUoMPq0tY3R
qkNu9ZN+te9nU/bJq22waJxK5hifbdZszOPz3fvetTAoAE9qzJKIAKSRRqcb8XQl
Z9k0cNpRgtPdARke7Y/GDgETlCmQ/2lbOgXAlZoicFwJKzUNVRJh85Mifx6bmlid
bW4lV5t2eCl1pZjWaVwsn7KdPurwNg0FZDrjYdROMEPwlXmz4Td1JstboqSZEGph
6tLrPis9zDHj7zmWxNL9q8tnE33Omfc65rtMgR9yuc/tpnRarG8Hrn3fBjC8EWJ8
e4iORd7K3aUyMj+J5KPP+pMnKMswD0yv3nOTOmpQOLCBkt+WSAfHE4y3BMBiCG8P
Ypawf+kPV9UtgxuKKpTvZ7EJabmPqA0jrxqnJY3YmJJ4WdwacrkEvpTR+KQvY7aq
zX7ymjlvRaJRC42qDjjbXmq/q9RJCMgQzviS1XM4+Gyh/18Vi/ROwMoIpBAJbDix
d3lZUofigJScd/hjtAspKqE7BmYCTLbM7Iy/FTSss2SCdat8RPSBErbQ2GguQCyP
TB5oWQvJExgN9Sotwi5thGlfWplyFZYYfyosh2yZkPuzsT3AKodNDVFKSzPrBeKM
aoEndQzHnbzzAtabcJKueLHRPGfmDTxKba7hXK3Bsv0CoQrsJ0DBgM9UDDxuWBkI
IMOQdvDIMUunX3Enw2cHK9fvdosVx8hFsnUsxdhHRUFOL+zV05ISl9AB1Q9BLoSG
Q7Pr+SdBzBLOLhCTD3Bsb7ATGa19P6njV1mdJ2J9ggygKaaajSs/b7m7PzVYmT/X
OpXTkvWk9ICn0fdVlDtc0unxLiWHR0xwMWyEIY7fs36s/f/sNlS9ObPy86xHGu6V
LOevFiO1HZh32CO5RwhiRQsmWddDgiCrLLwFZM0wEuKikHr4jb2fGbqJggBdFlR9
pLlnOuiW9Jtcx3UZ5s0AxqhoNnW7ZadgcknuLRWxm9wm0VZ/EJ6MT9yXh68t0QpX
BeqIdq89aTZM+jcbgRKiilgez3lhnW3BbzFvef9Q9JfroqoU6J7+xpR23GN2dt+w
oRyzu267sKtNflfKbKvW6jw6zbidsGE7zZy6bBzv/D2NF44Rl9fnrqLe1m4k6NFB
Ug5TdWxvGAmOknSO7lj+zW+akE5Uy5WEXRroQyK5m24L4cwNsefFnKO9JWi+QmWL
slqhj+rtV4nbtR0WuPeVOHRDCP1YhzP+Dj5TVHU9/+dujegJw3q2vVeg/9AR0p0c
1Ll/ozuT7GJ/xzrdv9jq8SPK8SGTcPKg2qr/fD8hox3o9Yjp7MIUvlWRomOk/6pE
U1wpDthRW92xUVZa3o7JYDismB+iF31U4YsoKLyvdJZDkfiKdQLLNYZzvCUBKAdW
cu8UzhvLERpJgbRreYbN6B0Odevm4Fu6YnLy2hip/QhOR1v7Eh7B311zvUMiPCcD
+mo3zg+iaY9PpuebYWtYFC2hJws4K0JgG4Vo00zhW19kZDcFhkXIkjusy1bI1BOb
fqsYeFY6mXaoJrzfy/vEqnXKmwSGBWJzR72k+KtpLZ8YLqwPAoiSqcstabkEniwN
HANSRpFvmsDbKTKgIbMzGXOlRFiiwpO23Hk4jn8XjW8r2yU3HAOlg39UytdNccpm
sAyOrlwvf0ENsHZt1v1ZOuymF4LqH+GnWQV1oXRdOzdzQcudCjpdrLE3f68FJtCE
wfhxvNG9xCKpcrjTzGpDxaQg15Li2z5LIC/bg8VK4ymFBoy2jtg61L/Hi5qjLo9v
kieS7Y9yI7/tyB8X18UogGw4Sy5iN/fivKX/ahv9HEE28WXysXctY03aGV3au5F6
4qPNuJ+cm3iRj7ilCQ6yP7780ob+LLEUeNCm22r3xR//NDrhqdwl50ISq0AUF2EZ
jdqQWsKea7xuGz2/JsJGI0vIhR9gMERxJfeKG0s1/GkVHH92QAxe0Q+NQEd7QM2D
PywZ0SQ5MILO9mTV5FctK5zMT7SbAIyo3QBkceRbPBph/wtkVSFv7Mhu6ii6I0sp
E1ZPd3qKWAvS9RmThejdPiAa8u2uqBZQFolDwaORGzITuycp/7/6o7WdcH/Th0yx
vmAiXodiMDJW9Lqf1Et1yeNEzmLoEpjyCM8ddyWUoJ/rFm2SXDbIiPG/Nx7G45dO
+9u2UViNzyMvRC3ntui8MXeiYZm2wt8g3qDpgXsr8gw8eRtwte/F+RlcyIeg9386
nRjpCgy4gzm8XZ29PpqDhoWtC3uCTQJ0KY70sGa29R7B1LzVE3Qy15u8OZIioNIu
8UUGGlAvig3YFesTWsA7TEcdPH+RJJcpukxIXsKiA2ZlREzB1ZY/Vby2Sdp2bEWK
RWk4m0Vq6bl1obyjZBVzKp687oyY3c1e2FfijaH4CWmWPbZKZFsIwvpyRRuEkpbW
cim0MXF1kcVygwGFf3k/7XDnxY6oc55UHk1TFz9+uuDYZBsIE16QJzrNObAydYUJ
nPc6aCZSS56VceuMJA9LkfdFx0iDQdaGqBKPtUTIA494/rNxh7/mrMv02UcJwXz8
a9PC/phM6RE40zZH4syaT850uH5a9pMcWRNxWCtn+w5qg2WeMLeuq4uPa78u0Nfd
mtzbEnVItWVgeQm1tK8Ym+aVgVZOORbrY5bG+COl/dNGGe9nEZv8DYhn+hRTTqES
grXSYd4gjG+gnYAgDLHFaNHSqOH+RiCuseAuX97EQL4VoE+TT7VvN1pkqZg90lmr
RYsEkHQ8Jms3tVlu8sWxRaidN/XpEpJQBTaVw3+Pb/5IFfZ3U3X6YaoCJrtg38gs
q27v7weagXV6B+tQwYRImBGVqq4O0NtYUhlTT/NCasTzj3jkYE/qzzoKgzh/Z/6b
0JKIGlMI7DiwwvLSt/eXvwYCCDESXNqnfvRC5Ef32TWkfUoyaKCu0NhWU7zLfIs6
csUVjVIShJKSkpbU1iopPc9wPp3IK8RMlTYbts3PQLpLddBeQ3m0r5VxTZYKs3xX
MpNjO3yh7orfwwPW4WX9f5nChcg39d7r3kRjLRjnWIjvaDeIop0gcTDKcjZ2iYGI
/g1gYQCjq0Zo1yP/fYkmwz+nWeCrTnWPMZ0ZJxDTvxR8Lh23YaQqvUreP8DWYFm1
JfsZRGkamyWP0T3Ahiv1DbqE5to+Dwlfxup38yAe3Y8YJK3WjN7nSE3xwcCSRT0l
1MOwU1FT6aScVwfnIEgWqHLDeJVCUNJAwHv77bxxvzsLovMWPdVN03wNpywbrEhV
tNsCA1j+hlLgHJlqBo02IiLWch/QLcIUz/K1Uf+EY/018B0oPC2y75Z/W26tIYGx
g+QlGl/4ICncfUVTVuIlKVbD+sQoJBPBY83VLV95STmzDfZBWAA1eXsXJdEMSnYK
GD1bthUziYO9JXaVkrGGbxJqgsFzpJ7RZoiVdNjtBNhkmBUvDRHWeTBYDsQ4IuGx
Ye+uEqoBw5uo0GyMhbGqAks/BAuEzBj96nEeYNJ+R7iBYd2q3ACBbtZRHz9IvHj+
dfoDONMurRepY+3UmbNWEQTMzgbUdvaNk1873KBv59x6lh08QMu9aENfLtdTI9ug
uCOxVC1ErRyjoTSLeJC0PM2QHFCciorCuqE1b5FSZPRgPmlbIyU2L7zGSNhhu6Am
F8qdGHurHwI+l3gWKBOmy40u4qxkVt6FiPReQFrm1wwLKFIOvR36K22ZVDBtij3B
jnU0Eru5zVw8IiuPTpAlSK31f4GRafBHHXHqia9tH/DQi0tKc5+zNEuvZIHMoFwL
2/xsGKsVWpKXoAsEC7P2R5AgMN1ulN0Sd/h4vVcjCXBDdqObesrsawAyYS524Elk
rB/YDMgl4nQgySOvuVg3eH7CSiJqzEojmc64pQo/wyJQYRN5YLfSTScCiHo9MsXD
sGkXg8WYbDo9bvSWgzgKMI0t27pZEdWKiFqIMutvmQYKD3e60CgEbIeH+kPvj82v
Zu7jQLgEGjAasWRbI+wAk7lvoZHLoUIguBrvywR4LbRUori5Pa1b1+7FK2SnSl42
kD6O5lpJdTGf9a9o/jifVT+pODm6I5VzjtIL260eZVQZ1vtXlIOlCqW4xrlnGc+U
3k3GcyvA93uV/p9jR1Oy18ajvGqKL/u1sqc9x1vnf2l6dml8VZZlQtMn8xPbK+xg
ET/yeBxdgAPj0Fql3ouT+U22Rymif+txyKJKaJHvMkMPjvsUo3b3sgeed9W/c48X
LhVIfrxmaWlVok1buxOQMl7mvNhsMjjRhJtoZuizEG3K8Arqc6W5JjeuRR5pBQiq
7SUe23bFtO2sh5bypKkWcFbEPmYwnpq856res+mo/MB2q4JVUHuTdivrilptOfer
9o0SHSIGjP4Ta5CL2aBMRCPVqt8+OwNSz3e8UQx5ufW+7fpKR4JfEt1k09fGg5oS
Xlnw+vCej6ltCNzc4U7c3MNx4bVb7dpHK1/gv2PRb1L2v5NkB65BxTgBMk7uvZGZ
55VWhKKxjGMl0aQqGSjn7+fN2jonRD2WVfBCeD1yAbFg7mAgEciNjJRSdcmj3+3o
kOKkgLcHA4qpqr6py76CfE7YDHYSgpq9fxSQQsZBRC4ZXU9E7AUEbOhT0Y8BDJJ2
eslAOZtL/eoYnIdchRu4fx+1UOGmtNPhiOfdVVGPfx+OIg0oAI9q8l8h9brOrUvz
bF63reIfhh/Xha+vZFQzoGbo1+yKxZ270kN7crNwfn7reTK80C78wXbKAGQ861eO
w44kPY54yhTCVIWTKhpMEiHJINbTwrI/gO3zZbXOLYN52iMXcVwHaDDrvA6+SMDN
fSU0bCUm2ajJFZE9MJL/IiSgpzNC20nl/6/1g0WdOsPvcv+gk70ic+AR2/Rp3eWl
9zLtoVGVgc5GREq3j4JLdZaXkfCx4v46QC6rs1LHxxSHVXbMCNMgpR4kF4FBeG40
B/J1zQCubNQmBYedQzwZpVZn+gB/Z8VBVFEl3BFT5E4TWilO7NGFcDLKwAGXVyLm
Y6YWZx/ASiVTwwmLbkZIV25BMqxYqqceL8lJ89RzWWVYQ4vDbolXNOl2jUSwenqM
vfbiBkqO88VYqGZHyBg5MeD090aydoY7ju73SRpXgGOyhLDwrleIxZq3vfSiJsPL
GmqNz7suqSKGqBKxnfZxnYmHgWvCHrnLPZ9Midbu1Kf3w6wQvA42kzESoPfy6FIX
dg0blUVbH894xJ6VNkMUbwyF58WnSHQPYwcYrdFZldzYSreMfcGHnrPyfHMiPGg9
bnd0w8gMU6KikjzCm2tbodPMWN+yKK4jcgugja4T05IGZdwWwmT9mjbQPK4lpHto
J8siEuXBEqwDhNKGNZc+CKaHS0X5jZlzct2KRmZ1GVu6DFS10f7FYTN/YB9M+zjo
rhX5/NLCl7/S/HRwfC1KyMEQefAiXUL3zixIU2qCNVA4fzYEG1aor1rDTmrU6KQU
cP9KcVxIA/2vqt5O9gAy/M4+cmSmAxmAZJUJDNZjr4jz5fcYFWT6pgPujDpqQ40L
FZnCxFznfDy1A6FSPh4gIlCdfGkkGdRNgGy1dqp3D2vXDmm9Qhg5uZkCTxSE1uMX
uJAs+lyKHaX1JYMeGXkRhhFDpob9O77awILZjYTohS6GWc9HYzjOQg7y1OTALldu
mW3nM6ZT1k1KQ2NZJY1XPuVmUvgc1txFUDpdrSux5iZshQdJfrnJa/+q0zI+Dj8h
BtiChkPnUD6yLe1V8kHPBePpUQSiyYXEXxBSHGCpdhCK0zs5gFwPxVIrpNqZH5gL
OIdxhT7PZIR0wV8WD8qoUA0uwICnovvEz8D52n9lfE1lxSRjiM/52TbrTwbJrWgn
9EAEGdYoyArz+wAifw3TCCkMkRP5PRnPdCISwP6uWDbh/xc2yY+Leww8+zI/dFTj
sC3v88Mxc6vKaozSeWoRFn4UGIMwDycFI8r7+aZ+YFkBtH8ve2iED4j0YrIYEAFl
CNBFXHSJM9UBh0Lqj4FsVMA6EdJzMRl2Yx0LQzTic+p15Pcf5dfCr44l1xd0sekh
pEeeLq+76dH3bZLEakADrWF99frWs/hhwOe8pjD5MlqLCacxMUDeOs4UPZzJOiDy
YHpcfM3imXG9u4KRkLJQBb+qajs67GoUQ7P8UddlbQwsWGCCfk0N+bsgHZqAImmM
jdynGaQY1S5LUgid2oqUDtWbfs19AdKEiuCRx4T1MUUPvGZik3a5N/BnNbQLAwRa
e4vW3VQZY23+Gb5F8RLWu0rNR9SZtes8IAVUNK7Rr0doez2cxIAdjC/2OPzfOzn7
oR8Yng4riCtln+Lt5j6eIHGdehpc2sHHpzO2B68bbU/hNo19o7dlRC0IJAIiFZxe
Qt0yvcrE0sn9kPh23V1akXaX1V1bI0L3IfNqN1jUtlYlntaBeBe8rK13P94Jggv5
MPw+I7HkAhBDzydpP+uaB90i7gjBw1WOeG3frPSyVk7P4rV1lSwidWvWWmijsVtJ
Gli6bseil863N1JoJm/2+4ZD5X88oVM+1C6435138h1oWYarQyhucU2sVpYcW9WB
cPI7HALlb5XOfUqM6BOWa/ivWb2Za7ue+hj0BNMHbvq/KSOCD9a4iaM6xqmjr2s3
zyBQs+17twZBUZ2ZvL5Qy+ph3O+sUwS3iEeTanegJ/abdqc+pcuynucK4n/PFJm1
x/4k3JVzmIJPGPw7hhheir3yaSCYgsMm6IZCmhUIcNFh9MYcih3OVE3RR4CKP/1h
4s5os2w87jOiyov/lBdUvdLpZiFq/PfJJBRommDMZ4sO5HmLW94zfJ/UCjfNmiuf
Ta9vg+aaoPDKnCYa2ax83RfmTG7mqfVlCQjR0wadKUIe/9QPshSV0IANPeBX91Jg
FmLSyVtE8RYEEKzZ6sdcL1ODyLGKN0OqshxEegRiWwVuvSTlOQIwjAUr1penWU8L
tkJH/HTmTHX+3xNkshB5UZT60E54qfJQmOYfE8NzC6yDLsMqWc3dG2ky0QK3gVqw
ddXrQUQM9d75dz3vnd6XSznHasrSpAwxogQv11ibvobdasIUjVgnuYeBnEoH3cnq
HHd+fAYzxWSlTQ/wo01WcS7D/0SqiiQQeR6NOVg4pKK34Mg1+InD1jnEYxqb0gpt
vqECfmFSoI9RnKwi35ptDaCXSsulpwdz/UYCKU5+EXczRooMFmJnHeAY/+emiU7t
zHtZcNg2DtZpvvG0Djlypx5ZSYWR3pZttblvxW3yOxF8VNlFADO7q/ZL8sE6Ry8/
//v0CGikY+KCDHH2kIPDbNq4+WEYaQ8UNOz76ImyKPbklfUPOo3/IK0Fiw2SftKi
66CGu0Sl7cv51edIm6G6CzUK1N+NPSra9BTQa7X/bIMT8WgzThROC04OWpqiacNG
kQUw6jZrCArdDxMyKULEWAF76Xf1vQa7vWgpwRJHdMjdV+Ba/AwG600Ju8/674SX
hgALMO24RTKUuzRB3JossKVMI6M7vOP43SwmR1Dd/NUSX81R/y7UWS6zkNZ9vjG0
FL1qlwPVb+zXYtfEQNVoHWOd+4CEjB24kLvvljlQ/z++NYJPYFzSeWOyNM1i+Q28
RjLi/2FcTFpDp+pvyTBL3TCnsBi3FCRIKRo+lmD7ES76/IABwPTLeTk32B23dlKD
rDSdTYjzeJyozgRH7jfamSpYLMa7HErmkRR0RXgd3yRA5XKHpzHsPsR29pSlNBJT
oQLLHQ+vLV5MYM1APWcWFvRuEDzwwdu5gLNNZnPZ86/TQpKcKIgvVpJ/baUQIALK
+/ZKqJdq/GHGHBfNWswGWM7IY83oD9vRr6PNtN3ys6NhMeTKCada/kVz6Fug/v1R
cbol19OsnwjaRgBgFMO+2rCGqWQ4aiTiMDDO4u9wT+ffKBFTPOw5HKI0Gdza6vFw
2d/SWCMsU/ehDNkj+My8FKLrNiBoPh77lmbA7d2UVJ6o9iBd90pZJ1+f9F2B55GK
52NjTvQWLMCz2NfNNAVKq6LXVePwpebvP1V1VKlCXlzn8nWAdE8k1aVdpzwMIR5m
/ZOegmd/kStlsrPHEnLYWnM67wufK8Yq1HQlNrHSEP5RyM2nnXWHiIVzZYjo4/ni
5SLibmzoUodXZrMHX4TZVNl0VQIx3mFtp2ch5sAyPNBEpEPvUkBnzejb/QaOtGSE
MDM4/wynRaExPEiXdgXdt3idZ0y+fRCSOVvhCJEfpqqrX9a4JXbdq8bXaKkxnoej
XxgwzMaPMW3p5cjJvjKeKT0uiOPo1HngYSB6EY5H7FzoYsLqNNBkFfrOO8/Xku8/
rce6Mqh3b4tIDBuiIDhY24wZqk6WxCEg75YnPp012CyWBwGNFH36eHm7dvRV0UTA
74GqB8uwvIrTMmvtMXjkNWlxr/HGFLVqzvF5urmRXbexY7PqDKvm/J8w/F9FrZq8
jbK74UFFnQXwbdV8SnSVADg57xV6mjB2fHhNU1hZpmy7kZNU5tdnJzDbc+Hym93g
K5heg89tgjIrbA0g4AIk1du0KERpy1nIOP0QDZSk4csZq89R4nfPlDQgyDLxoe3b
2iRAlwKZ7vYePJdRHGTKBV34pdHr6K/sWy7dp9orETli+mPGfgPDBdavibJ+PH0h
jxoJQb9jNYkJhCc0bcKWce/k6fEIyOjiNsoWGt+XFK4sA0/DfJqjE4OyEZCjLJih
BN1UyzUZoAKu6F0IfBn4C4o0oM9KRzKVkChO4fLRGoIln/pMUp3ibqjWNnEC1HG1
J+c9QQy53ilSYE3jy3mUvnUEMgRh3uxRoqlHnv1aiLzEINeBJ0DcegeAgowbxQFQ
G6/c428dIYqwMSSd58iZcnz28GuulIcWP8wV+WY7jYCZ4WTy/Odv2kiSfea+9VWT
kTEVDEQbFazDRsWBcFFaIICYYt0I67P5WDpgWLiElyKfTiPF5/MDA4LqPShc1H2d
b98rVLVGBBTDKr+SZhEiZ6KhBAoOu8m5QIiMTjhIz4A5NKF618yIlqUMYtiiBUJt
WWA5Pecp+gQ1FuC/vXXQIsVEbHQ/ESzoJRVMFGfRhiTz7GEK5M5IyYUH34F/Xbrr
6vTf/eWXNaGvYPE5yL51bWOtImsaCk6Yp40HGGopAyzfJHj1WIKO1FbWTrNCDB9p
yrrQXi3wFCnBoeKvuAjJDu+IkDkmnKNWqGku9IAH1qIZBJcfzKkgpeaakiXZocyF
VmaRITDthS8mgCA2IBAysNry9j0NhOyWQT59HW1kdNZwzKfDWw0x1BJ+dkW3ulYF
5SOLoFDmGrJXvlwhap/X69Ku/wzQ2Z4K6+FqRIH0gqJZM/veOhVnfidTjjJOUAKF
WctSjoZOHPXbdxhMLixZ6eh1hMIF0n/zT5TCs8KCNUllPFbxytCMYwzrvxOTU9Of
Y1UiTZ+pgUcUpjRaAoh5CX2+1CCDF+d9OieiI5zQVXG6TrM4xyhDFQPYqlwcKKrW
OJxCYSNU2HFdN5dFNPrFOduBuh4ImDRsK3L+IEvNjuL/5Tc82fJ8W8/rJOQjD08x
G6WBkj1w3vfPUFOYWJ19vRD5vfM+G/QyrDoW5Uo/WkBj8q+2+PFtXGQJKxZfq9Cf
tqrh2eFu/5GuTuo/vxAbuJ6zAVUhhjjEf0JtIJshOK5RNFPNXRxapgPaBIgpg6xN
Su8ePhnXRpq/Qh53s4nwwtoIu/hpOhi7hhR+6uWD4efGoLgUhRgxOWNEeDmotvgE
lgjCYeVGpTKLhTSDwVcOUb94GYgbInjO8nW4ci9/pq7cZI9j2C+9QPSD7bG5KbFe
zf99L1TkB1ZFmuMKceDhn2f2Xi2mkrb42PXgPluMsZrskEo+UKAXG1xUlcrCPDhs
Dt+jeASEzbEC4pP4iaDNPRvPYVu5SuWoVR6hqI0JuxNNeHBCFPFko4X+INkcpjWK
xKn+Kmt//mn9MI5IWyr6adK4ntVEBw64pcw81K///Yd+m/uh9tbH9s7N+a0MQBQv
iarsQEj5GwWykTkcHZIObqd2/ZUU58ikYGP2ZoH7/aaJnZe+ZvkX0G5n037peq/e
TpONMUDwBw/feKy66TplqwqtIVyi1X/s8+pbjJFHvHVa1t3d36drbB41V5ts8K3g
muIc8muGR5zIe8pMUNjX2+ML/pfu5jwruRkqTdB6+HNIWPNN4JDy14hPRskJKCi4
kvPXjVf3N8KpzD/gv7gsTIEfLodXQhtRZHOuC0NzKvhACEChLGLq76uvBqyjdweu
1oXuiVtMP+BmzA6tSseoGilLcxS8f4L6eQwqSVMh5REVos6j8+/HU75iC4w1gMej
n23jtlQ1YqVqibCUS+JVLLTSK6iwNQQFnMqv0BomfA5Vu8RzTJKQ7/2uCGN8Gx6O
JmTH1bqd1NXW1/0Kc12pMXYYWr4gKlmxh/G0z8FVzMLAshjmXCBVY3BKYMcurNmR
rzWQ1kfOxAR1dH7R9NLQuSMgVmJZHuXUuo5OQkI0wC7+rJGfv72mRlGoD2Lj3GXF
OkgY8uRyUZa8guF/kS1ddD27Wwk5NJMvzmLaiKGyAX4gKC0kvPIcSWQBswLzRA7C
kLBnceOnM2U4UB7APGcNc13w4Od1qJ44koKoDrB6gQIPB/c0toYfiBuhytDF2NMG
5p/KuO5qco57J8HrL8Xruhdc9eTiUnCBdvloJ3KWJ80jHJHrO728MonpmFWf8XU4
Ts+iP6jdCbOXrLP2gKQb/X0v+pQanjIhk+ppvw7TX69uUyiWXTupwliCXhW2duS+
qKiXWEr5n4ZqJSk6SywBcHWnJzTuj8KJyTRz99NTlhuemcYHbDhNRz854SnElgIb
YTSSo8dX4C+QeYgH9RX86GsU5WKIo+VQB4IpYhAnnCMN3XuM3JzaWFmw++8IXXvU
LW17KldOGHxsyQhV1dMxjZ9qfF92IzPRF/0LzCF5uSUlY4B1/zv3UrfdjrhmTbOU
BJmeoMgLzlHMOmpoXwBucnqGYMFcx211JecCTr98M7tRwM4d3GK/jpr3BA/9GzId
XxRLh7vrBt6He9ITciXTcWdhZol3FX+gnv14oWaFN4as3/ZPiPwUxajCZMXzT4UD
zsf2A3hnXb/KyJ1Lbv1Qe08xCsF9NgdCZHKTsEYowwy1qU244U9g7G/8LRYRDGYf
vz+fSm/8xKtTqCYbjZ966RBLN1JyqucBRad/cZfeqP7LMw1mfWZNH5pjeE5wZJhs
YwRuZMESkEkWa2csN56P+F46irQGXaWzzzdnspAwcYETf0PVIeyL2SyDcvw+OkRN
BClspS2PpIxi0jue/r2TFutywwlY37raHTmhRW549T/FHt+EaDmEj9tNoYvWvyD7
70dHTnXvYQMOXaq8RBbuHkb+eERy5qVIeINc2vWaIGzeomZgrngWtMo8lPJPj+ov
GDvLqJwBKxogZ7aXdb0FPBtYNRI/7ziKO7TnJ+1X6MBpOn+xjvTvKlQMKLB6DxDZ
8AJEcIrV//gzMnvmxgFZck+GEBNbKcE+dvN71GpPN3Hu9hteCp2sefhHNoYSkiO1
ir5E9bVTVkrnMVEEZK8hcjvpVrwRKb0O+Lou/eqh1K+LYIrD+yQssbefsZ4S6xNY
22AsJOYPv3gVZZ1/KU5yCHSSOwIRH5rbQqRwkU/fF22CFypQyDZfmofgiC8UAl+g
AVLycT8q5LhitmctGiSBnMhQOrTWaYY1VBmBR1SXZ6nvgU8TRLQjolnvgpJTsAdi
ApCRx7TVv7c5I07oeKs3EwHI8JKu4qonwhxQN01DSnnz5ubWLD091jLM901eRS+1
0ISygk4vog67ShSFr1H3BptuWfYWBeiWTAHXESZUdn9QGqXGEd0g7iQ4PjPCWjkI
KEYlfpw/NBq5p3g7nsQ5+Kh9g3/iO/vXhWDcaNJv4tXRmKg5PP9odiEeHx0rYXfz
6FcpLDfZOb1nFFav4GJsgQi1gKtv9OGI5oWVCK/GXftZ5XlFRzpOLgNTKQpmTYQC
UQQZMzQkhv6KaZzwMN9RGFF9gFA1oYfQgUX74WhNoNnyP7Vje4xXvg+q08MJ87E9
/YPFBWwqKiuNRzIzgVBU284l/znoUSERytslQKvTemtxsnjEZzM6zw43/cgsRAiD
L0Ed4s/1my2IeATunRgK0/qIeQiaPiIdJkZUZrx8Yc/LmmRmQBK9iQVmR1Ty4+1H
z3HI3t20dzsTC/2ssa5gYMHMyjTIbKJo2dBfaYoFy7A4aMMRXWE+YyhS6DigEA2b
4kYJjdt/hPPAmM9/CoPIzCEe3wtmQRG9BYRhBCHeZxYRRecpfaFQKAn7PgG2j3Wp
/VHf3cj5CeMpnCe2LJqWs5QM8qrPZaUTCew27s33yVDPez2cydfkjY5o83AlH18d
CyJhYbLmCnPNDqrzfKPyq2R/nvVEWAi/8+PViDysVKH8kMkiw19n//ArjmN63YtK
ESDgOfTQqO8ysRa/KUEkrV6hsgsNEzHcH+2eJc0IzKrtblute6fAbqcjKd0bYAcD
mmAs3iuRMb5UT+3QKuDnguOUtvkdXBWl+hkP13Y+9w4PTMb84fIfvmQFnDafRurV
nTmO904i4lAbZXfc3dqakzNOYtPbIQvo8tjeRFAgD01uelQU6CPG9czziBv5yDSM
fs68dzZ0T7zhKvM0FZdhpdnUeJQHU8tbO14SM220zR+wNtiULUj4UvSGB4AwduEr
+q2M5y9wx+PNFfLAKyXl2W/cHIUrzlPJlQhGw+Lr6hWvZu57MnVUH1w+MeHvijxi
M0B+okn5p/LCtpApBYaVc7RdPu+5Zl/1pEkTuyq8QcJJK5KdSyj6uhYuefTUJ1gv
u5CgBJjgjGOfCOmn1qyoS32Ua9W79ygKvbT5lvKdW/xgLZdPwy3hqvEWpr/Lgjmc
L/7+w6GdfJgy9v4YCCdTbDEdrv2uJoqwwADSf6LGAKO5YYp3pN/Mljd6ro/hG3tJ
NtGnz0NlPh2UdPuW+crxw0OrUEC46KGbOD5a76N+jEKMg6OLNlUvNMyvadzAv2nu
Oui6mwaB+H5/aXJzNk+EdoVtDjp/3Ag3adKCdr/m+t5IaL3bevxG+/hhuj+fJqwo
3ifJ8CfKwLqDyQfzhl3wY0IH6QBYVukJrzGMQ12yN2knOaB55n/9eFlJTkbbZBSH
TIXNMcgU6XRWOHuzuemVGPlPSeYduXCXNWiMbMEk04IOTG4+Bq5bfxfR0kbJtbzL
U59ac1Gu27Dcd+HuFYGejIcprkoZ5okxT3LwFcXx0lewBeHWJDnXb1AYo91mxWtn
SNkIRA01tQc/e3ASK+gAw0DbVxcc+6pEJzeNtpPERtRyC1NjJrZTtfbGMnQbrP8h
NMRoZnGvpS5qhkf0+UOGmOhr4H8Diy4RyuKOf+vEyGzGa18zSLHdznao3XRjZgcs
aNqqXGvGLrvbqg7eExa/FBPwxf3GfpOw5aoJ3PqWbTgWflka0KrbBtVE+kkMOJ9u
UwJe/uig1zS23OiLgxYUYA5SSc21QlYUPt86CpVdI6hszUDGttasHc6obWrKvJMo
rswa5L+BT/xfXzyKKrZG10sTBnAUci1lKmnDUHuOOLS2mrL3046lNwv/YUVcQ41d
+57pCTzHsgXMImJ/m18EVEgqhzwPOXEBMQ2FOuTA6XsEi4VelWHblWWbOaW2irnT
UoHEwMOCrKqAa4WOpYYhKjAXnyrOfu8EhBbRSYdiYm8DhDGlTwpaypMyvqSdY7Mo
o8CdedAP+H8mEJkwJmc/FkjN6Zw16iQUPVxBajv48Ul1J4jYlCEtNm+IDbSx2ERt
ihEOMO/NwB/J2WWmpeEhdsiZpn0iobaGCW9tVIUcIiJ0C2hhZB9dHsLNydtxXGU6
e1RzqCNrdyhAnlOPAwn0Bafn9tlf93JXFYRSxs+VbIB8csITonN+cgvfF3B3ZHLE
ArnEacPxoYUyrJnZLXVffTdQDnFp6al1CzI0ryOdsQOyRmHUnBIgeTDC7gpI33Do
SYPp7IHeuXqEw0STL+BRHggRxvW07ngBB6XfphLohbrEg5oOZmQiUY73R9x2hpZS
hOJS3O/tQE6632Wzk1GMIrzWrxVW5W+2U30dCGYlI76q9K9luIBOy3D6QqMBSiZ8
LpAxLOfZ2LONpjXQiLUeyU2QvcSa8+l7OOdxoovKILGhLgUIAnnIpTO97t4raHJr
ArMTTrBMpEMuwGvSH0NXIg1bPEKGP85u+5pRe3IljEBF9FrYcvR4bGgO6o8Beo9b
8eWxvouJpdgEZ9dJX9+sttDwbHZFgf/7748xPIFvx6tcMDYPDTtldHEApsIr3X0Y
6uUYf1cfgSoZPBTFWTpzsJFWoWCOC3aqTwDLrOOqGQBkgrciYnLI7jAXFLdErBMX
kmy8klLPH+zWgR58h6l820IFhj7MdQjxwyi13eI5balK17nZ11qhL8R5N6A66sNz
/thbplLwnFyg0ZYpM6nWSTP28zfwXF3a/C2wD580n7d25irMmmpL8MxqopLmrS8M
dbE4YTFWmTzZOUeZpZdB1ANq6L8LL7/hVGX5PmBZDI34wuYwhsfOHSp3p3p2GmNE
ylVF6Tvj8Cd+jr6famfJVH9Mo4ar0fXwuxITDihIEjjX777UIco8CV3bxbFQnr9+
Av6wTQzWJZFhVs6SH13FVgoqp4QNohv70qFcayXG7VHNRsbw4NtrQ+1IYH/BO+ZQ
rcAlvqLmYD0VT5TMIi4U6l1isl1PrsZUuWu8QQzLfJmT9IQNWIn0XgsSseeyLGVg
54HGf8kXV8Cbybr++4qlBAWC6nP5/Xarhr7oaCY2U2dSqHKrb9HGw1+TpMsW39Lh
fbJa2kpRMKzohVpmot/7MtOfnBEM03kvt6NekxdDhVzal6bcbTNcvmj5r1sZtCsX
Bp1iT6oN9nKw1wwAiJUbOSSsi7DESSh0XccAjJX9FhjicV3b0gq/HRsV6Hlx9Fr9
ejSraIVkFBoQJJvxfduatP1M1MkbCfoPEkuChBY1PUeZFwoUOofM/z5W37sqLiik
K/ONjQbeEkCSxtBcpwU966GUNJM3HdMy4J2Go7BFldkVoEouHNgjIyFVDlGL/G16
G6nde6c9WrE7Jj/HMSc4fPjpEQx4P1A50myH9WUIPfgiUEF/KCxm2r0qWgTSZr5z
Af3UbzUJ2j2y/X4N6Oqf/Kh3hgCK/Uo+iLZihlP15pYzjtJTvbaUugsw1OCQ2XHZ
yJMe0rdEf0pQ12+U6J6nA1Fp3YfWmac+jhozmlpr3mpXh/G7q3Q9GnKu15TnR8Lx
5DC2h36j14Kcs8RiBmMOyoflIiTWWA0sEh59SXAqA9pnMfFeW0vsRm1ioA1wFpGp
U5mNABtY8OooAfNzw76as0C1DIzJo8u6LDr5MOngsZWPxkgoryEhmwxpqRSb/mnO
SDhmW3UhzuOQcRhXCXzsGFhOjMIXdssH2BInR/8TvNkD7dPyC3bTKQORTP2iW1Bp
6scJTmbYh7R0gBG+MfIa2QhleygDcm6wTgaPzlVuiBdbqXoRO8EU//wrrRvvHJWy
N+aCglAg6KHvRjQPOqirUR6EJi9qkdRCP+Jt0toWMRK1yphGl3VSlvf2Ma3TI9A2
RkASrUwMWuZjcgQBh8iAQEhnqB08ELV7I3VUroj8GHzkXf8NuApQL1zORWYtQdH8
dU5btNrJvhbWajm4Guu8xu6SsFeoK2HVyFgkK2c7VPwICph9JUBskdWDLo/oWTgh
miRs+xWo/Pj7xb+eMkuv9mOsjsuPgJhCA2r1gMs4ET3YUFYziCsIA9twnOeCVfyG
vOgv0SwwskVqLL3dd0Foe2614BUkUz3Q+NPo9+PicmmpWjSPTA2iSDxRbpqNRmEA
5VUU0KG+r1l/xCbQcs3T47UC63gYHL0JdU+MGRfn044iNHYrYgeH7ZCr7Oh+dff1
YOB9CVMRZhEfKPe2+Rn4y2sZsF3H8cf41cKDlrhaJxeLJe7yfHUjC5PF6azSoYcL
mJPk126ZRcZq1+DjWx7mHJRuwF9cdpplffTGuEAthk0f7xf7N5wpS5dNCH3r1bG3
wiBNiKkmszNISydgOonyxOhNTgv+YQsIMXBQsnGw7kE2Pf6F9wTLTXCqSO7HPGT0
Vc9gNOGmGoKCzzjeeyp5RJASeKyik3nD28tkSCWjv1lRbRjlklFFGBuKICb4ax2b
qYNL4/rT8ggHBDw+rdsIj5R2r6q7Lkl59OLBlLnQcrf8Pee8fn0UqplXz9aPiqlk
M4fMXwp6uH1pNU7NF04zCNoGzBNud2/uWFcreBUImuab2VaeVz7AWa/LmIDheeh1
0e4ZuNvYJlSqJGxT1u3KHjKr2fHhf2mgJ3PJ2zi8vW6Wh2jHts4zKWAbPQ8Y4zBe
Rqz6AJZLhanOcI+DxiQHDK9pFkaIZPjaBGrKNT8PwPfM4shCNVB3vb/8MG6iP0KU
n1yOAIU4rj/B4ATjuz3NT18O2ZufbAT2lNxP5e67mOQBomeb+C5FgyzRQJPKhBr2
cm2To3hPeE8O1UCWZzSsWVzCkW5JnKKmE4q5j94AT56mJzSJrB88dpCmPFUDTEOO
CagD/bnuP2cZ95c8plMrrGktWsBhgO9YHWlhKUDHQNzWse/FUskNaK92ImkUQVUc
kcCOLaJ5YLkFCy/hyODVFJh9ooW7jHlC+Y1aUMbuuIRERwxB6Jfn+e8qsibJCaey
75ZUKSMcWCZR9daEvpU94ljE44TtQ6SSJc7xoOag4tAvcbigrj8AICex/vkQ/B2l
8UNzs9syVC3BQgPofv8B2dhEdJ/zaGECY6bdRyvPPSV6W3C4yPI0at9v3kP4+Z8H
WlGWXn1LO7h+mCcaks5EAbayo96DxDF/l2ahZ8lXUhaWlJPvfLxc4C+wKyHFywC+
D8wY1MMyUK+Qs/Zi3Hsinnw2RlZtJOLMPvylFnYc8w4/wmrcPP+E+DSpJwaRK1FV
TXExAT9UuvW2r/WafEUCrCR2MUMEcs+3Qp1U8nrSD930D4vSPrfoidbCy/r4DRH8
tFCxcP/ucY7XLxGufj4uLTJI2oUsjjgRuUFHjkwMuh+cewsm44OY/sncACkBBiCx
MpFyUn2s/PH2JZqWBPA4oDzuAjLcL0kfvS7qEazW6Ry12ZIuwMY0YJT1ObVSFKSg
y+KUHHxu3GLyRVAerFmyz0hPc2VJhr+Rjy4lRfXi5l1Let7Qi05AbsQ/LTpYkM0L
3+oIox5zTdrvTnNOzFvgqxSpB6+udG871vUYW2it/sm1ceQb0LDX1q7L7hSrWVYr
dMA9EnkeMrcbOqO8eRHt3xrS9zWvqmwiLSupHPr5ZSAFUBI4Ls7dpt5CzGSfzOzM
WSun1MFXBhwe+X3fg5Q4lWVp/QrMb2OWeXVcnBdnfUO/FOK2OlrllBIqyHzEr1BU
AaV8s1s+CPNnnhiPKngd+bn2S+QaNui3IZ6hPHMYXSZ6g+vIVpErnclGyK1n13vX
4WVdP7qh6ZzFa7dFNY46k5Sh0zRSCvfzbVj7YDwPJmYpsB2SA0JHpfJwJbBOsDOT
qpLwcOnci7DBYfNM0VXMxGCEdQzGkwuXf5n18Nzn3BPlfQfYkrsgfDp37P1I31Kz
wY2KVAMhEfnysb8+SNzFZWt2v1ne7bq/MJo0sDykuVYhfcXXZQ0m8e3RO9vydh1q
T89OuNhX83qCMLVm2YTNP2fClwVBzBQU/EctkZyGR0i4C7MrNbnILqgf5nVJ1qGN
28YBkynyYgmctX5+bUI4QJc00lGt9JbubTJwvYnSjs69LGmJ4B9tsaauMZ1Q826f
p7khPMsu6dkJR0qL4yOxhfD5FsYb4/I/39gJ+p+c+ZOCAeKqtC51cY8Sp8tM0PWX
DpVXb4dttf/RFxvJZRSPk4i9V0j9PJDaVpS0tk0iD1nMkbWhsKvYljDJoTVjbNCf
n1kB6mXA8D9MzLXG01rQwpZ3eyU4XLZAfPaQW9jmCSWAn5KkewUqTtYOkHEV7vgC
+USS5+c1/dywapYIdsypU5ygwxKoukgPwcMXQMtLb05o1qZ6W7p4ige0JHVf/v7v
nLl2bXoX4W/vzJdACpvrtYj/K4wIIP3Z6s/g+TvPeEdYuRmgSUh8/dbk2UT7Lkb8
qUXBQ+pINBbBOfVy+Q4aoIBMtAKplkeHtU8MPjoTIZCkcIa1SxLmI2nopSNubH6R
OGRzH9eWVzNMhBUL8c4Y+KkYWd5hQ3slA/pTBpNGBP8kILBbCLlwmOeJMzbBCfxt
iMa3Im0W1hGwET3GvuF6cTspiyALdZGuyp9Y33gLPne8GY//Xxy/aiEwImb/IKL+
EmCfmCq5DNdaFZY8ErpUyqxYx04d3Gsh3wxWZu6omHF37upB/KwyGKk9NDPckCUv
yxq2bxedbkopI6lKZwlFWlxQ6xcQzMtJ6H1U/5ZF3bx0uBRO8pyBSW9MwzNF9++q
QbTTm2bxCwxiq4kWvlonKrcs8weicizdB5gh4CCRzp5CmnE4FWZyjoTXgYWpkcF7
lbhYTYaqSR4lzX3laytB8mvHMNgmnvJ9a9j2XH82RESUSDAv5IKAkrPm4JK4s9JF
ER75owgwhY4J1woGUCv9T4MNkmQNSRUH5WvOnAwpRp5x9hlo1//S49NvUZQnACxW
eSsC98bgWCvv2KwL+I4r8YVcJYTz3zwk/uDK5W0LjeVdQYZC6nH4pIrmK961pbU8
XJ2LM6116aKDwGPSIZxsT829TyMGLtrTWLIOm9SuYovVI/dfxRasrAp3o/zXPPsa
4LtWiBoBGFqm/b36nzwQcEqzvrX8S5Bcxtk6qNJL0CEAlxSd+97xuGMXg938LXty
mDgcXBVf8G4iFEfebIHjFZ3JuB1y7axnVUBi4+VXbw9nJFzbOlljYKTdtOQ7bkF3
AMmfkQgQeaIX+J2bRaffOMV0xE/voHLsogeLoexk4i+IKylawf5LRyIbxjFqHbF0
ob+vuqZn25WaFMywIEN/RzqqMBHijDj5LdIR3h7LHSd4OaSVB0HHro2XKWPHktEW
CiJc0uWN0l4jxf23W0M3GLEqylkKrRUQ5On1jgBCeWPqgLBJgcJSKAiZvadk2CD/
bJolu3QdTK4fdoSvRxu8hzpaVLHhDTikZ01YsSjugBBBqNiSz02jGE3A1bjdNyBc
YOfF3o9iOKSD2t6GF5Kwwc4OyZiDFffRIde3wgnnl9QuSqN+BHjlFyq82IReUbra
yFgreBNTetFCOE9w4T6nl9QxuObmubjf2xywy9HokaxGoZEtMj3tocHG2rTNgIeO
3HIj9ppLjdILVhRFZTP4912uJPqlgjqB14kn6uRZhlyB/gjjbgC5MSXPHETVz0kt
rHmh23t0ZgMypdLJt6+HJ9nu0gr/G3JbnMbakgOoOolLRLvoMrK3OV1hqgiOcMYs
wVeRwB/wLSHzIhwM9BS4Pfwj4MZpULCQisZTbkyFWMkdLy4mZnlCQgjkb5op10uR
FPuATJuEuvWU+LoKvrx9h1DlUsEgXHj4/t8NcRrs2FnjHEPVgFbA9ly7waJmurhs
A+oW7Dt6vj6AOI58MjZl0GUF7cnigNUFPLzZd1Sb7XD4bTiWYCLZGncNvBH038VX
ZNeBlCWHmZB69z98EhtI+mmVmw4hBaYQnzO83YHBB3JPA1jTHDo+KcedsG9E06sg
3vveKOSYbwfU7M3kIuY+ACmdK2qQRj0GKgTfiOzFzReMHoGIbuM+UfXsITSi9ekW
wE/oj/TP2wDifEC733W4BZC+dUSAzg4rlrRgBFlMsN/fZ3h22CbnQovmSQWLol+U
fqhOngCaRePq54gbDq+RuHh8qHz7wWhiYB5hdAGPMolOvhDigltHnjeHSZ+3Skdv
i93E9DeWQs8niCquRQC0KWnePM8Y6qfNNmSTK0nLb74jXu7+BrkzCTlhRUOLcAb9
OKkAa/ITQo9i3QWidtmgMrcW4JE/GM4Q43okK72MRGCbcly4NHjoqxJFZcaH3+ih
hwW123DgYh2x6J7yR8x8JQ6q4q/A3dIFiILkrJ/SzpGnMhGSnIALcQA9PWU3OUUT
9nulnuX2Z4Ufe24ojIkuISIxSei4nx9oXGVbFmq19F4jjT7R/I6gkbAsdMhj3BEm
9/sQ6nHLGTuYDamwT9O5SEG0Gpeo8p1CPxLg+v8uFmNG+HiO8SWELY/UXLzcw2oa
8Rxe/EeGc+SnVQ3pbHJW5XZt+1yPU0gwduh89a/vay+EJlgcJoCiovo9izPOz/j8
ceGt4kCy5Vos5N0+9INQvr3GMJXA8wpIWfkErjvI80rVW0twiFxcg6IawO/8XtTI
gTZcShnJycrZkmSkzYZyPHjDRt6qCwi6uv63hprL1LLom4zL0EPrH+alKgke+YRA
hy3XLeDA2nxQGByugLj8hDB2WUk44ZCT4eKegXZ5pRE+309OnfK0DQU39A7uecm8
vl+zpS8HhYZVH4cAvmDR9ftlzMl1pJSxqiKObFZCa1UJO/4ahHXGix+iWtMMLeIL
dmV7yfiX2bcLc6jKmUQigSxeuYJq3geyU7r4K0zwJxplYT/VgHy5LwUDz3P27cSq
ztL/RTVRIL9nLdsoYOcM260hwzKcDTXsJB+w3Dt9ZIv1jPdwGekVWATQhwIWrJlv
csxoeu2IgmRb/g4s5FkvYXAhPyWbOfZVURFVzFTGIn+OPAJs+tAKsHABEFJUUoI6
zbYpZsDNnYnCAPP7eOd0/fdfXoCA3NlexeZOrAdvsKWZaPYhdtxaqBZL9SZ4Xme6
fWp0bb0kSU0MAjBY9+JXb+LCh2gWhPDESk7KQP5FdYFQjBoNoLe5Xte7m7HcWktZ
Rj17wAcoTVgYvrAPsrnolm/tPMUuUu6JsbRkiZ/3LHDr/n4V1SCN4zWR180TBR3/
e3DAn952RLHNJwBHZRbAcxxu3EXx/JNDiQ4nvnP+BVZKKfbLTrwh0jWVQq8Pbjx4
e08hR3fj6+8hH3m9g/Pgt714gkFdx/455MDHa1kMwZbiGChaZW5kK4ePFsish3WT
VLWHW3qUhF1Yc6k2pg8Z2vXmeoa8S9onLdJQ6NKMy4vPg1SkfGvVLJ+lQ5LH49oX
BSaPt3l3hINQ5J6Sllj8s/U31KzLPNfp53HkYHUiIR3vzyAw/O5ER7FvzsYGAKpe
JDA7+0NpWULsDnwhO+4QBR++QjR1un7KkE585RHzEwghnGW/NYsv3rQvOeznCXSY
IBo0mhrCHwLM/Wq0bFiSuDR4+RdaUI77ul4mrPzfarllOwhg4/xrtCoeIn14pKCP
Vv5QJZU1v8boEuDhckyU4t5Nb3jVo/8BFiPQM3IrCbGtkeeEPx10FWdUlpVtonEN
pal3yg8EDNNdTON47OE0eNdbIa9WE2b21tVnnoXup9/X8ePbsIUkQabTX6wcdEuC
/vyB31JB6rm5VVFZnvhELgr5c5X7NDGNdNXE10YumKpdhsUrpgLcrbSeBqLeQNph
ifUtDf6I86Ei0kZtMxVGpGU0ox/SwjNjDgq18HADDIt+nKsX4b+r+tEiaFkVNWbr
5oFbymmAAMiL8JWKaTozINaRTbG4RdLeDxOkFmgRUDWek1qAR9PYkTOVQHkGBhIg
jqyXbrd/8YC3zmwzayqI+gFksnkrlThNFGy+9mtgQm9f8Es6e+3DKHGv9JmIhGbx
PHb86Ouqro2z4NVc/E0jayiRg4AUtZ/QIhS6Sgmxkk4agPbBGeBMZ26Qv7tVVbyv
m6D2FZ0h1ftieWyHz5dibUOfx1ps89a0h2nKbo9xPPtee8CR7b1aXGd9XkpPD13i
daqowMK51Sd0OgCSo+UcgCIYNWe6fV5Ydtm9QOe1q5ixWZ7t5Ur3SDEBdLn0UUNW
Nf5xMo2mm5tkCgOdnSF7P46+4zA0RQHzekb6DVmiGWGouy1LoFCpJ2a/H+vA2dsE
tnPM7JWNat+IhH0ZKoosIBd9aqqmHA+SqQ5db4lBETxdTUud44qW2ebOFcyM/jDC
YkiHwrLEA/pZb9VCMjarpwOtK9jpLqVe+YZPkfeu68VfCNJ8pLYOeX+CV6CdKbd9
1+ui9h/90gLntcOVJXjrPSIfzXIuf8At8IVKkyY2FCfwi4svpnOZoKE3v1O6JMk8
1R430rSoSFctl+0aGWwVxrz8bL+RlqULpfKrOfwyb6MtweUuJGiRgFs1LEqrkAXG
2klhAErq+pxQKD2/pA4ZeMJW8KEs0Ob8rw12T8iM6fAyeEVB8o1bZ0NWaVco+0kB
u8otpTO43/cpGq86jgE46zJ7uSAL+6/dT/sjLgXXK3sYI84NzoL1YnEj/lyAGJ5J
/yqkDHyQntIYqan7VQIBQIE6LwKldXCAWrxdSzCkODMDY3Ci8Tr0ddAHG41fYy4s
2d6lDtCQ7lByns5hBvSZjfPlvholPuY0afFu92+qfrM0U+qNsQlZFyE4B+4IDtSN
zDEdKBuLdxHcs6Jyagal2synERLoXMGR4ssx5IUJnKejGV1paZxItjvrBpksjXpV
JLusVLIY3FMToR6etdTCJapfELc6lIGZ4Qerf181ldJmo8EDj5Lj3Ah9qvELzrW7
2ydBSUJl6QZfn3/7G43h6h/8HmSybzVS3AXD3wh/vqqvhvm1Ha9sjb1eEP1qP5XK
Ju6gGRBunN5nu3OF+e0BgXPz22P6KMfOBdVZ+sk9DG9LvnLcH1K4t3qkM6dufvlN
HIUJqTcd/Va0xuxAEsk8D2aDSJ6Jr0yB1PfGEeFPLVAmd+Lw3yBux6Nn2YYAqB/h
yPm4qeNHMmcObLzAVq2WIHMj9oEgapTHg/43hEKEX8T7U3hR2oGAv7Equ4Q50xdK
dVWI1z0gDvesG9YFjqhlvSzf3L4X16u3dUk6SC5tX2yfdMNCeBOYV3lRaA1UKxfU
tZ/7MM9eK9GVWRrYXjIuHd2xJ9CcpcmOX8kcy8UzWixzrbAqhnBBZWIJrzZpsG/j
X4A6KUGCLE/qxA6v7Cfzmx7PMis05vTgVJp1xHQZK+5Ev28Dx/0fxgBN8Z1/ApO0
HxLVaD9lyHhHGKPd4TdDFnny3c/u7wRtYQPh8MHungbo6g4hEujjMRUBB3GiEEgD
QzHsvxH4fLQo430kepWk/Waw15LzlnaF/4lJj/NqtVqnD2ASSKY0echj8464RMo9
aRyGh4gSsmsZI24K6gd7UQuJn+SRfCjW3uWGwmaFLQpS4stfxBAM78AtXGNtD4N3
I+uvJlVL4pgXWg3Ag3/L5wXwRs0goFkk8p3TxGQHX4XbozLBgKbW7c4dvuN9eMxz
TwWkyOm8vC4Ij6aEpf2HO01Dx/nmkGt5/OtNfQqSk72qNtRBwqlS2KSngISiClr3
XE1qHYmgTtPQ2Mg6IQ7JOEROenWahoMDYSjC9ojfG9tJIzjnczGyy+36jaDuLk54
9KiW7JdFIxnFh7PE870KNCkTkzqiRot6ZzKkz7YYyN31fvG58XvqQnVA5xkoJgrt
dg9B4DKL/xQlxq9ao7mXGgSsr4SXZTyumw2wRO95ga7WhGf/pyXSTTE8LrIYiS9e
0pjykrGZRQEK2/nYGIGrdrIGqYYBTcUz3NKM76nckFqgFCCufQtYdBtvkb9xVj3V
4lvUcVOzRhC96zJtCQSSMfm7G9PDnqaGus+cHtIsaqBxzt52ThXuKJ4TU24bamap
dTHonA/7N2c+phCQ1SaqdIJYQGcU/JJZV2eE6oXpzHtDVRR2yyVbxnriDAHnyBUA
DHu6gnF+4FuVu8v/d9Ty1um5MfoEmlpmAzUf1UlMRHEoCTNH91k6sOiasU2RqBIA
OJ2a/u4iPWBvpNdR1/dRePKTH56OMoLUJ0xn26bHr/DIFH7jTDJAIj9KVBdEjTGw
A7dJfJcZykTs6LyHM2rbo7QAP5bgrwnzmKNbRMvhd+rN3NrSqyZuQRBXrrBTg2Ll
8XjAuOM6wvDnqdJf43H2W+BSIJe5y9x7xyCXDY6Wp+4SfEsbfz66L7LyC1DUwVfq
dtj+rg39iq8fyx3dL+sTNtjlIa3jCy8tPfkA5ZiacUH79m2Gb4S3fIxYFgr0R74M
mI0pNp6ERicCrDSNztRm6Pk7F/8f//Z8+/ak4z+6Y4HXKE5hE2qHoM3lXJjC2Vny
WbsB68YQI5bfT71ZYQzepYgz0uKfISzGuRQMQ/pf2Idaj/QqrPrv2CMpZtUucbcW
2siq0T0dxcy1ggEJ6YnwYqhic8KtsB+iLV102Vw40uV1g56wMIBDi0drTCg8Yg0H
/1RZtlvwaeQoGvnUjf2E6fqubUec3x7Pr75nHFfot+YvRIlnmNOXVdG3ufsLr2lO
yP6XZCtkr7wgGrKFRMKAg9BFiGV9/1gbB46WwjYapt15S8OVdaorOV2u1XmMSUX4
8V4A/2R9ftpC6FpuDxHqYR8mgVake0mn6PtANItRLxoHLFruOIOdL/DHAfuWkGRP
9U0htAb4/g0CPR91fUzNWpi0CcWK0GIl1ddNOLqqeRAF330pl9qTptz9hHSvI8eN
5zPm1GG+/BduobJ+tP2JCGnox0m35LFZOsiEubzZu9KvaNinVNhww/UXcSPRBYxd
mEVMgsZlsImzlArvSEjRPBOPC4NJNqYOjTOFBh/4Rv1XGPWoEcJmdghY7wIo5GGk
UXydwT+p/YK/QxbecRX4X7yYm3FcTywafHSDFuhi3Qqt158wTTJf6Boyr8tcwqC0
SkV7uvuf5bDt62L/7654dwo/mQkAmnQpxPUfrFndEYog72pTkB+pZ5A2zcv50Vvw
C3DOuSyKgPqxBdLxNHEIz8QXVRXKjPbSMLr64RHhvcnPvgI84+U5C7Rea5bttX1d
kBKZDiskEnPVnD3NhkPFhu66aQT0uUI+QHPBuud6BI7mjKn4W2L51btnp+Y8e8WQ
yNuP5qFllN7+2IKCF2QAroZkKcG5a34xeezOff0QZLTmtDdTOVQKhbcRQS2mJnGS
BChFKyaKEzAlKSTZJZtuDG8rCQ1eJf5hyqgeArJ3paTAdR/eq04ye0tyPmWo5fTw
M190p0ehU6P2x9qulZzuwdGA9nRJDFsvd1IhHEtMjrVwOpIcw7fpM7gr81WjofWd
sZkG5xbSRF0dNK18AUxlufTBb3pkDPMYFtmVydUF6cXF4Cvt697DznXRn9A+h6Rz
T50KTUd5B+9aiiWqu9AN9JrRSUHMYKikPRzzmeQ1eVFv21+H+F318Tf67mfsvUDh
abbSdH/xRwu3rhM/8KmObNwsro0I6o9gnC8rUqXg59j4ZCi3QiwJWK3qrZG+qDC0
WVK2GxE+hlLz7ePm81yIs6G+iUAgbidRA7NXdqtEJ4QjYHDi+Rzowu2aQrKvWt4P
yMXjmGACOmjs6hjqz02GXNDCZ7qBUY9WWzJKBnkg0IWPmOpvbbP5wyb6M3Q56Vv4
F/kLl5msmZoTZMcUmWjTLYlu/pcDcTLNjJ5aJs8xxsbUHKXmNcrR7EhL8O0RkG6k
3cKjuQEQ3f6dBZ7X4hFu6RvFcoDmbJTFZiCc+uJnlDotUYFMCZc/GTCMJNghMHn6
zKObz6IubuBuLZGgPl+GPcXYehfgrXrPYiX9Fq2SWJ6mVhEXEtREpdIsCmpaw8tD
Qpg7ls8M4B8WSHwTNgDGuuI7U+sLJ9MGS0vpHdsjF4YLAwtygnMza2PdHfNPH74W
csPwnDEAgaeEjvbmGVRBeDHnLWoYffIIzB9lgPr0OaF47BcXohgIacZoZ8++9w3I
By1zjC4qfPKBMdMSsWBpVlElXi45QTYUwUIMusZ5y+L9lGElN+b8p4Pb/gl10s/6
Ac5K86+laayT0+K/DNuhKSlIMY0yhk4TLY7o+RHUsDyJO5StQeIAG6UCIL6GHwN4
YXSijdGc3th5x7i1MMJsiqYu5atDbtmoPoKi7ITQRK9J1sxK5IGxHd7Oomj6Um4X
hELJ11BZazqRsKRXcK53ZbKFCDA5yBQ+7iZvevdKmgHJVk1oUy0Hxi6VuSD2edcb
yhDUv9hvCk+tJHn6M8DJ6piI4liGrruRUkasREaUVYzlrC6GRgrGHySSE+dadINu
2GB9ULnrybqJDJE7+MYv0weufHsNLcnVpJB6th+XUljmFF/bq/kPwAJgWh2eK9s0
93lRfqK4zSFyFHuI0oDGowjV2LJtd9qWJrFKnczXoT7Alhj2pMsOynYxVryJgXQz
VZltYo7DXS0tjVw1tx+ISxWtlZ/e14XcN/UpeZ91EvX+5I4JENAvNVKKwXUOsrvR
DQUMhzdS4k9Y13YJlBj9RdilWnaN5rIDTI7dQAuakSks2mNeL2yOJ3DZ/us8kWfb
98pjxJxNZJ4Z0Nq8ecJewrQX1qtmleyy7zJAGRNVwmUbPTMBj/3YWwortkhBdySy
s5ejWtlD3RFi3SLqYs//sbrfDgomUp42gV3Rvx1MGOrV0P69jIJuiVD+QA46n/YW
xPNCpu4M8zWmEjoQDJ9eWfqVsAEPh8b5lFeMTAwJOIpr6BCec/tRNpjHtySC3qcW
kZuLWAe1gfXeSfK3aw0OuOEGxoRSD19b48eaeCdc/nGm63lbH688TE6nrwytabuZ
7d+lm07jHrfMES+a1fXPSnTabcQOCKqV3FVApHTxubau8xOd0qXR8Qlcnx3dmXiV
sard/vxbPZCEwneiBjoCTPA/AiCw3cEnyhy5EtvC8D2kMRi0w6/VzpLHTyyhZuMf
V0NztFos4EJS9tPAmlah41V11ftAQ0vE1IaLxMfSnmW/nZNCnxS3OTNqiXtP6Agc
6HfO0DYkC6YczriryrwyLA/5sVJaFWCTk6+KiD/Bbobachmcl0fIb5QDI/7HqOzO
zgA6CC4y0ZpSA6bq8f3u68s3tWL892vhe1D79aJKC3v0low2C8E/EPgG4ndxNSCs
bCpF4xU37kZ9gXJgNO/n4Ia2/8YjYkFB9Yv5zwGphyxujHeG1z7Si2P9or/N72FT
cEQY9PQFHphHIysYUhZiKONc9ngbcsXSqb2o2hnxPE0de/J+7ZS6nKTYw4iymVMj
qfRuUEK3mKSIQK+FBmFf3J2JJLZEL1Q/lxd3stQE1t3+GqVPa1Fj8+JjXP0xY9Gh
rap9G06Wyc5K3oapJHXp2MU2Zg6mciZ8rcN79qDZ7RPFPA4G3d98N3rKA3fst0l9
lXHyeD4yA6vvjy7nCsOJOm04SEPNQoleSLhe7AlpLXQk+mxhN9Ewl+N/m0y8RSNk
qsfuN01zq6cy159W28gFweH+uFxH3WTsx791ZLsbMbMjT1YtW4fspNf5kYfo16GC
z8UHPn/LTqCLUjv4ljzDJN5DfCyBGIUQ88AfoDKwECFin5hBsUQt8YVkwlWHWvGK
Y6kZPxSfjTJHWAgAGBxMLo4h44+D1uXEsfoHrfDpNJvWJFxDwc07c5Xbtj82TTmm
TpUu3OUAVBC4Gh/CLVQr1feCooiCaTr9GYoWqBaltJdaAIgy6UGKsHbkOHoczbs+
pNnpPTyMsDjkAyIf86bOb+0pu7oRzWWNr/yb/EiBEmtcie7L6Y5zNgAWa+BpPjHs
kZGJooOZ9gT1/s5jgKiBGc1hXUJxDmYadML3++fglhrcL5LDzRDB5DFjKbfbxDwY
t4yDrK+smB3kMGYn6whl+u3P3oM/LN3u3CjXHv8oho5qJOtBHzliFHJr7JIWaeRS
wFIgATUmEmtpZyBwas6i4WoGsz56typtKC9kEqN9X3fagilnj03eiDEwFI1uqz4y
oaQx8gUgLY32ADwKbrMo/XplJ4H/Xve80WCQFtg4CoqEjk29/VpggztUxctGo2JO
x8Xt4aDvfPif3r1qwDQyur6lheKPAsFOB8iLralYTOiSTJ0M/NGP1Dqs+8+flz6E
Rvi7kiVpnjHelsiYz/kRrV2d3hD6us//VaA240d5LJ1keJWdEKgDFpPjHI/q3GpO
41RFVj0j7SWHygeSVLaH6s4mOfNV8a50ahifXK3JHrPs4rPqD+Bp60Jkgxd7OZET
e0c3ByNeZfR6uY1RLZXJMOfn2fFPCb4VYsUj3ofYpPr7upWO8/dNA6al9mzTR/T2
a/2Qo/MLqlaWl6YwZZMguhkofXXUmG+c0cToV/4QzkHz/PRkr8ar8XW026HX4mWz
qmGpWXpg+IdfGFyCZj9K9q7MpFTvNGVYh++0ryjBYz7SZ1TspCfahS/KiUQZt2qU
tC9BtXHalagA05IGFhjHNBRDk6Rf//Ai+Vk+oPS49cIodCVNm/gq4khF/hQQGyiP
AzcvKZlY07J7UU40Arqwn0H1CkbpywCbQTWD9e7wPlkGgVZNK6CzIMOW8mg7O6BX
HCDi6Voi7ildg5gU0d8NA7nXbHRS4nLBGRaI/xBGq6+HbK2E23cOaky7lidbssPf
x56bMCnXD1OWJMRUGoUXFMI74oFtHvq8xoOhajkUgQt4LWJD9iFoKBQehBSgMbNF
ktMRSH9fhbMzEjlh5XtdcYX5MsZ3jkQjCH9EGcRuw9KeY28phMWFbetZ3Edfel3/
OltuoBtwCVR6cXW9td5qxaiYLoaW3iXN3Gp4nmRcVEp7JFqR2NtFNHkykt42vK3I
956LQ4qBCM1rIDqy+NwCw1py9SV6hXENX/2aUDwH8Zsc9/2xep9/OBWP1KKjZUJx
0B6iRUIhqcAaNM1ZJlyt+ozKpR2C7MDo7J7CqXdtEWHuwArICwyxm5gZq3pJD1qO
T6JaC7ODSJdSpPi8EIn/08J6z2l0zECYIMGFdSC15EO1/cgr5A1Pw2ig2qS5hUXS
WXQIOf7Tg5H1OPVlL6RBQ6gYCsun/sUWBmB+k1R9gsfEYXBAIa7cZSKWj2bcZFcH
dtnLs/9f7pNLwvx3Se6Jh0xx+/JVtBExshOX6QDkX7sBazQ1xnYTj4t2xQ9+Xsd8
FWCre9sHExhn4z4RJ6Kg0c0sMol99k3gwWLYZJFZ+aFDI/qAOZdwH0Kre31gqqLC
YEEHq8KMcp/9bzkcTpyKe63G4bYhp1B2U/B4uC7d0LQM+ba61HRE/9tav10mgDeZ
ksoHg8sVBoeLs93C+magw5MvWpS8pdlWiSMjFiuBxGeaucg9PLQmKHoPHI62Kzqf
r7SHdp5cm2I2/3glE7H4oXi5lCYH+t2lrB7CHTssTDS39FirXW7KoY7o5wWBkwjx
jdqhZJGWsbgG6Tna9yCc/sT0Lg0m6dXoQEp8DirM4RKXImQOGWEp1kp2jgdq/saN
Bt9N7j44mAjFkIQqXUIU03qDgxYB7kVG8q7wlTh1gkf0wghiJTEL6sgmDembdOn7
y5Tr/NMM94/L1VKKYTIUE7OgWm/xRRdXmk8Wgtk6UKYWkHrilwSLZXqJJX5hKZIB
QRbm9trtnRmdbhFV9mev5qFDlXNllM4SRQVGuxY5Xn872slPKuLgYXGSXUTklux7
N+vpDo5dYL0zAuVWhaVS+DfKdJ3FnZTDkcHrMFISTLejcnqmloXu7KTq6Ke97cyM
iMqFZzr3lclSmBn4ArPUQ7Xj5o9sJpDx/95fl43J/BQ0MPpXLRBZg2xz+2lycUyj
KlAJBGmDMS9e1+9aKG5o3uWiNqlBpIFKuwhWKfb7B5IWIzEI4+Zca/W66C/Z7Qfy
bITvjLqoQncI+Y0chRanMLxXyvE3gX/0UOBknpYgcnqqbusOcYF+mH/1E7DPZ7qS
NaZTVRacquB0uqUMLzl6dM9ZDHX65WUp6DTiu+tqwz2MhUCdjErrDEMaCD9odT9z
EtPdkHf585bcrIQwuz4nhnqA7Bg3Ya4IN6iS8G7Qi5XDPMgPCUrbbJFX6zaacU2+
pIYaHiWPkNYHi/r9sxZW/UWIpU9pd+8dgb9QoUj6o62vphAGn7znKQcBRg1gm7dF
8UB//w9SODbQiR2Yne+n1G2KpBbu4728RTdSIS2q/yYQs+t0NOYyIsdTYdua5Eic
scwvHWnimhDRbSxg2jRrOZ4LcOtDOESkECBzquLx7H4SbO18EZ+aorJL5HVSfEFH
TctzL483BLyXCydWk/ccxSGpB9PW8BSs1XV5qRA1w3iHOoD+6zSJD5bYoq1C3Y4a
Tig2mflHKrhuj96NCsM6NtUVpTK+67eaRyWx4Q+M/5Miu4xbvVDqh//bpAjFiLv4
C4HcAvR1oUKN2olRTdfelSehi2bKgrMe7PoKYzIepe9WKIvMx4xVrmv6FLJYeo37
DoNeyDBzBDmZAIHGB1w+QG47S2dNQ8H0tbiSuLL2SYsKEhEw/6xGeJ2dWnlfdSKl
+HABWlcvzAyWgTgSPNtE6Imw3cegfCU+r9OJvbQRm/oXxmBsM7YATKHwBeRijIu7
7xYXCaGZ1tTk6+fpnntdNchIzvmVIG7uJCkLwgYxCq+7L01MxWZYyUL7N3Gd9dxI
gDiymX8+0AY9dl3Umqq0fudFIyFXxHD9Gl4kdBC9o3ViBCsMTwjEnUF5fDTrFKL8
bsqP+7US6nkD9jkjcRt8DitlvLKxf2qLIBWaGhLvkAM8FOWwkS1A+1yW0uIcq/hh
+ODjLRYzvaVsPbHbYMkNqVSJH5n9vIW2NqBr/1txSNcAbon2rxRzGeoL336UQzXG
wGN8MDgygt1GkJ1akNYBSz9KJ+jG3cO/bxubbdR8ZMFPy0RcNznUZ33bTVlr4Shz
J83L+PQ0KJUN9F0mThdNB//lMHvmpDP+qsTKuV78xRK+LoXKEp0zkhvmNA+V3gjE
uFKbk1piwVeaagPyTLwKRps+q53cuS7u8dA68ewcUYEwnqFqePPKtBRwlyaeQUzj
Ey4ybGJyxlaE9vEFgQ5kI/se7G/fF8+wvW29Ccr7ZDzajFqLBXyIcU22ewOzCpP9
/CGMBgyfpu20jYJ+i5rOo1IeWRzi0nxViP3/L7gwJGOCo0l0A8qtzQlJPOKcBY+1
aLjKc+xLaiuGzDR5553MJX7KE0Sb9v/T3XJWj20UsHJZCjNiIfguIHsRdPkdma21
igLS7kDW6hLdIzEDlUo7JHKODIzSFGs+EBA1ANcCfCX/Dw676GZ0IpiJBXOStFoS
oQ1xPIcvevItQi5ujsPRvIf1yFPRLPQyi3nyvL8lDs2lWw7svYuI4VPSpAliN+MZ
WT8pjp2XtjWeWrPgcZ9O5xe20MyY9ZvM4YWJXHKzA9ACyN0lR52z8GK/pS/SIelm
sJ/LCvu9LEGYoZ14Z5acG+fHg/euofn6lbbPq5m8TgxLbZghjRYEWDM4QT1UyL7S
VPTI6+LM37yovcvBwJaYOJoLa4p2kHveqp8FIo0DKnboGKZuPUNj40WMor6wEJVS
rkgWcvDzXk6Yg2NPzbNiUUVaNar3OWXJ66PH9PSsLp9NHI0U6Txfp8pgOonRNpKL
3ChFDbcF3YywPo07110uteGHFN/Ak32c+3zIys8pdfh6nptzOy1bm2mDIIqZySi1
DE1HjjmRxoRJXs/LiBVuFnXUM2GcXxnkyLItZO094cMl4C7TAZG9EwQbiVW9zrZL
cnSi0FLQFHUx+i0RbqP+MAvTiZsRR50UzjOq/LGFOC0/C5NNVp8pcdF0YC5rsWTh
yxP2umdL90jHcs985Um3u9A2OmMloym77OmiDPKwH8WtRX58grLKp1FpL3na7hui
XOJ1IxsH1j28rGYUI6uQlxUsD7pnrzq1EAZMwcN2Xr/wNP1wIneI7T0nPCjC2Om1
XsYak2IGTvPJzXpEX3RwPQRvs6egih555cb4OXLU7CcqwCyDvOM6/4+LpVM/RhnU
GarPx2vKkPUYtaomw6k3Zgafzsgc5kXGF14vO4Xy6PjHeb1lPg8GE3hLZVZPOaiH
wzKT71+ri3XWRyLEtB5MwdnDVb+UCK9iiezQWGEGEWi1eQCvfPrsY2QzjYT/h+or
M10cH9VJM1i0pU/RHeMLZTk4QXY/kZZdIMxNsH/JhLWe+DsuwGCrQnM3e/pHG+dA
IQcL3FCu6VJPhbtExZLSXf/oSSDXSmxkG3MQaZoUSiN45mls4d8kPoxq16XiScF3
IdrNDiDsmGin7ohSOBr0ByCTZgs/0BaBfq0r7Y3H50sRYfLMTrz6d6pBAPZo7f1H
bV6maQttkRwck4vtnjMmiqvuZk2kfSjHwikcgZEGd2+pS3a/bZUNMjUGMBl7SNOd
3tHm6ZkYbhTAq/sKafrbLnUE1SjB+N0+s2vgjHh72xL2KYXqz9mn7daX6CQmu3il
86PkW31RjVyphiuTy4S4R24SnujXhOghAwa+I8Lb2ffKsmqXck62ASZSjY3hL847
WhLhQjNZn50kbAjpT6/VFfiOodGIRKempYEjASl5wt9xTV6zrHbSWk9+JFnnGTwX
s6kTJwHhShY/newIziJpJQtg86gwJPWAVaAHkUZIPL9NQrujOXJZM1MyvXAp9UUi
r/2tcDLZTnV3vhy3+Av4oBoBmhVbptFtRawWPXgYj0EJ88qv54kHKAu/jN9pvIIH
MmI7uwXLgPZsTVyERgTKZpADkrsJGEQLGokyGiTpHnoeB0U0lhYK68OiHiLW8YFS
fmW7/0pdNawGrXaV8cxD7AxOBov3l5op6yaE0GiNb20r09Mzo/kkLfAksYbJ05PU
DvmOWpr8OQqwL4vQ7SWy1bP35erWamZqB+RGvpYE+REBLwGCZeAemg3ZhIerqUZB
5d2FPy1x/QT2L9h5l4KcV/rpwft84WhhiPcAzR/II9wCL1CDRMzqGDTu6eWgMWet
ChP9um61QCkk1XIBTymyCDWOOGEDzO23t2/ifpbdUV/VMHYfcPRL1ImO5ytPWTnP
q3v8zpIJHuW6Wm5zCG7ZuTumOQWwnUIYuEc4EBjV+jDE2fM7mXYG4SUlk0nEe2Fp
ryjZzbadpuIEiJ6aeI/pt/z1fY4ilfSJPqop9lQ89en4c7zM6S28QM11OOHOs+z0
X4HJNJ7CxZgcj5NxTfZb5Did3AvY0a2iSkIau0dGSScFP7x06ds9zvAvFOI+PKC0
wf/QQqfy0XBr6IC9Dom1qy0b//cSbl3iR2byoDhsVaqREp2tWopn+ulBn705mJrO
PuXGhlHhSjPJtT2t1AlqQ/80VH+e9AXMFs02tPVDMOT5SJuuXmWwP3RnxsERgS6P
MviWrjMA75I6Gp5YUgLhwwYO05acMo8mft6B4XqEr8BEDc2uh4vJ/RiOZyIgMMjA
qqhgV27KeyG6Z9Wz2iJgKK8gtVYy3bGLjHBGYJknjzZZr/AIuiNuE9KaqNL5MJO0
iQqOc+YiDtgYa+NWo4ijzOtJNfqMeep7tlhPf+2eHLnU/xNKye0pRhqgfNLrzefk
fQpPPWIeO6LDrkXzVOs/dfQ6PE3ez7+2nfSHGvJUg2yQEQfbQeTtpyRDqgy+rPof
07dBEy9Xal4Bo0qISquF4e1Xu+QAoMxAz+WTw59DK9YSfa4Pf/Mf0ko73E1ESQDb
lLS6GDsoyAkz+z4sd1zWiqtbGdSPgXFjDhuW0NZenVeM4WOKWvt9cMQSHeRgCYCI
4AK/bm0BuY2PN4ED01WzC5OB8/EPb7Km9fS7iddj8nNmW7PNSYHNYwC12O/wtGaj
HxSrXAox9yL+Q/P2NlbVUXs9gIQ4CQGIl4aCRjvb8h/RjtjPePAwstqPtoo5UZV1
GLdUARUyBNnyxSNyqdG11O3kunDCfG+ufy/wm2Rr+ohzOxMhmcNun4JxvJ1EyHgt
DW7tROxJKOiTC+ZW3xwC8X5qwBx2i8VBHWCkQMtetyAMYRHDJXBISlM224IIppPW
9rDUWMZw61dER29ZbazTFtj1+23UkEGPtIXyGnygRaMqcm9VoArfTeLJzVNJLxO7
ldmaHt/3Q5iHYtqlz7EO5AMf5fYrAXacOkXUnPjKV1BSWeigy1wSkE/z6nl9wxV1
pwiXv3tbhYfFF7MjPkhKDpphKhA5HgThkU/+I4uTo78TQeAcgoouyPGmluh+K6Bw
P4cJDTn7Mxj4PLBtjx274hgoNdz6nfsQtAPh6Io7cn972/GoVAh9cYYCvq9uM9jg
gdV+cQbeVRBf2kSmystklouV2wdrFqj7OZZi8zI+LBgd5eiS2x7CxArs4h/6LxjT
lQ0bhU9khpdc5SaFw2zyCDZ2iczvE3OUwdXAu5rgDG7tcZI8A20w6wmD2RVmfk28
dbT0fw5R4EYGJtDZpPVwbOQ6yciyWDqiDFEKvL8zraQUJqGIbdKFK4Biez4BVUWi
OI5gtVlFzO9ZgpeaG6PjFPULzwo6z116vtEsk/tcckiYKWM36+sxLyTc+kdOo+hY
kTJ4DGqnaKafZAosFFIxy6q7wAJi79SsvWDA4z4QlLl/GSCQoVabQDDPQGsDDSBa
XlqPV7hqo8929juUWZ4D1ss5LVONh7e5NoIdoX0HNo1doju/FF56JbmblId/LBQ4
RAbbPpZCIIvF24/glWotaHydVvi+kCOoibv4K+g6TWc2U61ssPalI+5oJMow5Ljm
+DlpJ81nWYtN78O7LxpoDQVei7l+aobtOwIu2UfFPnjwQaFeSfKOTc+kkvJYgCJY
g0YipPrNlv7LJL4SgO7Ox3fFm91MzI9pd9lQhvLSFImPlInV2imspI3CTHYSc45V
JCPHjgokioCQSxCjrQOprTZbadl4X0OeVTNwR0EU2jeoPJxwZk1pA6Knyj2xANib
KTf+9pQzfezyDLxoNTBrPeEx+nA89jrOnE77NFwbCE0cUlEQfCnreErsYVXNKy6l
I89vdfGE34seHTV2dTqQ/q8kRxgAXGXrM/HHnPCbI8KPz2+qNEWKk15Y8WRdKRdK
LYAWHcXkFx0p5vGERq79+1oqzuF7F+QYlHGrtToMdjP7cBtRChcjaAsEZFwnAB1Y
1E29ml3btnqAd4jJ84tTDHofhFdUs1+vZJmRsnGYpxut080HWIKshyfRih7Phq+s
DeTF+W5flNEaRiq2ojBVgCax0ZOqAIwSIYn8Ecq+4J1umthBlpO61QUw4S65eFeG
JtP9TAAFa5gkn4WRRidag/BtEmMVFVzzMPGC7djRToH3tSLnuX/zNtyhcAosnd3g
F4KRPpybDF7BeNYjml9E5ZetwujQOaKmnE6IPZU7VobLsbPbgjd4c5868Z50/dwK
9i6mJZ8jWzMMtV9MAnpFikrCOgMVoUY0ShWHQP3Inim4G4Y+7/ptcMS3l+xjf2oK
tK1jZGFaUYEdtZfSwFvAX6XwWYVdfgVDCP32bUM121Lc9f9FZnxh6qzQwPlEOi53
R7vqMP6m1HGOz1B205rehIFNhNKYxs7DU/aBKWnEg8YoW3WMxioumUhSaSS32GOA
pZJUsGrDqZKVZ4MCXAPGATWFbm6mbHnTeCYgGN6A0x8WnGLd6TSoJD/PVx3CwItF
Aq4HUjt27bC87AjkBI5w93QKHdZiir8eELiXA0m5DicXj3cYx7MSVvEwWSYLuU2X
uchq6jdx5rLdecAJ0WmVQrDzY5XbHElIr9wTY2RYJiYvig3BzEoMnwKJ1zrxd8c0
4o8AsqW0Xvywca9lE19RCli1qAx9FWxHujwJxfny1Zi5yuwCUjQNqZ4I7OEPtzvi
nW8ToE7DBlnHT17ZWI6iUPIiYlUnOFrXt7T0HoS/zSt12G6lXa650tLf+zOvof4R
D5rhdxNFVg+1CgwYiL6ScQiAnEe2lfJAljwcLhDNaO4ZzoSmwdF+ZtD8WkLDAbUg
ZMkLJlRL+n2nrSBx5fsQ3BXwD7J5JVLALwDG04sBZFs/JjfUwaTL8N1DZlJF1CdY
RyhoGSUDMKfpiu73ydF+XXN1RdPBauKkW1Hk077dB+9GKN3dZBGqP8x9u/WX/heg
C3K0yo5DUhFxO948rsaEMPsjRa1aOyO4ii/l5gTJwMquChpjduvdWg7uwBzjrdpm
5MRKanMf1QP2/+SIm3jvQT56SDBVWPX+al2phqroIsmbc4vmvXk0Oq+rufIPXT7A
Yq4KGgvyK6JtNq1qIxHIEPCa6X++iS+jCHCqQ2PQWXWNJ/T7KgNX+H0TxgGi/TmY
ilzZtCSyxfDElpdPm4JSQMrLZPlDYjiSmdeTlUaLUED1M4/U7OwN/KntWxV9z+Xd
s1G++/Invg2DJ5yk8x89wW4eH4SY0ar5LPdXVuK+xrOCGTxyxoT+M9eGdgURpusl
Fw8xcb4fK11RB6hyby012DgKmhUsSgP3LmAoGM85MuaZtQ5DTmo+CrpHbFVD8rNt
XviXe2jVAixEcrlCm0rnoUNevsEsW3oHP8UyQ1N91YNipSDKJMXhClDjdW8D8PJp
V2scw1gt56YPaFJJCKzoZsWoSj9azT2EbN638RVVbbyUsdhDi0gfRK+lG80B6Xtp
2UtZWQPMLipW/UymVSQtT2dKAf8OVEhhmqSAecyX9Vohzhv8zNXUqrkwUDLVR/45
gwqmYVVhKlXQ8145kBq+y8eS1Y8HE585djK/iGib47mtkdgJGgNg6mGDmju/7ZTS
ZTmp7blDjrXVgcNzgsee7zoskNWC3dqtbgzhDNhh++p0aNLY1K/NLzM2ch7hSk+/
KFASDW9l0d80j20PkXYnvrGsFEgO/HzUHx8+NwkLlgvaaVHeX135pnLTZ6Zca5Ol
fkAcGnfp4qa/tdx9h2qYh8rGU/TNsk7HFwhRGawwPHEhOQCotOT/AvR9zwju8afp
phzuiBoLrYpfo+wSsmU0G2chIGuOkRZOnL1vXXeBijUsa6G26wyG5gTiULQUOCzC
Rz+FfuzFhDR7N7nWc2vJTLGcBne3JmKxgS3hkJWfFqxbm8ZYeshgE3ZPYy/hZkMM
stYX6Qg3rEPvq826h5iYQRatHgiiaizACUxGjydrzGeOhYR9UOUeCL61nmi1lnKK
GE6FIvYTM8fp51NAbMp0v4YDA2WjYzVy3W5Nz5dnALNtAoNoIxN3dvecG/rTXX5G
U7HVs2FatLzqpFPkV2hv3YrJ5vcMDxoBPiiOnXEZNbD75gb2TKSt4Stp2b7kVcxV
f3bn05P5M7b86Ke+v5al6iLwNaL2DI9gVi1q46IDd45e5WzRRbLnRqUpWyd6j2WV
CY73V2V2zKAvj5PmkiGhECOfU9dCEqchwAjxEyf9f51Rl/GhXNHDvJ6ao0WEIXZ7
99SLk2HNBUuZCIWMX8aDbxMi8KB7hjyvQHUBPavUvty3+guJdht1Qx4vvgK6dXuV
o3IlthdDBFHq1XoGup3E2PHNbzHYF/SUgXc2ZFlVl2/Jx+dh9SbOijb7EQyZSQD3
Ju3N15uU82ATU9pPiMv3X249bY/BnY9LNDrmP6mjSmIiWIBCQt5gVeQIDdXG05vF
xGnqOoV8m7fHuEfPOYvlthfQVBZaZPzEBXD+dPq0XlXzaVe4+OOzagxG64W+6w4Y
3tzuHcLDomwcVJphjRowpES063YmiNgatwBirul60hVvcENrddqba2oABNa8OxKR
6j4mphDLlF3fqtq4qdn2r1yHhAXVE9hxfLJ9xqf1VWWe6uMmH/a2EFjDt7o6uvEq
NuDp6yuCQRAcyg6YEdpbDpbGAnA7cRan1WZFnkku86bteNUWSKQc0x3OZgAkkGhC
WKgJrBtgXRyeiy8s7cZl9vaVIFgNlc1b6id5A0/kam0itGuw0kIOhuf2FBffv8Gl
xuO5/cACrf9gOysZhwrsbePkuiYbXzmemLYcU5Th83EbJ9+JyDK7x4cD+bSi/D/v
2CtSc95B5rE9PayAxTdiHbjWoQ/g/NLfQkoZ+3ndslWE4qgVqosywmIgrCyn2rBk
OZiZ1lpA3HPKSBfEvZEBYXxKFACtDCuA4zFLOG0axZTiW2obEZhRruN2rvkZPsAb
C8NXbKw4BQjY9M8YbyDdBNiTBoy7kmSW7mUNbVngcm5cNdgA4fAESsV+skYgk3PF
OuuwF9eSRBFms08yDamFnyoyE6n0K9Z3yDmjydPtrukgqk/ydiw6A8XBBl1rvR+r
wDy6tLQWVShQ05YEN3nVojEmbHZgAaIPkbCMBxT+9K2Yo0nJNfjo4TxRT5OCGuB4
oSFZxrkybr0yHF3nl0WAKSjJ8EtHkw64/ze+c8T1aHlfNfxjqjjXWZDDiJf7drMz
H0GAlLu1RYx9tWVCUSYzhAs6Lh+WazR6okFPL8xs4cAbDCPB6afEjHrNKP8cUdm9
IFyKFQey8dqA4RuM8AaT7sIPoQD094OhufOuPgHP1ERCjy76GXHQmG4iOzK5aprP
PwZlakc1382b91uqMN40vpKLsNJxXcgkMOfmklMEaPklE2pk7N0ii1Nfhs+ueY0r
Fct+MzQAYIQyD5xJ9/CJLVhaZsSfaSjJdrLAfk/tuDQh/1xs+Q7p2CNkjHiQast/
OmOhvqx741etYatoSqEQJDeEfihnesmblqlnFvIE2bQENlhNpupIvd1YI49lnOCa
wAkM8K31+9Wry7DW6QfwlFdHIbfHKdwehCOmVaHbZabkey6xeRiT1VH2KVelr8j7
bGIl5B9kAoyc325cZjAEqwvyvSRP5SceJYY4clfyiFzEAywp9lmjakQO9vLg7fAK
JvCUZIzul47CfZ3crGtqOfSHqxIYuEwsD8Lfto4jivBJmwj/Ads43DMjh0o8sBr1
k9tfQVbl84Jy1rCknYFTIiulgjM30PhXWyN4LPUDNkcS77p/puNlsNI1OFYqNdhG
zE8yMVuzEUYPwif0wBT9EmT8K75BX6ZpvgSroHq44NKz1fh8nKGRx5gtIZlktyOw
erjrs43+KTJSVFPFS3htfmBJlcLJNMOY0601DYHEHafMaMcCFpdeJn0aksrkGPXH
UOF7RjSG544h29LKOWsxZm34D1BMJOCHtUUaZl8VND1FMKOU0l2wbQVg+sUCErW7
P+s5GVSu3OwlMPx69vHIAmlH8uN92tW1ablSp9xsxmIu4uB+OOlKc89XBcuJYCM/
3PbYG4NiwgnDRH9mZ1TF4X4qNmr7egEC0AKOZZe/fkFa5v+v80Hzso0JYTxTe8jy
htzK2cg5zoa1nUuAZEAZg8s85JqYq4d5SlWZ9w1x96U0XDd4gTAxRvB6Hqwhay8b
IRMdp4Qaoey4bQKewZGdaemt3OT8tP8sfK+PdaIzYvVYmt/qamkA0l8KazfJa0VH
2/K2arJudmA4E78tpchD8/AZ+2eGwkM6VV1fAEYhawsixuTuTYlTPHSNw4aydVZL
DO7x2GUybShFavUrOpA9wC7xoh3GRsw7C/lAD7cYV3zyrnhbJ6SsafhOOAHcHt6D
CcaBWE0KFfhluB7CG7Tq85sLqnDTMY3sm5u70MIPr85Bbi8yK2boiECmc80o88DU
sEfz8pkhT2J0JcRCEKQGtS/othfb5KLS15xAqzLw3J/Pgz/v/FrsZ9CIpzMXSWxT
8sVXj3wgBRf/D1q06QxWSopalz8VkrbFGycISDL13IuP43vvrtE2iujTvg2Jzm1b
DCI0Gw5OXlgXJJuF0t+y9sJ2jWgFeE4HKzIA7MpnDODQky7KPZVMIAE9Yb5KtPCW
cRHrYVXyR0m49QKqqzFoaji7Mzor8ALmto2363Ws+JmBcS0EcMOHZX5KteayXpI7
t5ixh75jUMnZj2wORTzw6CIWeT3NvgVW0o24VKTs6ZIBvGW9t8oWOyBsfEEz4Tkl
wxZZQOtl5rFr8F7aZHswu45lkd1C9JQcIJqQ5iQsGGseJjKngWgdFy/W5iT8oCWM
xVxZhcG/JbvvJ52TpkiKWMmAiGXWjXrKjae63f/6WKt7Sw9JHzrzjgBe1vE9rw7E
/cX2o5Iy/v8VaVI25i0jEO0Guv1B9pZ1dG+Y2KMh1/XxEvDrqh3c94lylKHGrHRG
+RKdxMRV1pN+Ty8hMscbkyFSS1OYKAxL3nSOjsD1G9fJmR1HDLhjVMHT7hASxERO
BIB5yUvyPQA2mEMDyUYuNLfTAvc5Nj5rRtHQPNOGSMgBzWGWupZzT/EvoTsp/5EY
6m5X/uN+6DK19eYCDpD7WkaOvdzIhOeCFHIoW9wbjoGlKdVskI4df+O3fUiRy+6m
aflUoB/QTxjDIgTNPCtb/1rSg3FUb/wB+FQyuoln1Ze4ZZMCCb7XWsUKyTp541F4
lUK/NsTVP+kXHWbA2vvmhpvYX/IJMf0IwSsAV0K7Px58le5S5/zC6FmVn6+5UPD5
0ZfGO645D9LuhV3R+IGqHkWh0WenEEVpWneQFsYNY5hF8z4rC1qT/6klphSZBUQH
brPo77Q/F5IFN8FKpoWWAu9BIoAO7w+Ivgg3U2fsiEFIGYeugOtc7AdPxTvx6vEo
LrPPaWyh9nNV2ZsqhPu/t77ySoH+COS0p2TyxPMa2kEBxN9M0tZOi5d3MYTQXRYb
47Zq3fmW87D+4q1gNtNwRE6s6Pf2ZYPRf3UpXgROVCIRNLZQH2MH9EIu80NMTAfG
bP4LEqb3q4j6gqkI+ptUuqxlwh3nO1MhxQfuUCKv4v2n8RvzvRF/z5PFYZboFMiP
Y4/a7mUs8gi2pSZCBZwB6yb0gZ/MHBO24dq8XHrFEzcyTKZpDaHwMjtkTLtkt2aq
yxA8gbaLRIUU/EbURTF/6ea5bhWbPY4RH7B1zWp8uPbsCvJiRaM32MD6UN8HPtFw
j2DfkDO4LFeoZaZpkKpeNx3HQ8eIz4ZzmEfb0cXaIq2INt4hbY1tXqoFJNSlhF5U
6Uw1TQGuCNsHxKTw94iCV4vFr5fT+rK4Erweinn4JcCEXiAWzbU0E3TjsQX49pOa
HIESWiik+3zLkjvL4OUAKDcptr9oucy6hfZIjse14XRHAZtAWOkXUrFm7F5UbP1O
QJYODgP34eUYa70sKRfYmRHVUvpMuF357WbwCcjJIRt8DO/RSWD5r5nWTSOXa4vt
Rb/DxrY0LDPDF8kiG0OHugz4FCpKutJOyylKm9yzxDkHjhz7DqHU6HheWxMo25m+
b0V0C52iCsXmbKMi8AMu5+dEYWeN8eZR31OzuYYMFwmMeQgQaJFtP+nOx3z37Na3
0opeTxmUUjj26WLqZmpan7K9dVWTDbrELDWYfCd1Mm4LVWdShU+4yZ42z5L4r77e
1V0oBF8uqcgEBwRsWJxG40nVevXot2wtVLD8FAKFRcx8zwhzuGVUnmvWnGdxjgaO
bsjO1ADZ21JXOCObvIdhsTY851DeOdG47ww1yIIxIX8OOzdM9AeEJGVR/bdjGinZ
12ITbXLmBRhdxi44lnnlp4ItYIwAke2fHOaVsDRzz566kCDH/v5jNWzYBNeQmtzk
FCGz3lHKgtyw0GrTIxZiZoInlbEN6ZaCDw9agg1iFVYyBw2A4q51dFG52FLvp4FU
LWYobBnA1InDtqWYOBRBxo5uiQ00Ej31jMlIpmQWCqQyVfgvA5e4KUf0054FtnGN
HldFmmUVFPp9/95jf1LuKGIodPkpZGNV36Ly4LooYzyfZXvIcx01M2R+Wu/xKGcz
EdzGRiDRweTbpBGh3ozGu6tgdoqfCe0MbAI1NKb+/dAyEmUL1u096VIfseN5nsT5
AmUBcVuJySEVkm1mJvWdm7sZTBiDOECGeKEj5OEodDCfF5/9CCLoB4fK3pgl0U05
lHRvwDdbokqhaF5XMzeIAE9DTEWFPRWuG2NBKTKLcceVqbV+Xup7RqgVlEUmMcW/
NrDpeOA4JDqesPW2dJl8yzEYgz1dZSdEu3h4U6NPfETl1qk3le7ly9QigNt8tAgC
3DfNW/o634050HUAK7QMPVduQ5JTCmmAdrvcoZ5tMa3K9tY5hdzuWUWx/GAbel9Y
wBpEtXuPM4NQJmgXIvlyXnJhh91BxBgPf3ARyNiMuef6fsKQZSS3OmHGSvVJvlq0
VoeLdqsRrXZYQSDSOvkRbb7lOM6srTO1A/prfRXC9KGmjiAZvZZO3/LKpugPZu1F
9PV1cutk8Qh0MbL0R+X7pW7aSYpRG/4MZKBh/uIHQEutZ7RoQ/gxRXUhOes0VeZ8
jOhmf4TcPfwZB00J5K7PbfDJj6nKgdcEP+mHAB6fMbjtewhaqx2AGx7fE344Kx2d
MHbCj6JVDL+2k3fNSzzpOF5lP0nku4whobfojND5PwkMIcYs0pwXNGmsBAZ7SwLW
0yqC/w1T0U3SmgjQ5/f0rLfJjH+a5mbJvrqw82lzq37Px6XnNNg8co8immytNXP7
Yr01LJuZ0VvGOHG4O0b+a1IjKC/2EyQfN0owyso7EOSx4ScI+cTTWDqUWnI6QSOW
M3o2+PeQdOm7HfETOJu5kurLnm/s6nRtbQZJGaJYaMcwlGNoOv1L63p8yQoR3E80
P469EJJqrQAmanozIa4GtckNFqQ1pdZDUhv5UFZ4xyI/D5xGKmaECCzmMsZs9pzx
Yn9S78MwVHFskXyJYPVq0d/LJOznDrN0lozRBCw7MWnCgLU3XfBacqyto+Y/M8aF
G5ehvpS/iY4x/QiDOSQSkXAoC4wNWfr2nAHEgVr435aIBSuRZwwFXGyd0+rIEQy0
JTnBKp1c1UMiYKNxgHUBsQPW0HbId/i70NGwN7TUjzg8mgLkdpLBzfSXAl8wdHg/
JmvrGKiNOSejx8CuNFV4gdD7p/NvPuoR+wCL7dwt1KHnyf/Ny1gOLfb6IfOOqub1
FaXmW/UomNTmWJ08UgqhwLkLHbIgObhcGiOrRiyDOEpL8SpQq4fhK5yRHfaVyTwQ
t0QiS77nDmyxZEMfwTpydXrdbAz4I2EJO5fOe5VNaz2LLWL+t2vcIGiAEYEZdHvu
hG62UB+B32XUxoI0zoNbBsHUWLWfGZ+uFSm2qrwyS3KmbhWlUw95Bs0l2zD/X1bd
mmrB63wzowC3mtHvxj3YSMHFWRxZ4qwX3JJf9XvYUs4g04TwetFMAtUDQD3HDjFE
Luv0aPkgTuTvINLEubgpyotkIkpC8WDgQXGHOTURjAbaBoKfCA4Qmxe8FLBl/Srd
IvLXVW31L+mKDAyY5JXrbZb3a4UxF2pHZ+L7Iw++gGFQ8YV/CoGN5KuJvn712g3x
A8/lu1N9RmacAkSr/wMoe1v73DvYvCgOxYSH68MCEqhR/sy6+OzSBHeeDXjdl3J/
BdQJ3l8702BbbFkdMrmiSmXMOrS88v9jtnycIc71HBOL3iKnybOrhr7GLe8zt8AT
0jPP7ohveu0JSIMct+LcmCxX/dFdNqwhGRhqz/oqyK8SokJbGECGyOzQSGUeul0U
nAG0SwJ2FOXjA57Wkh9kR9U+DjXmp/4exCqT5hJqM2qr4eAJQrPGe8zkp+1zlo5d
QlMPyF1PTeTVHlPLnEGQ3WlmGS5xT4AWjX8wdcBNTA8+ybs9gENgAvSu0xK6f3yj
RY4PS57h/ywGeQdTpjVNm4lg5nxOWncJKKPBchDeR9vwe5GUiYeI5/XofNvHAQLI
JaNlOlTMxyyuBJgEIj6kM2wKikLzFPygzvS+FlpvFlW0iMml0+FltEJz2nOj5rTs
dA347csHMaP2kOUE8geYNdAN5/XoKyiU3bPJ2dE+zB9iAwuAUxrp8eX3vNwAwz1e
5JlrCfpw89Ynj8rEe2Ftr3WvslhkdR+Gy8khweZH5zlBuQAVB30SUshIcbju7UpO
k6tW3o6hs9FUHXZZGEkd3HUPqSF2M4qVgyEo2z6gOaJu/TcfsmYe7TcwzTlLA7tm
L37tMz2MlqlCcmMMrJNFmK3Ix05ufF6FFPSPphWJtI7GKpetjfKBuvF3fViXGkTM
jL4HxLiAj96Dnqedf5Wi46Qa/HZ3RR7t+phyLwIt1VCO5ffeAxo55UDrgPo7jeCx
YvZM3fCBvwqM41C/GbRjWuoTkGKrMDltmgfDHgaid29joPB11hhnt1owWNanqaUK
VuFs/O9MEzaRU60C844lMoaip08RqGDNBbHweuUy0TJy3B2QmVpY7aEulvuEsl7M
MB7oC4Qus7s1+maemVJj4tlGz3hoP1PtK2hvpIC95cekeiN0f8vgQx3+cUBRWzSQ
XiCrqmwF4e+SJdOKVf4Q7BZ7M6FJ9fa1/UXdTpShMZCE6Prx4U0XB03BIFRHd9bi
lXKiwjq5gkLXnGG/yo8iKWU/m5HG+tYxrKi5JR9oMbnZle3w1onGfiWZ+NcUgkIr
YnYkT2KcbpNvvZdzjtWb9LIh51qQcGNOtosxjdvQmLsW/W8APGQZQ3/1qWGDjJ6k
n45EAnk7dW/Hm6rPKoa8+pOr+zjGUSJPIreCDPER8vy/aglAJ02Skt5Lwi9vdSoI
9aNB36L1xNf4yP+eI/P7/zrZs4s2kVFtrhPtHVH1bJinqdL7lkt5De3uwwCR5Z5y
i0AFuGuQaMBwhrUcAdDwdsx68GOuYz/aMw4E/Dn21pDzZaOBjtUbWm8h6nrQPwJl
OvX6KqK1LGly9GsP9Ynr+Iy4RjfuBrg8aUycDXBH3vNOyDYLTOkUWq2xrjAwFzK4
VBkaDwr1thjZszDJ+t/GXDpBuKyYjaXRMXsoxX638CDCgHxWGSrGQ8htmq3dR+jZ
9Cr/XDHUL5SrUroF4724NpWTbVERNiW1zWpyg4EMH7tQF4kxNV9Mw/DKE1HAWjTR
AV13CE/oDr2vhgcylvnUacsAIAQzS+v84Qn06DV8UfPbiECWxlQjk2chmdaNV6t2
CtpjY/KRiCXnyfznIf5JjqIUdMIzovTXSjyc7XS3YZSX4qB/HLBbU3kddFghsTqR
Hb40KXYW9LNTOw1WHCXbztX3m1vrXBfcfNpoLqdKmk/rWuLmwAIeOxn6XgCwv8CC
Foy8lW8d527aFJ3eNBstoGzboNiVGRrJrv0T1DIvL1IMUHVPnr0Q/u7CN51A7kl/
MJbCD6OvH/mq1/Mo+mrNQXrWFev9PSUJSkfvC+nXylVzMUQEu3gVzVpqaHfi3hMu
h4YL2EANZkK9ASrVd6J8I/tEUlesQNr6H/yz6oC8R5DYwQaQlzLWZrSsSpwhDUzh
/dZofvPGDkiFBVv2Ewy3qWdkVKYdOH95krP/p1VS84HTQ8GscaaGKLUX3ydyAHN8
R/pXX1Y1xNensqcDB+VY1JLCdXb46hqg8ZwPbFMBNwV7ylipnSm/9daPLu5OrOKM
G5XH2LnPmdge5JsZmfkZ2+xdeWjNYZPfMv6/I0qg/NJ8Uxen/hQDPfvlVxQd9FTD
IuJSb0MLoeByGg4ZtjEuw5xSthUJlgf0BQf6mCTgASBKhDWqZByUbiZLEpWroYTv
QtP5sKIsz6Ol0C3GVfJcXJ/pSfNtOZsQBo36eEJVFCgV+rriy6azF/GnoZQlV0IZ
Pmt4P7kM39eky72GbXg1BQgbNKNjO5PY84fBDdrnAaBoA5d7XhOwk5mFacxHgcoO
EeO2milc5UXGOGJk3J0mIsyQYTOwNGkD1tADI5QpaVCZpd7lj11WikOUgjPP4dPU
y5bIP3RpoI+bPp3Pw/NS4LOL2Ub+FvKIilnWp6IreQnNHPwQYUNNKUrJBcdf6BMo
1v2TGqeN94/w//tdgySwO7jacG1QXz+hZ+8OH7LDcbMMWQyvAK94eAAmHv5rApZC
eJ4GHB8XDLLPEhFoxBgjxgVYYJboht7oIz9ro9FNSkt9hIEETLtpxHPCH6pHYGL/
jSQaaIUxuowlqOIGaYkM4gCKjCRySOeA8yvT2dgyN5oXW+Kkn3Ar/v4wAXg/6CWF
I39rKqjUVS57xcfD6BgAEc4pOfFOHzBzSfbtoGh22JBA86F9IgDcGnF7czP64pxJ
YR6YVAMsXGWTJXChiTyrPsKS3dLnZ5FF7hn3jB1TxM7PLL4M5y3TWzBMxtf1YXfJ
fEXvPhk8rzOijAtdmWslXrqeBg3h1DeQ0POuLSni3azHg+RE5JgXt5HtOTLaduAu
/+fXf/lpjwu6PyDVp5eReLDVqSZwpDQ5Y0g2mcgOWjmzU85o0oaGbNEP4DEyMMZt
WCRThpWo98MI3aPaSnVZvgN35QjtrKZd4Q0/IuVgGTIJec+KPcEHQVggH2eW+DKT
/FYYUJvCkpzn0NP13V1iVVCvPcKu3t31iQDv+T9NN28uI/LKt1jt9Mn1VUbIzdpX
qegE2DCjqiE3B0AasUkx5gZk0vql4s8Rq3X8Dgg5/7tlVgLRBeY2q2FDzZFClwDN
uc+2SXYDBMlS3x8ldLI9jWtmurRbEnsM1dp39a79A8DjaqcLMD4fpWrNCDSPM+xG
Y252ukr9Jn70GQ5ghpec5JksjHKmA37irVPhHU0/oM4fQTByBY8u7c7N8MpD/hhj
4EB2QK6Z4C/JxxYQ4ALeOl1bQSCHDkRy0q+zydf0bPT3gf1F96/qiD0PTfaPW+nD
zCrv8OYJeoTo3uxbptcvqR0OMo7vx2McWh5mX2zjuCBxRZ4LqMbXe+RZs3rbv9pE
K6M7otGEVhku2qZr4nXdWRIHDUnJc6EcvQP9kuQlCltcP9mA+aoNmnjkiqfi4ysQ
Vdw9g09SZ9lvrsHgwEFhQ0nR2cNbVSMXzhaHcrI8msHYAFB34AWU3dIXHbVjcPkX
XffRu9919ZtsBAmrjivG3zVVIdtgfJ5cYsmztz6x0OCeIbVRbd+eQyb6hB0Zra+S
dg5pYdthR1GSLqb65SRA0EcjSJjrXnSAqqqjGNdV7Vkb0ze77Otx4tmm+1r6YOUR
BnYbTdByZmUe/7DTOkTJ4+k28J4kwNct/ZCgjxbeIaS1dzQmxHljWCDNnMATUzpS
9mDH6B39f4jDYEvcSamsAcv9GsxaxMHvQATkRUJK67Mg4RO8NGJVMNrJho8Ae8ww
xXBn9DOVkd7gL4Rmfmnz6oUoZaOBOotE/G02rxMEtfKxC46JxKWrruI7THRHtOg1
IEkVCrLHsfDch94jcrdp89Ez+Yb4hv0XWSIGVsoeRsGQRNp+4GYCFNYOvIneKlYF
GMcmP8aU/DtWEY0FmHLQEaP0uhOMQ50CxWybN4U3LNV1UaIg/EVSTv7rp4uxxrUW
DQ2hCIVW/v1WosdE2P//1XdwEVsK86imUr9Rd9FKsbtNM+/LVs/un3dtpOUUYQ71
yScOWikmRICptCE4zM8N9TdyNRLQiQ7uMh5Yv8zcPWtNHpGYJep0OyTusZRgfokJ
wfvchKsKRJfr6xnfMJ0m5u4V9l5Hb1RlCjAjrRQyFK7TP2b71lv6aGw2eSy+fr23
NXqRYkVdZF4K9H71OqNFTWDq8snMH8T1QxAyMOhb/icMRBauT2iM8Ao0jScJ+EUD
S/D1sGUKB10ZSHp1WCVR1xu2GnU5avH84okhx5C39aL7wyv+LDjx2EVIimLCe5yV
/REXaRJ7qOFKoPHXqhJXnsicHotQBUSsIjyn6ZlOAV9WCN/QSFs1cH5P13ENiRt8
HJ2JoAq+Z0r9rQ15AChDCooRqU1kPx+MlMDeCwmHyc0I0khmR0qxsVcLF23rbjuD
4aB4W/FkBZIyeqyVV2zeRrv6CDmgGzAwcG0PW29pvHxhZWtrcYWo8q/ZwOw2nWqY
pEL0JRvJrQ4EcDP+n8rCgBO2f17PVfpwaS+958uApn7CISHpbjYWVPm/vAuNz3jd
SmAVd8amSAhBA4fzR4SCywIvIxyRfYDLS7gCiE9b/QKby9GGEIe9N+vawMYsQRbn
8aSPFDJPe1QcymxrN79gkVE6xhWV5R9d2CDROqZ27RTTvMOvogJqtXsb3OFFhu6F
zMq1DGaA8q9KaJE1hd9Lcea1vSczLTsVfaLRuaR0+WiJNvV0GGpSzcnkEs/6uZEH
dBb32gPgJfvApnXx3t36awKJTU3mswaVETRbY9DAgQInrmVYGsHr5+DVYCc8vmaq
iL3NmgCDijIYpxc3iZNZ3fMdelaWInlqzXfTybFdmUlCloUFXQsAY/0rJkxQG0w/
UGE7YF54YsV/f0qIzPiu6IZvrU2oge9Y8tFn6xa2ScU4jW33Ft+4/Mv3oh072/H6
VIn7YAv5UDkepYgQoiYH7F0SnVj6myfIbpVF1D9VsPLXvHIGZWFZZ268nBAWaRfP
1wG08atpv+B6Whk0FIsRmYoFTxQ/VEQEdCDr2Mq8Vd7zA56EWTTwqHZDYeBEOaKb
TQa2D9cqSr57v0WrtuSkhH+35W31jcjP+rrKPQghd9h/7muPAe133YNx+CwLmXdc
6sSNTyWxs6pYf+EIhDrej8kWJldpgPIKzF7ahQ4cr1/0RwjJVUUC7pW8JY+pcIvE
1DVs7pdtgAJGd1dkjW2NIfRwMza/ZOjozILAXZJzBgLfPUuiU+mg6WjUf+gZEb2U
BEZowIMhdGHjWKQDlCSLlJJ6zHpxOJda/YAnuuwVilBoBgUSxcO+ObALQjFGq9eN
fcM4/jVQAKkC7l8kjeB6/r2AqgWeo41akHCRfkkVORYClTaSjQ8yyBMpttuTOJDc
8HqD/1ITdT/Rd6R3ZI4GoURkW+4F0ZNU/92Bj+rRbQKdTMd10C73ZkCiAwIujXhb
5UCXcEDAfDbXSSWlg6BlDdhzrpMuo15pa8OKbccArKs/L5z8TfFDL7LGL9ckhUx/
MjUWKY+e7E1m9qmv9K6H0JFIAvX2gIASuPSIGsLAG3tlg22+9Qshmg0PVofCOX49
paYZBtGlZoKiVDpxlfGDTwEo9j4xmA75obr+C2tpbKcdxTiPV6fXqL5Al52b3Tlm
uT1ozyP4yMWvtOrgwryuaTFu0Ak3RRKXtxhMZdTnNsTNSXS9Igd+vcjrVEtxabxC
nHeXAbpTTpbab6Y0ROOtKM1/ni3aglKsym7Ys8Ss1P9zAV/Zfq3e1G42t1dWtBaV
9xqPWq7bUiGe5+LAnh0ODE42E9Id5d4Zdz1IusW/nGlDYSfFZyxdhj9+z0Vg9hWE
+QJvZtaaHUas5Z+C3O0mC88OIh185XorYXqED83hAC7+GvMCyf0Q7q3+mRnb5U+b
CerOnEKWThnobdKgemWHQNyWGdCdwCZmdkqMJPvgB9vbsMZd+awmM7EW3J/jAt+J
j+Srj/wd2Mw8Ku/Fu3ayYEUCdjbfkG8ZmYJ0i3XfW5B75oH5usZJuImjBUgZ0WJ5
2yAKaMMnpfhrJEiyHbnfVkFRS+VosCLXTTAHHwv44eXU2RbDJKTzYY4sD5FXmGjL
`protect end_protected