`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTMxKdsgGXJg7FTY8fitmuVSWO3GiSp4yzqeEu3xDpDfU
Hg2NTTZIua0+CQIAVJrJuFmzUc01RA2Zyyno0q5N6TL8XG/wXjzn+xnHPIvlVkFX
1AqVU3n1a1kARkKsPWs5zpKy2yb5Xndadkg3ZT3lPMQbQf+ZAaBy/LvbY8WTNduI
Y5HL0tNe/yovLgIK6yZLoc8V9ZYqgxhJLCcaEeVys+aZGMTYTa8Vc2EpgvWMT0Ae
EIsYRVZ+8hpLhdp/iOlPClN15Jb7llYPT1ILutwuVEu/gjSpKe4+YRGA+5m7AinW
Sk0Pti4AtgDtKaiANmNLcX5xsyhX9ONICSsj3bptHfSShY7ygvdHXO6Whc4603Om
/rJ+bTLMnD/VGFECXa4Tiu/bzdTT6UxRWoMFB3ndsipvWH/r4SxTfBj/G4Gm+H0q
S7YTWwxGrKKHZIW4CNPLY/qfy0dzBkYk1cgXZ+VqSbdUCfbhNgASlGa5yBHufOSR
CSg+NcVf1Stj7a4yt9tiUDzg+9T0u+2mLhMOncGt+vuVij0jCFSapSU2QiJ1J49V
X8PmDMzH7QthYS9899JZl2ir2nklqHd5FpNZAryllTcoh/A//JWF5972YkIm3ZIK
CZCjeQG0FaC2rr8vyhG/SNN3Hn0mTzLQCsPICQUvlBGKfqDrc+hITjBngz4wd4eT
qMgRTBe7BpiDnU9nLGcz5cltVf/KApkFf3gDGVdnXjKvA/rkwo52CId7vqCMfGlY
tJVxayR3OfJZL0M329LIryPOAQUAxPAFONUYgASiGHL1DpOTkYX2FlgDP+z/ShvT
i6AFgstINwCIoyMRFyiBegmP9k4LwcGBoyEjOWHAUrEjHQhqUoEU/PvxP96F1VM7
cPoBSOdrFax7HWP/v+rdcS/gRGpCsjcDCDEMozAEoWrMm/NihuQ8XI7r6F8H/gLq
zcJ9N8DdvzJACA0WFg4dZGmlvDTHIrfwoXQSK6Txhp0YrDtf2uXNEkycJfhq1OZz
WkYXCk/Fp8T7fAw0WGiiNz5d7B72yrTE8S1IjX5hEIblE88nvCnq8eAJiNvn7KgW
UgK6Tng9FZZiBTKSDDrdV0ggV1VRLJ8G5guq5pf6iH9BOiaHL4IzFysc025HQqcb
Hwt2gCJFLhdEHu1rg2T+jpnb8F3mduEk1Zqqe3Sqj48p3rL8d26evTLN5798jIbn
hpaM0ACAmgW1YZ2m2ACQXJTQXk2C4pUyLv/QQKSwwpHYnH1YidyCmmJuYWK2GIhN
8bpm/2AdeEHPvT22g3ptbmqMLVSOKb43++RHlZuCJmSHooTyWl+eSENFF2WV+Pmf
hiElF9b6pBaVY/2ZHMpBi3WxdilFZ1zxPUoNXnVUudyg9MW/U2M2Jay4Ii8X+PK9
LBEyjHZl6/XzwnCV2FKWBneLQgGbcUA/LNYTaDiuBg+hYtPNMZgAcrhVfQyHpLOY
rk8aD+x0r4MsBROVyvLjpK1hDDzgK5W+iDZfMPFgZgVCzvR3Vcu/cxpQWYzLL1hb
PWZOXlfQ6Dk8xrv69S493wgbOl/n4OgLMEGo4v/QHuSRl6BmVikbaWUH8rmTyxWc
C5kkXpKp9mGwmoStvhnm+N2NbweCPSTClXI9YrbyeCi7KuQQZijXXu4fzl5EMsL3
9LFVuHiRVtdw2LJrtqn6kgc+8S0aKZXeasu0A+Np245o4Dws2iIaQcUceCaNdORG
q8AUGZ5zQnDrOtNrBcoq/pjkSIFFe4cRC2aDS320Mt8F8qF5CKK2LYFlsfKg9RAB
W6oYscEeUSEbRaDD6VLg7poyHX6OVMA5viKWt2POTjPFumcTnlXlEEPbwCxYcY9k
k08+dE5a7SAVjfSazXqW3EU8IAWPXaecj73CaWtoRVHxOdsukfmeb9uuWpsMuHV9
lcnw5lACgQ7cAbaf7OlkMRmcVBYoYyK7AXsfjTKwQMYLehSZc4b+k1FOeKHq/ryF
a1luFHsNbncy4wkKqx0q7USUUCqubuGypUMdUUdJjTkkZT2sBqkmtdQf80X2UO9e
kfgTWRkWFcMD2WqQBiDpOWoP0b1qLjT7jpPp1u38nkBVjZfHtdsvcAIOjRQAwwCR
n8CCbbjyXQO1Nc3Fw3XMwRBUFqVwV3eQEsW4k8nhHq9yTEY95GlA07vIHU9JiQkU
Vv4rpdxb9Yxsqjs9R2dV1DCxXHDMNfXJ4q+kC/Yy6Likj420FQvsXA2qhwyUQcAL
yJhpG7viue77bIAMxPwYHIzHVoUdKBGMDtwUc+TbD9617THUWoNU/mSn5m9QhzfE
T70QRkmwqBQmmrAbfADDBzVDqspfT2UXj1UOoyF2d1caueMl6l9V2+eVPKwJMiu4
ZlzOFh0HU4nf9Yy8p29W/y0vn7MPgk2Mmkydz1RT7/7NYBPYIELixdWJd9sGrjIO
zK0wwc1Z8FKah2FBQbnk/4NIGp5V2G0rZ32KhiwuBEsbLKl7+MppQYQhX+8DFMSQ
zoke0EqzRmFvthz4PRGOSj9B+/59XyNeOloWdVnmaFHQwf1O3biMZY4WrkRs4zW9
ZhDIdeTiiom+i5teCxuZxEZV9flHE8Bdmlpyd/9Ah9KdTpqoJE3QHZzkH3cp4yGH
QfiC5uusns50xz2D+SFSZFYuMLqqflDvk+Z2+Vjt3J3kpjpOQaQ+3N0fehpxeKpC
KRLC2QSIJ8SZEvHagZ7dkW4yaRRzYslY4K2WZHXQJ/8hq1sbYFJzA+y7bZ69kY/k
zOFQEM9S8XujBvi/IGiznqLQ1PvVOp8Qq7A1ndzo8GJ9dtJhPWTNXMZz45wG3l/f
c+8wm/kU2Vk4tMd2FIG7xvqGhhEa/X2T0DUMM8zd+omEW3Yv+ZHpkjxApMiC81zp
rruPrtyvFhT3fVffpmaUyrE0/ORI47Vn3cfZupl1aDx/kK4NAZQo7yp3bl8dpGBx
U02f5OyfoB+ZEgVZaUF+ddhTywbKCuZVnMTgHqObKBr1kwSG/S0duxaimNlI1rtb
OTdb71b1sii+kGT9CmiYNteJft2zNNe0m+1A0i7IGQQkYnH8RQFa5HkMZo/y+nul
qPzfP0WskqIrf7iNnEiBzJMKWMhUVpL2i1FvnfJ8aY4JVPmoKhoN6WnklZvnNRan
L2iN1qr5EkCECHXhg9NpDWPIxQcv98hB+EUAd/SP4m2cpeGs+HXassT1sw13E90m
nEuGa8pYiY3YM/8AbH30HGgf74aM9nP/8TZQXIceMPlqnBS0Cn4l2DHgJEPwRvzG
tWKk3yRix7wX1meeA8YOuk7EAtucZfsPorIwh79bPQtdhEUcFyhvexrgxERN4fgU
+O3x0nnnlKd09/nzRF7eohUmYLdJjsra4bzkyBTeMEuy9cBv5PMW6a395oZ95kWV
XJsrobz9QBEY8+SSP4Dpq4KB7d+mgRjj4ev2O2yXhC2v+d2fIfHTUj8sZ4VDBKSy
PkHZhaxKyYBHIH+i0o3F81sRxla1RODoFxcxrLfnpdEG45ov9TCjbEEggdS9EF5b
WI38Re/6b6aKBatZppjlDrR98hp29zFWqN2x37T7HRqId9nxZIRAP+oREy4xb6T0
/c0DZi+A4256ZKPDzecLO7QpViOQUNdS4RX0Pnc5vHdmeJeB4SkoZvKCn4QpkFWV
bpPVq9hjqBatdfuv2Dpup6mT1XkD+S4M0rbMGX0J1t9teiZtfgt1nr2FajksOkUX
MUPgf5E7MvxkMVT2kpVcJhvvvTcuXMcBap5U87/4vyMwrRcsOGWpqfzhU0SGub9o
P2wcJH1KP75oV/SC4lkKeGQGBJbp+3yD93euCyoOZpbeXEnptlxE1z4ZcEssj2qc
8kd8KuLHWmrJYyEob/NoqfyNwAm3GAK3bFEH/gJTSbzRYW/PbcC/47FUrhCb6410
32KPPM7RRZKT9PTf8jslvtFyVG/yVZMUGnB/V1BmJqatwyNtlcupaD5LMME+5icN
kcrfdlQf9BLD8KvsFCh3VOy6MKtLV3SQ482HH2sedMjhfgQEk/u8L5/JzPDpCcRw
eZuqZPuB7P/KbswRoJ8ab+ECMBQivwYbjggmkqO7xpav6lUxiswrHDdKTv9epkvH
uc4vL/rZKETJrsUTsVEXam1seYXwmZfPMsGMlGHUF0vUATJilp06ApQ+MKl2iLri
0P+SF2Ybqc6Mh8WvO7FilFOdiNyfNovl9K9wTcD6z4+DlQSCVdOlb5i2NvCfjz7L
GR/aW7f2xntZ+7gNsPaSN8i8I7qNhC7RhnDWF/sivmXoOdpal4ydH1yaHNSv8IAt
eV2vmtAOOFGWIBsaZdCpED40TdQMdPLoTn6keBSdJVD9lDkwjfJtz1p/3eMKF49q
OSo/4WszZC7ujTGRZ3yUdigbi7Z4x/65Tlh5DPM8ISMFQEE2Wca6AXYWcjS3J/oy
NCiZNqrRPf+/6CLsWcXlSWfxJ4DryUPVN6UffKrcujKX6E6jbPILROu8Rrr4TglU
BZlFgegBC7osI1x/cJd/wi7B7LHNcg2yap4gCtEeqq7U7GNdX0Tf38jRTIiRWjg2
3wT/uQovgfYEX3L8ynKmFLugBqy3O/Inq52UZyNwj00DyzHYhCvFkrUVryQay6Hi
WYO4cqH2GQew1ZtXktaVM5YGuZQZF9F6qr6SRMroNKTegb5VPh2spqhXq0FWZoke
P65sjzLEQnNkGWxPKNZs/s2cmXpwjaQjnN8AJ1Jk+/tsWjhfhbzjhVD/5FPoLaXq
Zsw8gp1JKzm3xbgxWODlRTdp/hJluGmRxKSlg8BD+T3ECNOQOdJCFXw8C0GYmJJn
qNcpKMWM0QJ+5YRczc8/T5ur81odaoFAEx6qNwAdZAlnuzymqvVwPjJGzwjmJCAs
4+tlqcwiMryvVLzX+DBvN9Zof5curzYsQ/u1NWpiCuh8BCUnCi4KMAxBLqWWlxWt
IYPFL5wGr41LRkPFHP2Zyjy6hUoD5KEB8sQ2pRr96ic=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8uRJl2tNK3AzJpi773oe4yU82FSDywpRmPZyDjSf1E3N
UEU3+m88BDdr0PQOz6TRSs12bz9YJq/npyApn21stM8W1Nr5bfHDX4sO/yu4G0Cv
6KG6ooluSFhbf2LCBUE1v0DSIYiGxg2wBzkRgn/uuJ/CrCBr7qLkxDrV4l+SULIH
/78S7z93j1PiFfXCF+tPKE8XiKQTcCN2wq5gFItn/0yUvbsBymvHYoRN/6e+9iqa
3JjcIBin52CkOoGWnbEtir2thDh+aUfPsSo8mo0HiZJyQ7newCWeRJ7xEk04R3Pi
ed4qeE1rN/pIeUZhl+6COzaWLZx7nQiAt7EhJv1bp7e6Brm1TIWb3AYq7CXSzLNF
kt6l458i7HEnbb5MaMZ0ZRdLoAxKE3vQW5soPS6rqHmFYqZ76HT1jJiQw7tvyNbv
7U432gLIsOLbMOv/I+C/tHTx/IHErY4JkkKWBStVQhMR7sVVQW4FJhHgoLdZsPuJ
EZPg4VTo6CIKMVmbyLJIt9+i8uhB/+G+B7Zh6tMxJd5IFkjKM2dSRa23GZMHwDfN
Pzpq/RwlM8oV/ETMsqOxFwRBmcXPbHSJXaPFddRrPe1lpEr0Sn1o1skIwxuERjgj
ZVMcrTKK237J8f3Yw5cbfLBGfzLiB3zNsgyBEO4PvwD5JROjja0ynmphv1KrDcyh
QZ2OCUHIvq69qO5vp0nfcQ/Dcn6NkpkiSJ8yyi0npJ1iuFw/s+cYBTWWDPM7NbAb
cU/60VrVISkc7hfr4fxpbM7R7Cz2TvVe6o+39aOCq/09yxQMm0x82OnZv/z4kUSZ
ogH2KBaMLYzWvTfPIc7i2Ij+H33dQJpC7DrBMiSoPHZbGrDFra7cUA6SHv9fmNFk
KNl/9+BmqU76lHtO7/dKGeD0UzVfXMHZ9HncDNWmwI0bd+XUBAt/C3gCeFdnHQrQ
HyFV+xVQQd+pXtebFgwyscr6PwxSJmTEfyIKPw+3HncdYp83zBxBRHpuu1h95aG9
t8qQV5uz377+sUX8+MOqrWVBnSeQ2GFlYOk9D1zaTM/K8g7WM03fICghnxUPWK/O
Ur/tc/Mdk81QAOz4+FfAzxN0EMAgdRupYymaZyMQV0KoTl/+onLTlAuX8aCAtRML
XOJbkGlc9XeBcOA05Y/oNmMTZrHK4U/Cs0xcb4Hk+SpuOMf2tPM9aRwAvD3tQcvE
DLbiXAO+xVpcJ01OoRJJb3LyNAe0VpmRYWI+7+XPbBPJdvbF1nPWAFs2GALmYgKo
2wsoDwpLLotOIN+qUkWwmsbXpwRAkhfZagBhhXVm/mdK2t6mv83Uen8QCNZs41/W
Li8RHHN1twKrx90SFIY3KIM/l2Dk3pNmWx2XBmSPQvxPI4GHZEA+yq3tMKpVCV6l
qe9IdG0esjM31K5yGYmdSJ/xOkRuOQzadtstE3lOOxoh7IBDtwOGytydLrbQRf37
zdQ7Ekdhfi5UcPVdxUvHRrLh2TSLFPBeIS4ewt0Pe74yJSdr7GzKqWZ/NO9UdGO4
dMSH0kXqP40C+L6/r54EuvmHDR+ZolbOUgDaVDW/cHK6TP1OhitbsCp3UG+J2VvW
rHlG2RSZ2F1+GwEvODi7K9OLKBQl+0xd9wVmb7yvGGicBPo5Iks0WNru/zG3Xmis
uZSo9SOGWM7bOfMBqJm97O0VOTUWJgCyhBIjHLLIR0FPOYgPYF23a7cMwGoieInJ
UrbGDQLlscSvrZPh+deD9bvXSTOTpyaz4N8H/D+kQwLPF8ee0E9ucVpSWCLiH5sy
M3jfj0lptUR9sftYovgHb5RNoe+nJKjJowgixYYDw2A6aIL48XISyItDmfIqVqO7
WUS6hFwW2nc+X6w4aipkBX+6R4McGdrAMqVMgVuXVSAmwhbW4dMQHeEL0iLjPA6i
g4BtFzNVvMPWJ4lD+QnCCMtojBaRTgHXKaMzDHgyYSTXAXt1kyHS0JQ5p/BNjdcD
hsqf1o6EvvJo0qm//5LlVBfhXslPdvv7tWpr3I5fyKH+MgX7sIsHIbvijF4x+0mB
ph/xRNLWXNd5gLvY2JpZX68vQF1Swfg9sOyOKq6rK5HCYBJT+8QPlbA3di2HE04d
5Iaxjl8rU7P3jA+FWnTZG+DQe8CX8sf+TKSBBLtXRNufEC/1LGZWqqBCR4UjMbDa
M6jCqiemNbPJpNdSftifQwHmNR0TGG0AYAfubrKE0hUq6TcFQ7QdR+/nbhfeQpkA
GqRpl9/WR+d5LpFUMCpfGzqAxdmlSNNC1ol6Gu/Sxg0iiY9JTMvNJq5GMbuwglyO
wku7hafYlCsTafBKa7ULGKq5FAvWYQwxOASNYBL2CrattPmjhT79nYn6K5VYYalL
6NRdsB52OBw6dskCFVPa+gSZVRAg7y0luLwijFtbNcP7VTqWL4O7PKkASobGqA9v
mW1/K1AqwXBObQmCKqQgfEjpsTyJluKQaFvl4WAA33uIMuPd8s+DQ+nbkZTJTFkx
onSfONycKEiBQndBvCvgzZC958eqc0zkrJxkAc6JNyhCOEBjBr5QePW3DPr5pG13
KRuefv5Y26NuewOqGX3UoUXwgJBk3zkStULgNWDFl8cV7TbfGetI4JTgI9ojcvk5
DR+HFOvnBm/a9+TM/KAhNiEl3/v/vrrtR3GILVaD62hJHU1FqClH/FIgLwjhjpFv
JyG2ExPMe4u2hXhqTemc4Bhlu+KmBB+jzDnzoXv9d90CIbEKVJfflxb06PSbDp4K
DseNkaXPsIG0v6OnnG/ueqJl4eSgiUFCkNqb7bUHJ6jtjFQeUROZIQJA0tr59wUR
lHkZbsmJF8YQ3//dhE89+bfhij4lO4/l8D4QtFKt0Y4nXgKtIV4ZwBRcMiYFjPsB
AoIYBg1+fi9ZPV+VKcgKvfHFCMXiqCyM4wuoRZeFBIo+m16qgedv2THb8MaRGFmL
4APv33x5Sjg4oanmXQjoIbho06EqBKtZqAGp68FcvnMuFiLFnOjrUfdIExLA9GmT
wAgpLyxLxVAmpafcYBsH3lMAhxc7qI1hURTSxBv9mWT+oeP7obqUzAq0EwmuLw0a
JnAow3BCPMdVCDgcF5YLuqqvQezQmy8C85n13Xse6OKB7Q0hdpigBt1PhkLrpiVS
or42spHZUiuYMhaEkqsbIus/x1N8OZkNrPGHmP7jJOM9wSH5NN4KxgAvkRbZJDDy
GpLj7a7cDLKR5+QoQicyAPuGDhxGhfTuYQzFoRhuBVKsSdtMNOA90ykGY2tm15hl
MzN1ywvZc67vtgqxqReDy1jBG/EifAQEasjXsBxZ1LGs+c3bMYKU0U2a44RHU1pB
b8IklGGmEuISzY1WpBV19xlrrNTOjgQrUTIYg0EiQR4igGVCzNhQc883pEMGgjaY
LN+x1jYNL3xb7XzSqIj2fYFvt+6dslHRuqpjcl38NU77Arlhom9FsHvTXMgpOXcl
tIzPrE6odlDVykagxkVAR9HAA3UizoVACuetAAEbQrD03CyW/I77VvtMtY/izPbq
pu0lFtVQe+gcaetLWd4BvIQTiRExTd27KQuCeMVzpZfMLXh9+H4UJ8YYH/Y19twX
I7SpWx2tjgweRgj8ADXawkS4uWubLrxCXgWO93Sg7diL/pCq7gRsV6aVBfqgpJ4p
nk8gl7ZIpDLenQHXXDYbxpv1ATLDkb6do981QBZBqS1dWRxNEnWtGR0FQ/JNpumN
yEAtEilNJ2a6/un1ywHY3YHovmgv1N8y/fSvMrN9ccjVKx/myDMRYjrd4WglPZQ+
uX3U3TQNEEo9ehqwwMidae9RMI8KpNJd+a42ZMd/+UD0aiFSYHYqXm/toYnxmozl
sKEaAWKbwspR9GrS8O5N3Zz2FDUw5Rw84ZlWtJ7YmHtE39W5IodQcPnqhotoAPu7
mmK5rjTmOsgqNJ6yAQmWgqMigY/3ioLDRLzYCHDSkmYLSm6x1RGAlGtm1r7eOvby
93v/Q23hHah3Gl3B4CEogb47a6mr5vOe0F2A3nSDhWBeTpQ2e7iqq5tdeH/K/7Lh
SIvocs7ouPNd4Oc14q45Z1gLIBilNR8+UizLHq8e2Wd8bK4G26RDFIq1y9J9rZUn
T7sa/6BXQo5WUqz4vikM0j4yR1QlKGS2j4tZR4mDHRNGNuHWaoxDpwCvbrzGZCZG
lT+tDsA7zXMsq3x9nXqRaaEi8jo7TwPRih0fXBrAft02cOQ5uiDaeQGPKfUdb3P7
3ZCyv3W9o0RtSWXUaX8AzAWvsAK2h8/XD5kFCBRtQgD2LmlxL2dE8U0qkyy/KtYa
kggVYKbNPCLB9JlRWzbvyMXSVj5ch3963Q3nyvDlglVyvfxICiBAvrJkSp+RIaAo
TemXhB8mX0VxwQAwnTGmILX6yhjBUCg1er6SSIlAJzOZ232jnf1PRuJr8U0WKCSH
Tek7fNHSPqLNGYrhSIwJB0OEhtZlRvJV/EYOCCq9PQI2hrCgS30TOMOcdLg2nA7X
1qWTFoXNdVK62BQ30vF7AEHVMz2evOWEfkQTpAfeaB9GrxbGrYjjFci3DU3UmEAv
JVArNqAK6shZat/OJ0Sy9wIfVGb0+X5UcVB89tH3RhsMmJunOpz2TJa16MQdjh4B
MGehb9fOPCmwsLTbcT/eLXL0kCisGvN5407k3GZZKK72f8ZaKfrYMP/6eAmqtJPy
TCbGV9Fv+O/YhVFu3epLb2itFffzq5scJXEZx3jAQpI4AKjXa2UkJs5egqoEthoK
mwtQCmoZxg79PJY3nkm4N6rg3Lzd+yVfWX9/eFPB77YOEF5RVPmH0fGftI/9s9sT
Ru4TxZL5mI8xbIgwxqRLkh/Hs+JztGDGGycLydC6cJHTMQH8IlSI4StBDp5b3ntD
Af16jEi3klWkb+j7CTX74RVfoZT7XIgeLSpvR8tRjA3VjxsYVlmB+ptBQ9jfrmAP
PgvM5WQilZctYivMKSFStrxKXEuPIn4LJeUDtykj/2k=
>>>>>>> main
`protect end_protected