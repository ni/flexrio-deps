`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
sD5jeIt/NS2+ECTgxO9JlvlAcP/79Lki+rJN3Rb2Wknr22ahAgu2GFf5zoPhIcGW
bfW+VZAPaAj4row4K8vIsoSLV5TVK7k6upvBGW6s4917oM1VIvbtFeludBrNhPqI
oNsGm769P9Fl6CaJDke2Tsgwtt0I3UhajQBYhp0EC1jZgEv0vUYOHh207CT+CgPu
h1lzjDOJpkgC3+KVtwRvDcPeayhoHFBBNCppk4j1oEL7R7eGMDf/ZlWLQy6qKssP
57b+JA10vcTMEpbviNbAzBU+fLTv9h9p0aJxf1NSKFf8joDgZ6rlBPIcigNbZOrM
a3SLydc88U7Av1PE3hmmC9zU6c0bHj8D/YYgnzf4adTeDpKWlbr1TtC1GghiJZhD
wD9Vz6xe3iRoZArNl1ImirKpoGKbyoUWEgL9DklIdLUZWDQg3GENBORLfdzxPXrb
KnOMI+flHnioZrN0A92EWH7yfkCJkFIn4U2Pp6ZEomKryy5OEiAjBUvNkkCmE6aZ
r1fiPROLJgu+OZ01dQMLmJzzJpNYRMQeyKoP8Yy2bHKLyRglhEFinHJL8MmD6rfy
PDzSIpbz0fNNOj/ktkL5xtLnStR9GhYoEnDYeD5QNsx8kKRLNPj1ES6JCHcbW+fw
1PCQ7rwmpV/Byg0sDI8z5/3CUp+L1ZQr1Yl1NAryyfW2nSNcnjRJC8G7HIzgXSpF
4+i+X+lIXi4uluzg65nds6tO4kNmF1cq+CXXM5dyyPB7wXAdv244c63gaZr824D2
l/8UQaUNfELRsZu1iNgaty4dhqelrFvVkXLQTBMZNE2KSRpEu1bcH4hTyYe2I/78
TMMzBmLEcIR/yOLR/Tbm7hN5+NsyBMfwlnRNLZ80GYcsmqn87vXmDvERri42xP+Z
WyezyMXsFBjn96jZVHR3G1DovgUPhqG1sQSfVK6Pq5KQ94Ndf1bj4BPo2DuaDfCk
Y3W+5AOYKk0s+YvWTmaXrdR8MGxMk6J61DzCcCuxSQVMen6LzcsZ0wiMeX5i6JYm
o0SKd+iX7VtC/cmy7rm59e3N55ae9QoYdPjI7L3kKGClw8OS/2uvUV0ogTZ79u9O
AhiXaZDJbh02aN6UJwhP//Z+klsxMsE6PNYKKIK0xYSoJ9nHwLvoEgDqngh1TXpz
CVmcAof/oZ6732CItLZ0EdINTDZVZJeTZnfdzudC71AC6FforJLk9bOigH6ijzCf
HuXpMUfpwFVGw84mRtEln/y3CvXZjNK+EkTyEtLZbnQqIFcjmIIs0ydsKXH/2fTH
pZvC3KJjN0yJd/KeNVRI0ylE2ZykHFLr9+PLry10snl03923ISAQzMZHbfMHu+ib
LOHFS3wNo2vkeNCmSBBMRawI6wSAsKQyIEVEUN9tAg0uwmWO27yKhIXdNOTnCpan
xpmhivthCznKhIDdE0pgp2vzcqmE+Ajs92QKIO+eUuIw+34gBZy1p8E8XnlEtXE9
wl2mvUaI7YjtNpuk1PtSyu7U0HEWRkZRXquhkhwNgRJJKYQ9ndj9zazN9Dw0tNfr
hyDzleqDUTP79l2GEU+xK0EBn197zUztgcnoj4ZNNbd2qwwlZAdvt66xNvT2Ou8O
GSgr/360GIv56FxakSAhOmHehj78ARSDt3Yb8pF4Ufb21O7uA3ffaf2/L7XkGBPL
HKmehKFv/wX65YaR6HB3erpN7Y/Q+L+L/v3HnX2B2KFoPgf76ukS4NX4y97DOgVD
hblhc3MqY94Dy1v2Ix2j4Ay/gW2cB5oYVlkesUH+liFYaJ4hv4H1pFhzHMlgnM7S
Cg0rcZvaXZw4/8v2dlLlu5sXWZyrwa4Z16grs0k12MQbDiwQBAMbqaOl+oY4p3/M
/d9j1EiirX1T+SgjufpyYcPJGo9azEZMjqj+Y72z3771ShFnyQ71ZPzbMngG/ElG
mOZa5vYdNdDirqo1mQ/rqpV59sgFUW4fM4SC1aSUqcH0MZNKhKRFhPXJai9K1vZN
jHbyJSRQF6rEoZZ2LqX5/A7JWl351RozYGJtAcI6ktZzYHrD8k9fDucV0nnNxCOW
Cf2vmhLPmAVWzrEvzjliG5szp+FPGMeR6LNy6951OzybKtXPJHzw6hMHUCQ0SNYk
KNjtOuB+jcwZFR+BuMekX+Ml0YVPgFjX/Kwg2pZbPVY=
`protect end_protected