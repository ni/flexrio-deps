`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
Niazd3hQVzwxL2j/Np2ydj25NcNZTMvAF1H8JWf/9yHMj3BJlXC9oPmZKM+hic+l
BWfAEbRdVExFaAoyU9T9Hv6d0d+mmiN2l2ZIaGXLsULDLJfoVjhbOuICW6hBsjqw
0Lv5tmFNxK6C6b005W33BNCY243LvbaAnTr/5URiLjV8+4Rwv1oZAO4CpkMl4+K6
nYsI9KzipEDCuTXbcCPtTuDmHGFWfPuybxz8FuzIwdkTvfr7hafpIlLDoSbUqcD/
SImthQfRj6wGImF0vpAzJvrlhnLz/9jgygbpwrSUCVkD7jyhiBvctPe34uLd908+
tIWyZnAWDhVe97/R+cZy93OZwwokTFN7LCN0+4S646vWrkZW6ooUrMQHIbralVTu
c9K3Fwl2yCGI61TBTcKdPAJHF7oI7WuWaVxHnkO8aJTS63Nh2EW3i1mgB1Kz3TBj
NaEwju6vYEbb/icBPSNITjVHLnhPV5ntqSusF+wY2iGiyVfKbo82UExtLHrprHxX
zRvEsiyPTrfM46bjsBvYJVSt7FjwD2fPF6wloHGxV5gnBlAoD5BkTVJcZogY0mxP
8a3+lnWtrWZGIWXWdyHD7SAayMr7/97ZjYD6HZRtCH0Oaw1r4wotu9MCUUi/7nFC
Lt2l9Q/ObUd+Oytqoymzj5QbY6PvaBMqirVacOfb6QlcKXRd/Z6FJKkOmNU2bzWh
FyjGf7NTIZAB/5sXmdx9vWAlxjCm3tDtXg1IfKlNg9kiqbOjsi+TH9e3ltFHDeoJ
kyS7snJ2xgiKMkRWYNY5Lpnp+lXKN2Bd8SKL6/u/lFCwxDJR0p+/kh2poqkH7TGN
+5lkwbaE4G1HFdx/ZA+OkCTwZvvA2KU7jH9lHmFO//dEYHW8YwzDqaXNCG2oX3Sw
GytyxssBloAPbMINTP/GAQMc2PCInXHVAZw6uEiEvYfSSQqKI29FRRDmQCZ8p4Nw
PNGMGZhB8ZC8uo2YZ0dzwZ5vX4T1vLbhvGawDAR7axKB7rq9ZFPDeC+/KIJojj9Z
c4C5X9csuy4G/GA3ZGiI+pQ2sWsw2DITpVrHkXZQ3N3+VQNys6DbJiuFcE+jPLa8
ycAZunXFoiJp7DwYX9Cwv+VPY7VikApntsSrtBUxLt0BGLHytyEPM8+taSMVjqi7
tNVkEQrj+3gPVGBscYeQasZXKT2t8NH50T8z6X4JWsa8CXeceQr613V7XfhvWqIg
IpoQhEv2HEDO3n7gANNAHXWokUUbCzznQzdSEE5kfB63i91sMijcJxOO0D0TxjT1
B3jR+eyu5iqD9TGoBTAbomewqfHpGNjoQhGl57VugwiFXsV0P7ZB1+sNhnE4OnIj
8kjYCvjbnBLICTxig7mcm2j7GQE/68K8ulEqsqsOGYLxO3Pr1mcoAGc6RxQVPuDT
NtK4CwiPvPejgs9KiVrbl7FifCBG+YDfe0PatvoMo92e4gTiHCUh+ARk8tRYjxAm
HPzwcfi/pryk+tzPrDwhDdjxUs0avm7PEbwoQZdn6KIMqPvGIo0OB6xvIYgHimNd
8c6umE0KJw8q24p7n0b4FtFkYpq+zfnTFQi0dLswPEZNOp1gRiFKfbjT7keZ5fn/
NcAo9D9Hc0Sypwl/UjkyMAoc/bKuNl4R4ekGQqyw70Tsky/wW0xgUBfnIHsCN87X
Da4XmX4c9cy9UsKDJPa8yL5LoiwA6cl7ySlHwPlS0OOXBYuW8GYiA9juBw97ImLk
bRwwAE/nihPadacPBDOHu+UZSdLVhKI2SnXCFv0MhgOqXh/46+CDE+iYaArG9kD3
4wnAhIpj8VPr6EkDQzql7t4fxrhJB6fy72At0McPNKbHE8luIhK1rwxe5DG9LybY
elXT3zO1gzNK+QboKbthQ9N+rnwWixsC0WrTPwzchyP935/It7tSmMkC6GbEUL2C
ztLyG2xcUbLsIWXmu7abZR2qF11Kxk0Jdui7+J2AxMQXIS9jJy2azdEVs+bdnTvT
BzWcuAR8mqTVCTkPVKlxwVN6jZUCNtH0WYXmzL3RwGboknwmxzoVzFvlB/8hO9Lx
zVkXDhEuQT9IjqjiT6iYM8Z1F9mtgV1QsegPNmgeD+R7Cw/h+5BUAk1AxSVfjgIN
/A4IBBjHyKTclykv3KIt11nk0fx2cltcb3kv/IIY9mQzcAFltJe7wpC62NmAjXX6
nywf0PEwD8RXF2txGlrGrMyGs5S9VbPqMNqlzd+Z3gvJ3XwDuTzfRKoKO75sPz1J
SkyYZAhtptg6B22v+hH6ifY1ZdpYiT3AqPIk6eGUpP5vPkV1qSEIGe+wod2HALCH
3TTGoac5b6nAGQb8KIVk6kVVHEoeLcyQcaakTFfFAVzKV5gOas59qCBf08Eyp99F
6uGaMHhkt8zjXkV3FqM/wvdGQliBTNXnUYvRJSdEqLMxf3vQRC11sApM7HjDx5Y6
7WsHUh9oPELcfbitUx1SROcf67EGDXd9nwssQTTg88XPLAYXePFhdu70Vf+AnNsy
B3j0rkQfztnyvOseMdmDVUWqVygLQ3nnr2VShJC7oSLXJjTNK6/ejMQC2/Uj3lt5
lMrd5CB61fYDkpqqgSCVjBYgZNqXWm5l4HOhJrisEDDw/CNzqQ60i6ZZh/NZQsUm
3JeVYoXwvr6k2dGtrm2qz+u9cy9nG/0NdQ3ta2jCYvUpUOWUtBLqRUT5CCY7IqBA
+ynZGK8p9S+IDCxxpECgy4kEFnawrmRGku7pmDflMNf1GKydxn4h2OjYiGIy5vUz
LVq0OI9tb1HKDFxSLPGqKy1m8Bxh+6UNjx9e3SNzSe0WtzQYK2ystpsTks5q8p4N
FzU79Nc3a2WAaLBqPsZgP4xlEIi1Yqn6RwVSKM7UJ36ogEZpvharmoyzGbAo5xmD
vxSwvNPhN5gguWyFeruTz8JAg18WSbNi4DJaRrzXeX5I/bKB5Bk+8Hp1SUgDh0E1
VR0WMNET7/I7U5y77120tTVXDeTwv3IqmkCrkrObvHKH8VSBGEhaG0MFxIbmA+2o
zmzdhSCC79hJnes80TlzY41XpDjfl0x51ieZGqIchiehAleIAOqQb+Ur5BCIX5j6
AAkk7O+SsNmC6M08sQGbvg3K97exx7o3Z4x6cqHkgqAZjFlO12vSTCp9ZjM5GcBU
iZjIMmSOVVagJgFk81nkQfXjA0Xcbsuta7pt8lHblkqIytRUeZnNUwKtxBfdkUh6
NF2PoTdDoeMmrhrjI1UOjqQ4p5n9vglWzfc4OFaC4ORjKKNolQzNLqLkRRvWVy4E
c7J5KzBlAoM/KAdYOUt0mVbNs7JlAnXjlqth1HVuUc8U6W3hM3y9tB4+0GSSFC2i
38ka2t5uzeqww9LK9A4BtewXneQnO+8HCdFbbkKQhoEwd30fIZVMt4N/+Etq/nse
m4XSeCJCwmyIJO8iNmAHEbYeY1NaKuNWSpDVrMQYdpYa0ByvrHV4vBrvkNitV1n3
GEMLieYpCujl4oKK0Zlq3lRR2T1575YzNOMwZY+4unWMLfMqmjULr8GjRZLVR8u8
VLn+V8/brZIpiaC7Ukx4feE8Oyy0BobGOCsaWQaZgciQFPVeUBQiDpNzdnMvd44x
vt7bqKh0yFBZXvbuhoj19oYuKhGtkCypjc+NXlvGgY/pvaUHV7gMZF4gC6DL5cU6
gSbvTWG2TG8YpXSI2lc8rz737qNIxnUIzO1sD28lDKfl9ZVbqmFkKrvTePrxKEHa
yP9/4YhJyyFizwoB3JGpxd0QTONLgCdAeCKw4XMwanRbpOCzMBPGoRUO+8eRjS1w
EPfpa1O6+bVAMd4r1HtDKiyFXilPn3/rZ6M+UrrbhejWqdVqcODvkT6VvnFXiEdC
cakF7TLqsZRFCXtQVTy3XPzln0KdJzxCfmUa7TA8PeckfzAbl7tZR4rzFI3OfFr/
/bxWu82w0o2pqlaxBHVcndnTW86DiLWJGbAOEBJ1r1K3Zt2xXDZ8Bq4bRlkyJBOh
y5SV+dyaabVV8n6fm6/FSkZSHnDJ/U1erfNOnDRXl7phr4SmjZBcpB0kDwAtFsHz
G0jwBap8Mwoh8aL17trm6MB1W9yJmqp6EKvAT7bf6dALBFurlTrINMlvmZNH4BQH
SrKG460bCU+r1vmocC9x9GBGruq05T6EGgz9+00+FkE3TCGdrQCdKKQZtm9ug/KJ
/OYTGf/Bx54BbU1pT3ScDTkphg8g49NXsG+tBKRhvjkBiNmhc0J0ceatggjIjEXV
pAvIjTg7MCieNXNCjivS8fw96I+Jha8YAeORU+OiHhlibHI93VbVFeBsxdZ1wjzm
028N4Oej/wWprlGO3nTV+MZOpfaHCDz1eDFUsoqQGsYENfZpbeuMm9Y6SBnlScZw
xr1vOS9/A1rfb2CYDrs/Y4fp4akawdRy2OFhi2TGu10oIYwzHF7RLwlC8iYZCFvK
c2WYqscjwxuaYj+d6BFM8HygbOhkLVzSGECgrvKkeL+yOtRknVGwAFLTVsI9oYgr
TOZeWNkPiD5eS/nw8Q0JxFYYM5+3tacN9WPMRpwZlDDgzOLMn7d5udE47lahc1sT
jOVBQijLNuPyZAOa5nDNmSDK1Gmm9LBOWLO0ve1D1Y4jZl4AWy8A5q/2e2JoWbWh
DuwKSSBwwGC72XWi0GPuJSl8GnwXDh852Q0P4gd4jsujIEjudxDnTp4erz80FYrJ
2ATZD8vgVHZbmRFBTj8VXBMt9+2kDUgyKaQ/4+56ni+kpozmb+KzpUAaOOB9vLyT
Pt4H0SF9ISiopxGT0cb1MsLsbWh68571kqP8D3bf1RiA+cewG87iEoQHCX+Xq0PX
aknR1gbzEPlQvRryiT9x7MfC21t8yFADi74nF7AMriacgiYkyi83t+snn9u0x1Ug
8JpylYBga5GQba6CPOkKSNC9mGjzhb7hd1UZy7GKHN8m26Wnwgibw3AH0TX+WRGC
NX12tBixVw8+HV8P/dUdcv3rwaikv0u2B1kGNPGONmdwmqOdFaiQKVdaQbgiPn/h
0Ct0mdbWjLptbcQVO25zTuMNPVR+qZtKXbx0N/HMOzWUg8AvCV1bYZj/DAhNfqcW
6ooAORQd2oCbhvsIBO8aqxdG2ENNmGuO9jxKRvEjbKwAR/JTK4UewqeE7vm8PXEO
j/erDypODDX5Ufb9JyHcyftwr/jK56iT6CYwSn0jjh4PdqGc3GwUX909QX7EX7r1
8WrOwQTIMdvueUUfMSLQg8tumr3TYWA7Hft2LLNOdXqyooueM5OZt796T2TTGO2u
4By4o8s6Bhn8iFCo/kirZ15oCufClrmdX4hhQRqdTix8y52UUXUXq1609836ZE0w
Ubg3dZ4X2mV261JBww5hHV1L6FMEm8l9BvgjdglrgVqlwIGf8366StLVvOVhUrdM
MUZP+hlnVaIu6dtH0zA0JmcN5Af9XybDJqwHdWLf8NHzOhY0tpeH9TBXHNpGPNMK
ee9pepuaTWN5kL9uprS/mngol6eoxymNPxGIBWA/Rd4Jd7KO4kI8y9KjCMAkbQlA
rLeCzEVHNp9x8LPjxB29Og1zERfKZz3EZf52i9T033RGpBij+8gyWaV/+yupyhr2
rHgnwQ+MfvDX5EkheEmfhXLJSJ76DAohREHZ3ve9+DcHSQdIzw4IAZOd1rpj+Ryp
sPnHu36a1Iw8XEcRLIZt8O9eEMOyGMMm3NfbGduaED50SBmhMTS5mfbSslD1KKHf
OhMIOpcdOEfouTTmiVIJN5FSIBjCOvr5bc5S6IOJfAkbHR8+1T+0eT+w4O/coBB9
pfJw2Qhx5TN2nylZa+zP5znW1aeMENOlPNrxQYnRNjCyNEnBZD0BvTmqXvanXTKB
Ao6Voe+iygMaIcLBFoLnpgXyIkJSYzt9i2QyuGUjNGpaTtVeS3GClXtgspi72AtB
iGkHBDcLCvVBPtX+P/QTJsEVSGpDpoGtLbJIzNqhJAdtDKPG8gNN41vM1AD3iSly
B/sl9q5dGkLuL8BrNTUfogFARMrhiF+Ae7zIQJAw8DS3QqZV7Etu5t22ClWWBbBV
sKAdrgaGmqwRrGQNR9wRC0V4l6T4NkgCdjXSo1MZcDFOWWYSsFDGnKytCEZTfwHm
00Cg9y2VtFAmOa3somb2QyT88YYQeFufVnD9qGKAxLnMhVEqPjuSBF6pQASM4Y9C
w/r6Ray72t5C0H/ny4cOWhuoGLkxSPBQ9U+FRzRDJI3fB+artUiRARHLJUwzDXvx
+xHLxWk3Uooq3evX56cLFKbCcAu//+1CR6TTqYY9hm6+Adiu2C+EXHPnR5EFTJTx
oJIR9yst6oYYdfOUsk+1805el1hlMf4SzKjgs09Thz8B6koK5igofW/qmLV9O5PF
26hlZNTiVw9hvvT2f6arPFLHW+BzgCyJ7sWREJ52mBUTVDZ2rSoQ6i1OwMjuR0aZ
ZJrL5vvG7N2xec8LdV2pj3GJ4eUNySp7PN5RmruC2uHE3sPnT4e+RgiyochDArEo
2uOXOsPMR1R/rNf6eKQMVAEXmzHkL0ZdhrjoSk/e24P8mK3NQR6xmnBwoMmDMVSD
y8QCTupH0//lpgjWon+8Ohm50DBdmpwXyT0VW7LP+ZQvOiKADGQBbmHTSDTmqOcm
h4pyMWmXYsNpLNCjinBlln4p4T18Utyj/55AqSzZz40XqLf1Z8cgMctsC4yBXma7
oq6B+jnNtFAPeGkET5O49ymSQ6IDXozwux6wiIgIrMUx4ictWYuuDck6rKlKEhon
BFvkJiTMcTAxcZQywfescCn/3GpLA/0nOCDVPrs75SnvJxaX85bBRl1vU1aAHv0t
eatGCoH5IC+G+ojzaYBbN46UZreMFXD0PYezba4nIIDZLNihcj6mOtO/+71KbIOp
LTgUep+kK8jIZEwhic3VQweF/mgb3hQ52FXrBearGgH3CX+jYyyO7KALSBFTLgFb
6JdhUFBRN26Nnvc/fqfx2sM0x5vz8o5cWCFnt9+7l3vocrge9lvqsFRDt0zSluw3
JfJz71NuQn1LTMVeEqbgkEZ+9nm8BWFA2xKnvVYKwOemYNOcaBuZoo6+v8vj0MlQ
qtXQNEnnKDZEyOxAPhbcwG58Xr9pU8qgCdZ1peeqf2f4BfG9jQzFEjouLv3k7wZD
GOxGzhE6Gk5Ntq1186tovfCnqwxafynzG7sE6XZwasjhNBvgSaWBOJqt65H/9t8K
pVIsAJTGVumNWWXD7TgKlioJFxbUyeu67l3WV+PYf+bmMMHbJV41xF0zQfDSfi+D
UBcAZ/OKsB0cHdmlZuKCGzjhGXA90/CWLmuQhD14H/8PSRmU/n620kwF4xLtPJZb
6PhMj0AUlsxG2S8tHP21m9/onAHhclIhOsDjDc5s1Y8asbxBZuqdIVNO5gv2J90g
MsvZuvbxdJSNXeaOW8eK7mLXnuIJVyJtFm7K01MK+GL0jOFhRH7ZMz01eo7LSBBs
TAVgJyDZhAJAJCLw8Boz6S8fYp5NVjiNDZq+ww3sq22xGvagfo1ykNlncl07fOzd
50w38p3mz+Gr7qPH1U71+u4C7ei7vdPbhFJzbaCYwnMGNlYxXoJyBcLXntHT0dZv
xwPfTZAe528lI3FHrY973ANgZye9UmSpHgK92rfI1tHxi4DfIe5CULtPEXYhz9NR
CdznyPpBcKOQf67hETHT+KLR9XgFfQ5zo+RNTQ3Hj5IByCQR4jBQ5i4ZGReDmBLA
GhJH+EfxSHLd+zty/1w0FGUT+yo7goyltBLWRlRPpdy9imb58Q6E0fotg7l73AyB
0kdjjnoW+YvWWICn7zY0csEreLNwfXBxXw9tO7HW28My+sdHqDeTCpDFDkJ+4h4K
5La6NA1Fv2PC0YHT6FSqUVI8KmAg6Lw7g4KbvSlRNSYudsPYA+89QvGwdDhQp5nj
CgAWuZZYPs3cdelMF71VVRDzH77u9HSgeeaCUOV81RwNI/fbImvAKcu6F6klzR2I
cOoangrL9qLGakEWoEl6ZboisFTg4iAHVSAbiwMtJrFJXc7xstG9vVJFgru+RlCC
EqjqqC1KvbY7gMfc/DYXc+rox9ukJN+U2M1wYfolRX5v4XNtRIBaOXe4ui7T2211
MYQcLqE6M6UNtovMpqRHnbtOV7vwD8RPWxUf593uxAx068Eo28Ve6uBfQcTl2LTU
MB4JEUkjuk5ys6R6iUcqhHe2E3yb//qcK/M+YTqsMX+MR7s4xbc54fzY2IWA1KKK
TcugX+XXsG56sunMka79YZCrX0L6SvrhATOM9P/f5C43/c5XPbxEGSeIX+8lVJ5i
wXJ/OqDiuAjzdMzqH2qzF6xCoh2Z12Fo9rM8bpiUpEo0bAJO5FvBB1pkfdcZzeWB
MEpXKT0wisoxi47ETAPK2C46ZluQjGNUtnqN7pejTxeYaoBRRGYpGi1KsVFtliPd
fYN0haDJF59PpBr82DK6otVemDQhOKmAcM2GPMQeYGTjn2ClamCYLfkUyXGchEjO
usTWuwvMD5wWnWETXxvZGoMZLQbd9XkPQiPdMZruZ63NBblXv/spd1HAE3gzQCLl
qkmoY0xlQZvczmz3M9H245k933xiOCH6/gtrbhrKdJiSMSyOiH4CmjMJazkjRnv/
onpEPj0QKsRE9xUKBpAWy28PZHLgbJnLhNuS4goDon0ua+t1sLiOgDZJRVWJZraI
jJNGhQcUVcncFPn6Mkg31BZONNDmyLiAzJ7aSnTaUfsUnBUgGGUanK+Of3iBioPp
a2Xpsg7AgTiAy+dRHRmzGJYiPGDVWtDZXQ50rHo8u3h6NaIChmOra+d51U0Px1QG
VWxLyEMg3enbob2V469Pq+Zlfs6LphHiyi+F3+RtX+PCj7Gx+2J+sbebhXqX7Mee
LSL7F/FhJruV7MVIyBMdfwRc7DjKQn1qbStEkvyiGyxI/p516PAd+w96u1e91C9X
cm3ABqzYuq5NDZ7x8k0+Ykb6WBtrMvPOSYy2c7gQ66IK6wl+GjOu/B/6XJGH4IEX
UdkrhhmQ/EAcTjedehoZ4HbcHKccJ96IgYHs1tNufQXly5dj+db/YOLpGJf7RAft
iULLMe+6ltfeXO5zRzBjQq1CD6xVTvu3/m2lRFtUd2Iv0d3it2wUgo6++iKfkR+/
BKt1yCdv3Jl+6lFUY7HbqSWYEVt451yN6qOl7xOKkVSukNX5W2D2eXI9IQBS1Vyq
eToDGw6VQwzktcgrcBk8QUrqAeY3hdHX+U/zIfuHmQGPAtdNA5EWdNYS4o3r80q8
XDuvMJs6VEmY07WhOto8JeqBOqkBY7S+WIptRMCYFHY1yaPhGhudGVzgNnkzDRo4
e+WHHMtK6qNTgefYc2g7Yk+3tWzddEUqFBsSpjE16+bYSA5fEvLNaTvS8eOidnx5
qAjY8XAttg31A8UIgBDfpp0tQJa8H2T94EJQuX+5LWE4xzW4E++p75m13mW5S2cF
By2e4ox3n5WM6/cHEcwMOXzYg9m57ffFJf4Mwk8WxrRzEzbVxlYtuabrOaAeWoD1
j8EC/jszVx3D9E7crUpW5Sen2q6ibrgmjeuFlRqfDnj6fPUbZjodVvEYe+59FWrg
VNh1cAasRi2b+DymC4BExa9y2R6CDZLP6KoIV03GUrZWKFIX0zk810cXF48emIyx
lBilPFLAZT0cT9RrHNeXxKbEFctEHqQD+oGnY36W1eTE5ToqntiB2qk0R8MdOrLK
Ekwpv6GN+HZEBeeXuVOmHWePC7ewxj3Iw5rYAkTxiaOaZDeL5alXIMG+RerZpSOF
wXVh9QoY1FFRPHDrjCDa+l9ctThbyVYacet3WXqV6vZL1CF7ZNtWk4BxnA0HuSbh
bwSi3wUmCo6p1E4wIQXSHYwTvhjKIkZeOhY0rSIl4+Nxl3kur3VZ2yf4QyyaYwm4
CdqvlDLjPEc0KJivp1BFsO5tmHL/IQlY6uorEwTsRmQCmct22Dowd4hXzN2oAnTL
0S0Uzhr0S28ec3uJ0obkkqRg8szXwMbcYsef/Sx6kkHrpXVt/mPgDTgyzR2vRU07
Y3bBPcWUbx+PfUsulk7e0fPD54kkkBzSdqsSsrjpPjLvBp7p4p5jDGJCikuWsDfH
TZCypjkjOYH5FHwifXTDRWCXKHfgm9gkGvIYDreYDr015ktIQZqpTG1QPhiBp1ez
w6d5rIrtZP9cM3Pqr58R0teIH3nprbIRz4h6kN7vcD2+YFkou4Ne9dmdTOqaIVE/
wdM0bf+d/zeB7oaiay2pdbUADWjOa+AFKYs1V7ncNZJup8fxvm1C8ySQ1VKgYLIA
BJtKafys280R1o72j+Dbto82NZChbf7rg/r+DMECHktQZCnC792OkPS60A7ymluw
heBdB1lZ9hl5edcJg5PZfawK+xmKeGSWqWnRqiMo1qCstjOppm9OB7tFecIlNX3N
E3VW02Fej9YVdFcGGVv4gG/C12l9D+kxC0w4/GnnRLVigFkp++kbsMp83vukdJDM
tSarP5Q7nNMJRI91TNsHWdTRzwn2NiBZ3cd5/yyE1gNrjZ/BAe294kHzbQSHT0uy
bHBoKInZkAVoG5eaoJSyfx0WlHwXHxPgAHac/vUUTiWS8yuQJRQYy02ZVu9yfGyb
MxUSBz8K/8LLPQmEWhADrJy2cHYrHOgU85+TVRXi7SUy6d1dyU6JR0ZYo6FrSDHG
9f19JVzJ1aJwCsClZayxed42p6aNpTzbSq8QdEqQ+C32wLfTCeOTTI2nSgkPkmOn
fvWTQ9Fjes/c99QpyItqJLw80LjXrOcY5t5Aiq9KAvwXPoaaUBwY1Q2UCSEg09Ih
5j8KkWTwc2Gux2qC/+8Y9Y6HFDqcZhja1F6gizVy2yNgmMdioowkBoV7K666WGAK
emOGZivgmSecW6cbiKcW0iM2fnBrcQzQBbMSmcArqpTlXugM5DwcYQgm8XTz858L
nknbzOCh4XnTdBYUO9wl5yPcMPH7bMkh+GlizzhwJfAm67qm7OCoWx/jw9CsKSva
1Aw8L6B5Y2A88mHQhZCsEWA3+8NCvROnRsFlcnp1xDrj8YXy5LPBARVsUVjCi8DZ
xlGHP0okBQuEsdnf322CzYI9UcKZnAVY3Uaikv+vGfCIDGa15ZEr6dwtYSf8zVFQ
PRrSEKkCXTTbO+4R3SPxLARBf7gfOYqCqAPBT2+zfYOc9qp5WCkd5boE00yCoz/5
A4jvZNDBV3EN9VFnV6R7c6G3RDkYCvCYzC/A5gMYWIz/HTer1PndyYsWw492p9i/
NLVkwOSF7PzWSJ/nJ6AMxGmyQUjas5rSEuG6Tsn+a8fh5iFhTJ7SiEwgmnj3PnVq
h2OEpLY2ez694T8bch7vAZ1fOrZpVvSKabdJoZ7Wsu2GI8KtEpdO+7IkOo6yTtQJ
2XPyBkB/PmbkqOJAckaOklz8Oml2W01ocDWzQCvIKKhhg+4R1bZbS9D3b4I8GEc7
Hjwpf3Ojw6SUEekEBJoEoi8+KzrT/imuNMqDtlhKMhKALCfmi1JUm7QdX/f1QkIU
4kkkzIs/C0x2BVm8VDK7Mker2o7Lpf95ypGWxtC085PagpWalZWnrp6OMS0oos4P
DEz4RanmXO74euyPWnJ0BySHUpZdg2LiOgo8Ju4TUjp4JG0c0vE2tQsrihscPh6A
+LVWYuH7cK2lY5kzNmOcaCwMVeW8VXPxI7MLh6N1h/zsASclM38BgEYpiZnEQjGH
hqFInv6FdcxgcKjuAJLFJWzTmgf9tUnEQaZFujk7oHGrNpdr5J1ytoHyvXSySfro
dvsi3aEV7jbB/SpVjqm3ncnmLwHpm7TwKgu3BDhww0r5dcknnTrwdKuMA2cTW8eg
r70VM/RhLme0i8IKQG8b9qZbdXezZ+bwLGKUEc2kQTFiCafKDsy2DWJpANFQhe72
2n8zmOpyzl9qAITbUzOUXzQahwrLHWxuzIr/VNsMMHx7zzLPU2Y4xN5LdAGELu/r
gu8yyTmPFuWe7zqvFvLo+kU5ML6XmkiqcXS4GVDtFWagAZqADOxBUJX1WCBFxnc2
BbDJhKganFPI1A3qiExDsFrO46kIMaHmNKFXfd6dAFs8EZNQYbwas40mzkQeTwFg
AsFEhNd1Mu7N8BkaBaKWf5MrHh/prjH2KjweGDIe6PxBN9iJ5kHcbAKyZXxPclZy
24xbOxoREZgvO0AAtp9lftTj0qKtbzMtJaDHhvF8YQ5r6h3wdFjcc9tGdufJi1dH
M/IiLmlL7YszN20BEYpm3UURwQ0bdx3rzMQCw3dBoDaSFDqKZvFtqxEDDzOmKDe+
4fkUJrOB9ckTXxpoXyRm9h/V6OVjTaSkJPcIKgMDd8f5f5TbYW/ZLvmM7+q4O4DQ
O/EgTRR8TW7M8OUL8vIHN6LWdX/ZdgNti09cMqRyELGlo6FtM+ZSx1iz6MgoBipR
cY9/EAmfH+zRIfWXUSe2JSxObPDGD105pIMrclfAFTiZQlEHzUi/ICVonsghWXVW
1qyP+qQlTLGJ6yowlj6EhNqnsVmXxryfMb11UznbGT2WK5zIEpfvdxnaWfNb3L3N
xPZ1k7nftonveiACHzRYxbMNPWHv6on4JVMlmTRCifO+eBzot2XpXaW5wAGla8sj
SfADY3csH2obFbhp13TI472ARm9eDEejZ/cBXa3EsMiJJKAW63Wp7mO+NtXZCVzD
6tmvYg42EHRFXbALSd6wQGKyoRr2NCaXvXYF2z6+IiA9XmtfLBb564iQUrYng01G
oOTBvYEcPkpNYBN/HyG3CGktreaED748gFMQanleWUM3bS29xmhs9JOg2ZTL+o4r
qD3xEA+B1hFcYP5FmRoDqLSGxyUkFUqm/dOoQCSHV4nKEGnplXMc+6z/lXE+keiG
lsbC4kB0uOfaaLl/l8o9ExQ4DvMz11zmupJfD7UMXcB48UbSEhgLHMDxbaXWy+tQ
NTjV7Ak4ZXCvtnjm/wdBSbK7NosanHxrY/TOJgPPb9y94Lr3baPn3VbH2EzM/aPB
FWkaRgVmLSJU8vwU/KT4rWZHaIeoW9YIP8zgJSh8+xk52j6wO9pqb3/5gq7+oPRQ
J/WL57DR8bb+8nybNGIfacdyKLgs9nKs1UZETtZY3A9UC0mxTqzKsPpasiXpdy1M
G9b4PDZarthaBI4X9ZcpE9m3w6ZwqYdtTSs5fkJSP+zsPcW7oprJapEbJJpTG18O
jaI4KqT5ZgYd8teQ/RFvrLopCfTcRqtH/csfevaQoLloorrV3w69iXVnh3pRRxxb
bla1lbNdhhs45FjlPdlUlbZRpTpIl+Ozzvb1rHtY9vbXSpWOiFmjGzz5NvCfS/hR
HEPHkorzIy81BFeriTIH4eWAXpBdXCd9bOX67FoEj0zxWfC35aD4EFEENR+1rg3h
XGDBqWVgGsJd89838/Vyousmxa0RzSpZL2hMhElA34fCR8q+S05TiCURAyUQLhwm
I478ZhW6ts41ZHjAbTmAcMssEDd9O0wVHVYgKcZqozSdl2E3TBpdrXjlnj18YUWm
rv3RFgsIf1kZlZ4E7HbtzWuYLzrCVGs9CZxoMxCcUi1Q9sFdG4Xc4GXsrSs02cI8
9PdxvU3rbKe3RWQV6QDSoqUdaU69LVBi7OyC9BctgDE/8LRF+U8s6JZ1AGJR4QNd
ZbERdGzG+o9EV4pD9YNcJSt0f4UiuXvj6Zs2TTfZEk4wMbrbogu/WBk9sH0/0FK/
M99bHsEnNPQcb1SP4US/qcrmkA3tFJTbvb+ylBiPOHYpWqOHxvDFHfup+V7vf4i+
mtsag4626i2ZqcGOwhmj4bicDwyo5jTXQRtW8Hh9X0TKG4leB4OSHMc7h4BR4o35
z8qZS81CoyFvLGWAcZhe/NmPWia8EHDGbGQ890wwFYssnNh/Nyb7DgoLvCsg6DfY
aw3325pag/xqNHYDvF6uDMzvdI4+V3EGRsXXpLGLgXgh2NxONJGBKbCQ+NJF7KuN
6X8lV+uLxhXpDwEzchSidZVuz3W5rp08Drssa+kJ3BOgMNMPhk1K7SopxiIcYxjD
PHbnROhI42VOawV+tIHuvgtyBlNEfLP/12OAhlAj3X8Jy+pibMTh3jbDGVtk9Tmu
KpXGFrUMgT3el6PhUOdbSDf4df55umqjXOCTcp4C9Uf/WNvqxX6RYj5RktIDb7lm
vaw2yroIJnk3BjRA5kexkw95K4e09/3gUE/NvRuC4yThNWR8oiCafAx26IZaJl+K
NMm4FOzV5fs5dpbgH3lZp+ZE2kZk9j9/8PRd3xLFLDGuzEcEUKQ4Lk7CZjdi9vW4
ntKB5ofEF7Uv1qe9es1i5eRtznWvDXF14uMf+nwea2EmMy+QXHUOhC5kIX8vySgg
ICrTjukRPDqu9+AjGfTt4WWxjAnG5LEOkRO9G6a/5mL4VVOuY8HrAG0aYbVkjZeu
EWlDzQaaZrCsw+YtZ6gT/G3JVOMp8WkxCmCILvvoSqDqUNMswIwLSRW1+LQ7Oc+I
uCsW0JidaeYe6bsbYJef5MPT0Ky+oLBU9XnAUhRS3Gym1AM21Vn2EdXyPWY1rFUN
LHCO4IZGWpI+yUiZrbEsHNsH9Cx0wx6LqxPmLXmdUp7VafU7YgUhqA74qKJduiXQ
QU3OHgrN0tu4Her0KnEYEFBem6ftGPOXT0EWlocSapZ8HCOvMj0gW38e6Sbtgak2
Ayv9bIW40RDzChPgkPnrQ4rLlC02PkAdXC6qRNUUHucTRBF3PxygpDgBcpWHrsjQ
697Oml7ky1UPbtn1x7FHuWV5WBNzqo4E/yKa6n/QEoOwdh5Ds/gHPVRpGLv12XuH
9vMuquGJ5hMmuAWBJo1gjDbbDuZY9ANeU2ydVesuhTsfeg7SwagmWXJkWfijXm6z
LGADtnEJ6oejpUDMNK2NntxFsGgj7S2rYDZh7K9Ypj5188f+NFRvReR70rMQJa1e
Kk4Kt/ImyFER6BOLxmZ0uu4iJwsKg7vr+Q3QxGTiF5Kknih0PvHYySkxbyrA17wi
tM2K80c5KTSUmTV9g66KsIigqhxL/92wKk70oy5wOzuNGBcBOtORihXFVzxTKyi1
SeQfqLq1jRLXncu9wTc7g0OeKaZYQWM2NHRdtnZurmtd82iJHBh4bogDkdc5KuFw
vEDDnGVD/cdrxyDv6XcG08td/Kv7PfyPCZFS8Von+4JmFaUKjJ6HbxxFt0FJpzLE
vt8i9I11pRbgiEWprOARBPNM5eSct1aeRlURVqXtW1Jh9bIVx+7gqek66QA5LuuC
GRzIiR7ZZ4jLLShWN77fO87WsygaC08AEafggZsnJ2vJlmUN4PzFDdjqfWmqBrCj
GMEfRhNERrfmKMS2nHikHXVCIDtERQHkQKK9Pf4Ji/SCBwEp6ENp/HVknATBcrtK
rqHedSN7vhSRT7hpGwd4qqrV02+/NtDcasuVMjqnqLqo6bxLXSsHLkfsgoFuCaGD
tY8ZiDXuObfCUwHkivPCPiGqCB+yGFmg62rWenI7Zd/zSIlK2YmcWi4TMDQSxFX/
HyyCKp/MPPvb5e8uKLyA5M4nLXj7nm4H8tztph4/YOiK7P6F9vNYeDXpI77SKGkv
ChRFHK8i/9GPJEG1xPlR7SoVQcMlwufig1nhghv4eLjuZRKxmSImuHxRgxgABXkH
qtEBbF4vAvMr8Jyl8WqvrkgPmPNZVQfVkvCQa76bgyqUB9V56oZXsWgtGuNTgrkC
MGZjyr8NPva2bo3dW2gvvyRisVgh9E9P+5Iw/5OmQFrAPoLWrMw21ShRblQZK9GR
Hk6gHDB93SxeU6aDwB1niiKYEMbJ1kDhvRwejlJoFxbBMIOmrxZ7Dgw+Zz0Y+n2x
xox8XLSC4iyVdzux5vAoA/jE6DIgi5N56qXa4mAz84RnjtIfOMDmvyIF4lLSHQuA
qeXcdVwTatA+JLMP5nLQVnZnl3OhbVkgWmRc09Bzl23MK8uHL8PgLg5d3EWrAmkR
jCBn+7K0M+dHsY3DjOxQ146IIVbmU3D60WZGt2uvP46Nk34iMSDYny01gC2z5yvH
lbX9dEeyrdTsiWqYy5d3+RAwq8BDzfaUYqHJM0vcWqCQRG4tIhO7NDSWB4D96Nn6
udx87fs7QY9YGZe7J4Fz7zAw1lylrEG8Tl0qYldibj2+Zppq+lzzQk3tcDfsdjAP
ir2cajg8qgupqJ6IGN4ZIObCR6FnJT4wZoYPhayTycpPaZBsu6qDcpN5krdANkmq
LAmYppPMA17px5IB3Nw2LzO7vJme1a4/pymxRHaS/SgnnIQMCM68Dd9LesJNYBiT
b9wDBYxaKJ3lPfC2oUpUJtleoJmZNum3KCg6K0sCAxNSMaWKDJr8+wuIMvCXu/oi
8jMc1mX5HTw0tiMJtqbZJH6Lszu3Ha3JkuB2QjbPqM7FuMaIPE+Dl3MOC4QagpoM
wVyxrg3RZ8wyjLogKGgmNk99WkDTJ2J56RkYveOF+bdefzWnYVnx3qLMCMUzEVW2
7zXcqQ/3++LboMrQ8D55YbNwpDGrfQiNxsGJ8nB4+jWsO6wg0Hig36RmyESMJKc8
RA384TyPSRFAkfFbQcL1tW3c4g+cMqDNmQKSwINSuRJwivxScEIuiCNbFoP13KRv
rjvjr6n1017REF2hJ4MkbTi6aagAYzAZRSconk1HJQnc+MPsvb0tIa0cpTpKFOZ7
CGZsaN5hLo+SzQsq5K3KfSaMAlK9z9p6my9eyNcbTXommWMukrq4FJAGkGhURmMs
9gdzl5nsWnbGRhD9y3ioV3xr9aduy1SyWC/3iwijXy7lLrQwspHJNni+e450fzdi
NTeBURwiWfWxYP7W8HkcyWRIFBrdEyXmer4Ep6elRgy/bEuWSpqAHqcNXhmO9xvd
AarHHRJ/FBYKdsjJkjA36lpipsgHQcA5EK8eVHA7axbmNMqIgCtiCI6cfpXdDEvc
tqhcBOENC6DModC/FBx4J1Zx3azDo1+QIYkVrh2D8OIa3uLkmGSNjJVIFD/9iqgi
rjcbWhBMn1yRHPfX5R6L4214OR2X7IsCKwcDrquq6e5MIYifBVvrI8c40tZ8KKoY
CDIJyMrar+YIh1TRtEqLbCZdwNYQngIQHczk3hUobfASK6pzMWCgyS0JRQzFHs7m
i3GRzGw1x8hDstAqBf8gd/RuOdhv6nufKvcgSEFion9zuyqdxiituBK58RvtTj/W
4fWDVvv1PHWFMLXUD5uyosmEZRv146nRr8uE63psOQfLrQrxUIxpF3alcq/3eBFM
aMEC1gJbz75zAfzMMxudZhQHG1zWLYweu4s62mHmWZ9Ph+i4ti1dLPXCtsfbP5TZ
KV+M0xZ+Zty79zIIgpXqMYRL7ieyKf9prbroQblnrmNWr94octt/QBivyuLUauhI
KdyPr/LjRQVhF3p0d6Z3QceSzdtohRSQtBUnNPjToQN7E1eS6fDitWtbi20/3zlf
8vqqkirnlNlVEWVAU6bZT9qgyRqumOMbJFllhXRfGbDXyC0Tq2W0zLdNaep8DOIk
x9hUaDAFyQHzi2eiigy2jDXl2vXklYnFrVqSb/hm5ULZ6FPsJUydCIUrxhXBW01S
CIDBnTaWDvA/TLGC1FeedmnVzIJmSaLOakmx1g9oHjgTm7rA0qoCXXqyzsN1NDlp
dQ5q0+X07p/mKB3oR9Orkk9ik6sRep3/ji7wB9JTfaq2nMVdQSnE6TjSBMipMPHm
mCgXEPkgZQkEUlUWrddj/MqtfrFWoHknETDJT3cNzjGw9lFMgKiFbwtkI7Nw7JMW
IsNZKf3uLGNR04XrhEErJOLDtqU3+FeCYyRjK6Ix2nFNN4JtaowHaCJlWgu38T6s
aOaK70VWBy8ntmNjXcBIxO62YXa3p3txAmGw5qfe0D+gRvP+bBbX9t73F3JIiGjl
XXYDYz4OBVhcckaaMyPOu78LuN+DE2ED1E3MiieR2aJGnX2kMj/BV8m668uPZl9U
Z0+0+DAxy1wjBnYe1UWMdZnpGFAaUia9UR17mt5v1lvVlQNdPHTMMsFF2tc1xIZu
cLV4bRyPwjl/5weurL8KCAgSSZDqtbjG7B+NYkJoNaIude+uKAakjdeOqse0f4wD
bpacALUdyx4XNABqjiOmGG+Uhm0JyVHHR4Rpq+LvHUfR7dhVWj1KTtVJyCs5/MZP
qOeM3bc115Vf/MN3mfoN+hEXynXQ78YGV7Jkug0BTbtV6Rh4H8TLqPdLXJzYZ5LU
T83YB0OysnCvl6IaOQ+hJTYQW2oJIxM4IPWsfzWxTqA6mrX71MZHLui+BrzLSKhH
rYIGYEm4wY3VTKHADOfn+m9Doplcn8S0wLHCH+3gMxzIP+pbX5GnccNnu/Y9i2zg
gOLdAi/p5UwpBpG/Kd8CvnBjZO+IVxcx8+2waTfCm4Lad2d49ezuV/+oMlgfElJ2
nCAc6IF56yRxzMl2HnbE9npOXeW3kxpS7oDb6vQqSCaLtpb/vV4oOk+56jZi47mC
4zK2wZddGifmX0r92VMUCr8VPaP0JpCHLM5+0UDOjwawSrJAX2iKVo23WIJkAvud
e6780TxHyZ/OxBKNcP968N3nAuecIyyHprwPJKbvm8q2UQJJX/xfNF73Z+KQgSjB
BHA8ItoWS1dYkelvnhM2qKHgMmP2IGnRQIFHBrFrEpL1Sg+a/rC3HpOAZxjnQxY1
PoAWGrdNzsGylAUJ+Pk03WY72Y/jkCV+odtiLy9jL2mYgNI1AWJ3yOTgQVWZz1sF
1qfNP/zX3KEG6GynGg4le3WkWSQ74BUd+HGQX3BxNazKUdTFN40U0bLcaRLuqIV9
P4N4SRZRJ3lV8TbjXgBZZmX137plTwdmGl0FdvV6LQSquiVl+EQWHpuSFntCsI0c
+L/7jWAmS1h8FIHjCaQXwH7bwJXs8F7QcqnaUO7SvQGADpW4NEqM/z7Y1RXYX8Jc
sf4snhvVuroS0uf6SpGhHQIp1SdRLhDQtRTgVsjRwOTANbm62b3kMifWNaUJcPqc
CElSygL1GNnP2LKIA0Ebk/5hiQp2UqVyePh8FcFAq2GM0gq4Trc5YDSg4AGWeQ0P
UYFr5BC6bA5fUMVssxHmVVXtte70a+eZC/Ndt9CeLi88caHWn3vRZcKcXdlhkOL/
qKbDJND3jXLXvDQUh147XQpg2DNzST83DKf7iyc7L5QzvTR2MX35+RwQ4LgbnvVI
33QyiD2WPrZj6nzzYj/v7//YD3r8H5Ye7Ndlhy9RGUWuOTsNYbj3oMk05DDrtBOP
Q7owfVRrCLgDAjTSsk2UqDdgtJek25VSrqPMuHf9Odh3DC+y0Tksvmen4IDMYJw8
4/ohWujJmpZEjRfifsBYY96DM7flygW2duzTTzDHoBcGS0gR+yIBpeElULDrOsSQ
7Ppmy3AzWYu5AIJL//Xlm2yh639WxvMI/C8Ivq5bXOBeF0LnOQ6AJ9ghb3lU4Css
HbS8mBZtz5JKl8WRk/F1gzHyx84xJjBfbYjT9XWVyhs9bSV/YZ/+M0nkTMK/3dZN
blp3XS2TWMGKRjSJYPQZzZuHsQNxNCPvP17F5ccFcdj7qLB7q+6UO33aNpc/qDvO
BbQ3AVEzSYDUboY4+icQgolnZyBqU64QksFCaVLeidwKFzFxryouRCv8H/5lykvV
B6w3+5wcmqeSl4iQIC7wO+ewLRpRImd3FV+rDqRNGDzuizUY67/e3qDktZNLnMoh
ptM0qcZ7POBI+cf3FEer/WI04S7JHkwtPNypLQVS1xGlrdSaQNGY/8Oi1rOWPTLZ
A/pTNqf24y56p1Jp/K1RaNm/UuejBN3prC0xt4KwtFPmOcjV/qTVRxQYnMD4QIqb
Zl7t1E5rjn71DTdtjip2cxxKA38ruDcPX9BuTcs3Pyt9cXW7xBn/oW3nnNNtH2Cv
DFgNmHhSIiROnTrNOldtznp/j1ladqNKSVWXKfgtpFArzYSWNcoxOlAhmleiNE2F
YG1GtFK98c/IdWJ405184EK429UY2Mo+QZHEO+oyLzoI9aUh/2gSrO++HAgbfjsg
eGfk+WJcMvNPP77E3ylJCFlwO3x7cW45qLcGsoATU5OzfD489uQ5hC7mua9ZSSiF
n+gQWjQlM15PQhaIIyYvLScozvE/QGu9xwpUkP05D/sYhSAkw1dnNArfFUpFvOa5
Ft2qL5nEQc8f/uPZ1ZAPEQpuyylVPHPGT8nwPQaFYIN9tmfABnSisV+3zGUfezvX
3A2iEOm9/AUWT2iQKCMOBpb/+Za/1dTt8XB2XhVm/z/DwWKlIealsnZBR8cRLpxk
GWuntAOK9JLzIuAkm0UMvn4bhXy4oVFz3eC0FXx+54VDQ/iUiUgt5QEwre8MRbYD
vAFlLSyPGbbq9kgBJUWC9I4Ae+xNEJNKlNbWWlF8S0jnqN05owB4gltNMih16HuI
jW/H6DFEJooX7gVKb2gdJHBdcDdmBVP218J1AFwnb69kV1SdnFtVWmQ+cgRbE6aP
q7UkkhtHOuaRdit3k3wXsGsUc1Vtz9BFVvZCmHIS0PrOeA75idC5+VGga+oS3uJB
/L6g+6JQ/HdqmgJVyGvNUlr50npHto0pAlmOGIAgXew4L9DF/S6BU7/gLa2Rf4xv
R5wK2Fy/LW7dFbZsY+UU9DO071tAoqAuw7zWzVWL09UcpZ18L2R096Y0yYOX3kTr
WPwcBLthTSlL/kQQRLOS5ZDEjbofSTP8nfdjmM4CXGVLHn2TN3r5Q1DscJ+dY/+G
8HDjPNlhIPVEv8Jybqw8YOqJSpYGqANwPVrlR9eoDqJBoT1mtLMT83Apxg62qMIp
M9h05M7Z6VwtpOd29p/xCeZs92+cNXMbXfafG2D63PUw79lYsfJb1F8o4tSSzJKC
GeaXdDN2fUzu8G6f4cZO4LYhOXorxTqpwvQC1yHXqH34TpKtjiH5XSzOUaMRLDen
n6BHsGV9f7vqj11d3TJiQNcHLKGLOCrKGycvUuGphscJXXMhyWs0Sk4IZBoHyFL7
5INeqsKgbPcSCKk9me9EKsVoxiYizBb6SsF5F/q1gsIhrbWEftvA2Ug99Pu4Fg3o
czGK8zTNRPjYFGvdwIQ81R0PCmzKnD/OupkkTuZfG0AQwzwshoH0YXcFkmmFCzec
lFKizVeeKcJHtbNIgDuT6k6CocUZ1jj+nZl7b3mu5rv70xmoILqREYAphnFt23Gd
2rA8n+LnJYNMCPlMNe8/s/HXTTzQ0IXKXGiGjiiACK4H4ZpMLMVSHwMtDkXUWmMj
hnsCch8LHvNfviJ8tlKb8QnW1UyoubYiaYIRs4lnO/DkPB+HhUZ8EbaeDc3qTCGg
QxxJlyUrlsYTwO5Y57a2y4wDCcFJObCvMRtIEWoA+KVD4LofYGd2Vj2oPRsGRZ+f
g98XpZZCU+KAEGX7Daur7tOZBBxAjKOW7mcvTcKqMPc7lWK86VfXVP6NR+4OuqWP
sEpA62svm/HmuErYaDzO2otfsVD8aOp1Dywk/aHKONtPEO1rBDZ9EOK871BhEZNo
N+FxdoMt0ztB/98cXxDDALIO+bTIAlxQBmLxbREfNDb6Hhkzuj2auPfc1EN132lJ
nad5oRw43yKW11YLOyxXLIiyJw2/FgqyckMgQIO2ny4qJdfaan+6qTSQg65xhRQG
Azy8uJZH5RzfsdUxJ6Fd7LnM54nvZ8fpjnUg1RfDD1NlxFU8J94Bl5jB+LfmdVZB
vZ4fvVugL1LwXj3Kt4XHDasrMXtnxBF5+uwNJYU3WCtU+s+GeRwTIF2olVaeLija
uS1ZrRSWICdbFFdp5ekOHB0gXPfkwO8lS1aO+JDbb/9yanlpBVksaixmdDdrKUmK
AIq1Ar7K6yqofq0/yDLtrj5WJ3FOKj0bksb9BYvBAlj6LL+og4zekF2Vj54tlWtx
6WUNtE0/ezSBV1JtOX0nBti4gp1oqf/FvZxptWmLAGMi35HSN3RED/BbgucLz4V/
75DBFZT8uGFEyIcLnJsMDgFQfFen9n6e3iZIl3teON+xWsPGKrVfW+Wl6zJUDYm+
WpvrWr1l8ZyoemSkTchuoaQBs+zMgjFjft51mV8jlnSq4Ceb8fcrwThGSD4qgc92
XzgNSc++PSZWZq/oi+MEzEaUFn5BiKY6LeVh7Dq1hGuuwWJzUuW6xOGwuWbXSlu8
Dk/kEatJTY71CP/gxlUnkdAAZaEnXgVZEyhLIxHcdkqn9eMRbRJQfUu+UaG0Ap8U
yYZ+z7mlMEpMdAijd69Qk/fNHNAKLCOWHCbsp/u5RqJmNlqGNR1hsCnlU+NwNMK0
55/EvRNll1Kz45VjP38MAwcTaB8uXDbTpQC/4iBlEVjQ+3OpgbtLHmDGC/Au2Nb7
2dNeWkTCcNh/GVrayYUrLAEN01dZYnpXRjtY25YYju2hyutXhvCDkoACXpqcbW95
R29BDTOE7rrDaeADb2eCNqRVAHN7xbPYVoKtXNgCxKE4rh/mvUesNBbMQl5Kmz7H
K9RvbEb86G1koixprhm6ubtWAYwA7BngelYNU0gxXLFiv1aWjLNRC+b3hLxOgXOE
Jhmu04WTvwu4ovzTRMQlX/Ly33cmMnSQhcpZ4VOOWf9E/DGUFA/tiX/PaJusLahS
EZI5fVYGvaSgE/pGTJfYFzEV+LAFKbAacfEqQPgdu1n2oE8W9E9zc1F7SVzboFw+
gxahFnaO5Fgr3C3kYkRY90Z82T/R+DNxmXjIuQBxcXFdDhHu2v0u2mMyVkE5ANPU
j4PeFmbokROLYr9FthnOBalMzFiUzMRhqGr+5mEqa/lw5Jyc2/nUXyWfTDLKWZSn
9ObpeLxMpivkMQsK02bQz7GI6aef4HQq5cxIqW8RuArXZzkkoPfcsnJbLvpTRQ8C
7VopV4A2imbYDn0bZCmXrlH71eqjwDFZ1X0gVA1/xazZU5A8+NZNoLn3MgUst0NT
hGR6K3KPmxqnLpIPJppmSc/AyRr2Pzaw+oqeZCYp2sLpINRUa/X6fZv+uZ88ysti
BMAB2xhWkPb8ugyQPkRkgcDg31pQn5mrfFFgM8iyLtaoGQrethp0CVYtb+ffxxFp
dlpOUrRxG+5qwZ1i8IZsmqLx4YCwnqGOWDhPmhci8RpFiFz6kK8YzFltCWV80aMk
i+VSJkYRVcXlyiTZd3lWWWhQLYMOC2WIwqH4OrZblvVMJNXTJL6WuFRyr/n3SS/a
rhT7ZbmCl20IVZcHbr2uJarIHDhwAuO9qZhdcO0C2gLEoFuxkoEjxUbf6j3sBz5O
uyAAnZBICoYGpsMr7N8Fwo7yInisMMVKuQvjo7NtabVGfWu2dKqpQcEdkAwRp4d3
j6MuxFnPfEEOuD2NHjWBXWbJaQgTv/yfdrO8B/5+eaoscw7vubUpJehIA3Rcw5Zo
aXQ8zjgcL0jM0abTirIkF1Hde8B4MpCP/uJ2aBYXAVpKFY2pZ6L/jzmB0N5yBm80
sCBuocP4pqX3jX31gwrDrHrwPEE7xnpUq9pUSa8/gKjtjKz5siX51EFirecceqvN
3ALum86ldGu3EZGU2XvVYY8AHjd8vapmZMZ+AnsDcsgxiKmCzekLznosQBmnbG7D
usoiXEAGRGnsZ+Mwi+B54IvPp1YMm+XtWBET9DEhDtJezgb8I0f/doqzrJAW877T
dFgrJrgKAlojXAcKoxu0lLAfkvxzp9uYsTKpwjkKP5kFN00XKqpWMjaVg9HL+Dx7
WnyqI+Jks6eFWzV/ngSvcLOb5pV3qNuWTUBeq2g+i2hxiluum3joXnwVGKC5V/Zb
aBYcdLfZ8o2ctDFkacnRFhWDFfWGudldBTezpXUgm1ZXD5DRwHSAUFsIMgXcZrjC
hRG19Z9R9Ws2tuh2MNfQIrKjuWX0wIk7lBv2h+aJdRh94T22B282CxdKfjGiNqf+
gSvTDh95M/7RLx54DNwXdGiJggwhJV4xPv/KQTVPnrQ3HCVUXi1k8Q8XTfcZxgxH
nXV1MRHabBWnKiiVmyx05zbNgVLwNcBENQoShYeJPI4nJNsyRc29lB1ZhNbsUN0I
2ZNVxuX59jVWcF8+szr31ZnV8AzqXSpQfEpnSzCitXfiXb4XbzOKdLqGuXd6vvi7
ABts9k2OhKjsR8x09AsH4ityAeGQJNylunuSmR/DK6G51hb2e+ydoLCmAwgLoDb2
5mo153pADRQvdtrxJFOF4GXvuRJoz8Pm0tUl5mho/t8nsZnKMFfohGBYkAoYS/EX
Kif8L2uMu9qE+T6/AYi2kGE8mn3uEZCcYeu1YpJZ8ucqXPBOjfEw4TpXAphh6eyj
8LYSNWHuXrOjV2E239p5NBQRAJFQJa3Z8Tqg2Eocfh+UEFQ+5qd84laKyl/ukElU
Jz3iVtiJVvhGVRgMmsxUvfvXbdCeMs1mVvuvNDQ98+zQvGXuZ7NEnic+8fpFWfOo
YiRBdQfTz/Yc1DbbMtAuErAQUk7pKTWr1ffDMOIcUb4FjkuLN11MolQDGHmvrYv6
W/JUnFj0yrlWThpQDMgLgBHpvcXEmVy9nEwJ5pQ0NKyttQ4VglaoY3SwCbHyi0Yj
0Na1Ay7+6KDOfJlesa96722uggpNju5THwuMH4Jx9w0HpjwF1UyXck/gceHE2aV+
eYKzI7L8lF62Jr2Q0z/gv7nbnuuoO+72jl+WHqPDgl7GOA6LACWjzSQF+34D/hdy
ZlJ5ChJHprCtTDDEKcfskxvuW54YTm1wdRGcN45xMkgpzqO7L86vGQ1FI0MRaNIV
apYiysMvhS5YgB9FyyFnQ4oxGyewL11lS0RShUDvrnERtnDwQRuZ2v37i7DFqp6b
jUER+FncCGQ8p2tgJUhrdAReNovQDa0ELPoYuyBzW3RfSqySLNCFQ3AFy9QqR5Pp
LWzg6Pu/DES+peedbokjm2XhKIaHEPJmE3v/gtX6eO/Rv7jG9W4HLxrPFtaG+fSS
UofVzhwjHvrPIhJueA2Is2lkvCC29aDBskeMKMFQl6NBaEi5bHsBUEeXIqoPZpfs
eGBAyIWvgCAmOVNU6W28+tQ4sQm8UL0r8WGNHeZjvKKmVj7iwqFHNpONhwtqmM3i
E+3SJgFjezax0xTuU/xGRYlvv/QWfBRuKBadA/DvGvoGKnRyoLlVmSBodpKkycLG
pdcBUjX7WVEn/n6sNCA7u58b+0GR3DNKlhMeA/JS+FMkT+wyIUL5gqfQWGQSG9oy
CdyKThBF1WfzK9jpIQ8tI3vWIhwKA5BxpvksOw3YTYdB3s3QomZP460vQCnGG1Hr
a1ExJWES4OYKYR71sEbWQqMkG1HMdtORRyd/1n76xr0+8MDg03ES7c6I9JLED68f
FG6FwebpZSmfExc3F9blLBSqJpACffM8NQkpnOXinv7Jl2Yhc0G535qJeTuCWduV
z3tr0Gt/JbzG8WYsrXd+W/fokt3uL/1VzLv5TazhblFL+7HY2fsoGL/gWH9TGHVk
uRdIPmOz+nzHuKICFqf300qLq9mkAryCvf/dFdh/G2RU+vsDJxJcHGskhbB47W3h
m7+XxwhN8CVe7hG7VAg99F39Eq63vWofJq/7qH4GZUQXQJEceQ3rHTkDzBwQ2DVe
bpk2EJ7lsrNEUuB/28IwgJfCj/WFAhKu4rA/bRBffGA7kT2Uu+V6xAXexZuxERMD
Jl+snQ53tuijw4z69VThZHGcBOmdp0mRN+PZpohwGhJRk6fnYwR4l34M1vXzh/4U
wiCwaVCBYMT8fbIYdJlwhqnkB86g/Gxw6FRYsl68QV1OcbcsbY2UVkFVePVpNTJX
BodgDO0ri893uQPnY8eWsYjalSKvxsEbxYv/RI0aHmcPEs66bdE+kChwrzQjAomA
IajErDa6PfMmTO7+43EQQiSutnrjL8Cw9CpqKjF+RfDwetvj7MACyqzoZX92UjRo
cdU6mb1cfnrDHtHSX9VaXDHRceKs42IobSjpkzCljL6t9l+6DdgM8DIf7hWx/BqF
KY0IJLTcwNA1ns9HDk46cu+jOqRVOrGKteFd4K4PDJSCMaIXLwyr21Vnkm4o4j4Q
ewCxfkcp4/fVSfp9QoVndmydH7FsKOkboYJdEhNvUNXN4vteM8MK8jLu/qW8kXFN
Rb9Isebhx+yV8STl5ELN7dbh8DcKaGmnn4Sb6MkPaiTNiVO3wiQ6yoabI3breJ0D
PQWWW/Apm0Mpp7JRZsTtCzfpW76c1qzOLM2fb7FDwIEIlQJFejFO3T032U0sXw1e
Ur6rcxLunNrz59DMS32VOez7+SnYy2RRaQ5fsJwOjniYFv7kwUJ7Ph4iv+yCtJ7P
Vc5I0170YRuuXsg0Z6RFqPncrYZfGxs1dTa7LuaRv9ZpZEw/sI/R38x+Mxrizv3X
CoY0oUWwAD8lyQhBMBisLl2m6AsRo/TX3eOkER1YZu5siZA+dPfb398ROWLe56jx
f3SGhS3KnvmAs8pt6UdXQkutp73GiJmddV+WmGTLlEeHcUavRQo784fFQuE3aQ+d
yTdFGBDneIeKEUka5POVSLpc8d13m294dvG4GrMRpm6oivvRj444q/Z9einel/Xz
mVWuGn3eHrsD4dXWB5Z0AdpO2YCA/jh4FhP0XtQe7Bsso8UxcNObuW80hrbrMkuR
82jc5EYh76N/Nd+a/gWAFyvEsIJn2mVqsxyIBRKX5CtCE3htt/8gOa1sO4X6gBc9
2/OkFxwd0kAQ5BG3zcJSlh2XUFNP58b8ei/zgMU6p7xWRfg/KJ7WRtYED+sjkRZx
8O0a0gYzokq1GL8OTkv9PdAJWtKlxSc6HleUeWvgeNk+jFNfJ/98174YgB78Iu4a
Z73iMQIWWWP9uKSZ7N4oOM1cgvFi0Hva7ZpMvSzxauVRsemQkLv2U2BmIS8to3L/
qZjJEYnTl4e3by/2mFTAADE7GtKn+7Uq6v4/uJDrispy03m6CZ7r96EnttfIT+vX
U342EACogHA35D7NueXKOMCr5lnRIZ2WPu/nArZJSX3OLy8/mDKM5cx0gtdigaRf
9zQioU3gywEwVgBRBZTG1B6pwMXuqvyGRiOVap2n1KONGV+Q5GHZNHIx2/8288Fm
20zl8GVQ3JqcrVxumhnAFxZSJp85mAoIhM0hNTfnzDfjdvLropdka/pb4vTlQhYp
xrqj1cR1XYP4xm1YMBN5jVelg5imnfaQBtqfOL61wcPPYa8EeQOQLKXAmP6zviFx
Z7Y83U5nSZNeNpLbf2ciZ+GxLm2C1ej1wZVcRHe00adYp4CDosLEUrN8lWHMhEwu
T+sVshlwZ7vpCjlXXt9i9zAH8foTAhv4eN819D6uyU0L6KK7tuyVjfbH3Clxghao
qMCNKAPUY7BE9PsL3vG4/1GB2FCq91DwgVjqaWhp4WtPfkHdNLyIivMqzE3+YgCA
RBbwf+VEUvuamQosM7IvLmIg7mNYnDDu+BYftJZ0v97FpcIiLMUVTT5Uh7i+x5Qw
fG4NBE+kBFw8t5jp/6hLwCNf/xlTe2uqYVvBfXsepf0IHvaeRex/WPhm5vJTiiFY
LhssWCjP095T0SS3DmkCBYUeOPJf0YbN5ywb2PNvIl0Kz88vLt8Gl70XZ7bGemA5
Jk/hptJe36/csmk8ZeeMSMMcBLiFpfS5zalzG6C17Pfks39tjpZ8hONNDGw/wK3k
nVSQs2NEEEZzW26kTxoVT2HXAB1OZil5VBI3A2aoTPy1qXB46f4D4jIQvY33JzJl
7t2bhcSQt2yq9RtDg1ZaSX4/x2ERskWy5ZAkGP9AkrE5AGm3otBXhrwsR+kRypWw
oIFohBCN7lIrWWP/s4WWWeHqON1Wunc5wIt6fJTp6T7xUMItJTbMYbJviDAPLn5X
2fk6SmpYcEfNpP6T2D5la6GqJfW5jUcIzx6lxKWhHyUDbVkSZDYMKo7iytXzH0xi
PjvbKTJnR6+j/ePGm9XxwWlfOtVqbyuXCzGsEVNerthPecrHurPHMJAHRpn2WJLp
hkvsO+js4IpXuuE0w/RNOwchd58C6mFIPtrG+sa9z96DdN5ve+RnMewtjG6nzRyI
gldnSl+FZSo7hhkh1PzRn9Zp9KAEw2lfQQlVubfsPZnGDAJWASFwUw0HxquzF9fQ
TEi1aK1hDceaSyi6qbx5MFivzACsvVfKFLOFJLm1w8yTFqlTzhI+khaYaLhKJNcc
1BsZyty8wPN3gSAMEgXfL57Z3tK7uVEvhtRv4GQ8W6G0WMv72I4vAt9czQ6U5cC0
EakKai34k7yRFHFpvV/rxNkUyTBJosS3uBPQXyz98lK/J6GqDthmokIdyh2Jy8U3
WloujRUero2hXwXb8f0yckjuufnYPzSsZ+1MU533uO/qaEVC7BGnGXqZoF3Oo75x
OwcCGcSUhysPpszyCUXhrdYGn+rfj9z03eg5eoV5GZB48gP8dOh90k6xWgT34bl+
zk3orn93Xx23DuoPAuScUOfgh9GNoKy3MlJUdhfECfg33bVGzX741vpS+cOlTJ2V
B1/qEZmTaHCXClzAKyw16GM1MigZO+M8hjSWSmxzHJWOXkJWoGs7x6SBsCQNICAc
/o2VZaRJmQMex23He+1KnXPySJ/mfbzbJ3qY3Jf6tfAz3v3FqH3hfKVgzBFZQuX0
bu7R12A42XwfbOwxKtPTHbGpcz6XHEA1mz7IbtPOKX56vFMcyMw93mI2oPETer5k
jMB42O9VZqyE7EJ4t2d5YTpI6PEkv8NZeLDn3+f3S2ZzY0i31IPvTRyhIZAp1+Is
OMwtvNGO3Y3TouZUWsqiS8DFpt5qf8oWdXRupt4T96gGYRFDjQoTRN/wONx3aF3j
LRoPNlyf3jvox7YJOI/uzHNpf1BNBgqSbvCmuIkxaQu2UYzT4kIYo24azuE0VCHp
cXIPf12o/AjsCrvxiuFduus/rbgvlPeRdrmh5Jix2DexCYajQPHH8JpyoEjLBkvK
uwUypyFQ5+n6egJXmL3MgZ63LWRoTfWzDrwEnDhem3d2uU+NgrD3sBDq1aFpG9S6
liaiDmybd8OnqE+5L8syL2w5gEp+z2CAsrRYWNx3lncDqUQSXOA3153Nnb7qH4dO
14b6cQ6MHVJCZsH1bnpSowTfqdwSVFaK+oegTRxPmVXoGkqoXEzWu5pO7+KqZrBz
yb/wHsQ7bvrpxIV2myZmn8EthL5vFpo2UBauZUwq7GwQaQwfv1XhJ4f0WHtwbyuo
mZ2XSwj84bl9DGkFCrvD9TSr+HVGbJpI/K5OmTRpLI9TvcFi5AfgPoi9mNYCPMpc
DMZoKUb6cEA1XARPCrUL6kRYm4epnPY33Gjp6YaWbleyEQUQZM+ymQrxiFr0IlwS
Q4xrCDnQtBekSgAB3PNZYO60JTPKzZoPbtPVTZxBD+zeG1JUy40EbTyfhqUP0Jh1
EqP0ipRjECZMsGsr0fnvzVP2HF+P5vKWnLm1+3Ghxhc7lkgQTz5IJaXv3IzqkyV6
ysLn7V4DJZCXpoUXILluDPkKNNP1dLOQLsJmQKXxYi91IWc9DdvVt1HTUpTugC3B
YF64ZY198dJTOTALrS5G5e9ZIS3jQa9OIyzg6bbCujQYsAO4kivZ0b6BFzwREdBl
ugMpvjIXQcyQkphJPiVGnEJq+wk9NxmmVlTXrSXvDzZ4SWCyinlSe3TbWTnK7r9z
C9jzqdiXm6lIRpzhKNIKT6hj+WhaZkLXkWKOHWBve15mJNVpHcKXw0DbdkE7HegB
/qulyU/o72eoOx7sf6PIr0qunqD4eyuXYysgDMhM2IR3Z4iFunhmUuw/fbigUjku
FkwHJd2tpWnJIwJrIQNSOKrofrABH1Q1zkQS1gcOWKKaYDhuhY147RlpyPAyUU+O
d/umkiF3qU2+RMsnySz9mmqrSHLYjMYh9ov5PINGGSiIdw+RKKeJdpM5A9VOOJ5V
d0OrWz2mi3aYXzd55MTXLbVh1gHGvY3fZu2F0vdSTVc+pD3tBlgIkLnUylAAiDX0
d9bEOosmsCjTbOREvelgGmicAcHvTbXN3BIva5eWehocHBW4rgQ5T4BwjWvytSHf
bXDTRQZ/oSuGSV1W/dEk0vGR0LG6gMtHOvKQzJqBhMBe97yOHYHE34Kfy/u7IrQR
0jVtOuRTRc8OEwLkyo1bzmRTRHcab9IetuMozwADpXTjWKIuD/IVNCdil/n1hfWW
aXeLmtsfQyr46hW1NHv1GGpo+zIvRI3EID6bRZ7RSpRH2VJxiaWLjkXOiwxY53M/
dYG05Fcj6tfDzg8NkHy/1EBjIUhHpinsk/LcfW38bSXUVjUHdH6tz/Nzk9WOocdc
9t3qsYSVRf5Zdxkdoa2bxTmK+1afDLZNcb0GRlmm67b5Gj3Ag7wjOIQ42MpjgVRu
rU9j1CAKNJ6et/qGSgljCtaI66WFAlSzrHQHUBkvUCoyDawUsGdYoH9amL0pyHEW
auPP5Oe1KysKwLiZLdHXDcT0pptvx8+SgMRR/V6AqPGYdVFTnU6wPDnKpa6CQYdd
6UfmDpq0+SO0tHDJoZbEPqJvKcd/o6iMrI6cTP+Amd2t0OGHdo+cvKDYMI+FDCS0
7nhR3IpIhz5AqB8FJi+XtAoFDfQXf4+Dmwcy5yM5ZfHsbSBQ5it56n8Gsz1oRIT2
AtOYm2sG3uzI256PAHKr6ChKpgiVfwKPOz5sAKoJLCyH9aFOVfcptX3KOYGw2vFu
T5bUHcp8ifALm1hGGAeE6wnVihA4QcouCYvDaa0P96AKWq/TgAGlmhcVBZmOUTYR
UT5EcTa9IisPwkYhMCYsbS2Ztp7+n3g4dc7pTX+ZbllqaNajpGLi7UPMQj8l7RER
t1KCmx30nbEIqRNLF2iylTJ9AR6zwPOPlTIBAI8MKjBUVkn8FXvNHi9VQy3QOA9q
8gzY+ton635o11d3uMYMdJySjlKhzjUEFoqUfF7RYDrTR3QDN9LK4VmJo4yCspyK
NcWxXvwvPPHRn1sWuxo5yNsjRStUwMAkes6lSMk16EP9aQD41Kd2dueR291rrTlg
WMloHIn3Yy3oU2s8vzmLoGZ/OZSTbTYqobhZsDD1HpFLqzjs88hiRtPUy0fcfAdS
NJSilLSG1jyxsnM8rcBmTT4klxXSN0sqOyWBWRRxl7mplxXEzKOey2URldFgF0jx
PnW4t3PB0s8EYhYYwE42Vas5+CcmjFxO0fHL4jPFYGqqbyYQVq4PJ4uN6Lrs0lVo
EArEJ6ZOUY3Ov4X2xDkwwc6LFtHf6A4e1Bu7Z0mbKRf9UKOtL6G2PUMXORM3e5VB
lwG7tod4Je6vTTx2liz+tjxJd+kitPKAsAaNT15nnuNVZWcmtTldA/f6og2EAyPA
Puih2hRYGZReYzL8FKYUKrNG2ANBUc+KEKq0bdy9kQQvKkiXfmtP2a85I79lE3EM
ZoeSB0P24VhQZ/Y1YQC+LGEpg8CzL3tqpQva3pRFCjh5PHUZRGPoVh0KcPJWhKb1
PbKPrys++to5YJxhmICzlFPkbNAe0Y0YY6I/yfTKXRdU0ibr89rA8TyOLfrOzpH4
AI8Plfb26gi5Nn6nSB2R0irMT84Qg1pd2H6rnyPA5ca0bAJw6cSLsewluhb7RcBH
XPAyl1KyKGiK/QQfTZEyGGW/z6KcSE+DJrfCeTqKftQz0dhackH86/Zeh4SoeH5Z
IpI/8DfKDMl1RS3INQXT+2UgBXjmJ18Iet9h0c6BPCj5eIqgp3HmrD4DqPegqx7B
LjZG26We/47hgG+FPGPjrEcyX2W6dWoIM9kDbehM/f1czN3JpSLv9x2acc3S/Q3l
WFkxESh3ZOW8AmYLIIN9OXBnSdHoINOuyP+y2UG/vXvNTiI25g4zVEfX3vRCOTml
PHt8NIArlFLgMtfOl0R9cXujQEYrpzoZb5BySdjetBT4gOdlYCJ37Vj0KyuJ/zzZ
HrpAWAL95BRhgXzhpqs3OOl3MlLsGQkMcHmHg21BN72I/z074QLY37Czzxiyvuaw
64Fyql96isXTd1hIlvsP2viMvLkSqtsi8UwRBbkKD0iUDj72BSZubPw34rF3V8FO
C5zyvL9qq9ps8+tQRbmMrOns/623rWT3meHA3uSPd9txLmGhRrQqYSeDv4EO606Y
Nb7wIGjWrP6k7JJKFsu+Kh9bGsMPbIsH0qzOjrc4ECsrdWPzX57/27rTki9y0mJH
ichzDKJKVugavvmHMLqVaAZUHTjx3PwsXj3JaMTXo3j80lbUd5CHAYlY/X7gPt6z
Bp7ZIg29jj3E8f/JLRf4pMzh6QCm1j2fZq9QcEXuJj0EK5v8dve3zJlvhkGT+x13
CzNbogdIhIOPq4hpeImOpHXdW+ZnkhmZiKk29EQd31D0JTRCc9PY0tHxqOJRliPZ
Bbi5hn41/P5NX3id3Hp292qAHqABCVYLa2re5BI6gdVZfP0JUT7Bth4xylzVo27h
pNrZoGIAsXy/AEBX8CUri+6DfTJlNYC8xD82vILprnYS2zTkb2AlxT7otHK/+VnR
5kdH/AxkecKZ3ZpvHRVSMG8N6SfGmvgflW8WWy748CIts3bPBb2IteZG5UZbwYIN
DrmOtVCm8AVZFYFJmoethFKlNplITOjx1fmZ1pOR9gv+qdkCm0rd0PNpN7MILkkn
f+DuEmhdwUcGADdfo0cPDzOaTbw+alLrjTpoevFf2gYm0lcpqEJEO3VZ5Osv+iP3
PbCmVWQsMylIZg0TVu9jB3jXL0jnampFJp0Dtjlj2MITirBIXTiYd7k/7e4hljM0
RtlQCAdq/0IeCp/LdfsFaIrvjrwUaNsdkuOKqzWv4/NNWwcUd+jr9Tjg9un9U5Qt
m9CNzbfDEN7h7SAxTNo5+QJhJhjy3cRdFuzjPAH8M15r6lxhJ85E9VRqO0MwH7x1
cGZ1wjF7V7zeIoIQnYbquYxmoUWrPPhwIUoWBU0nc5PMf/dDzwHNWdKbpFhJ2S0l
I9lGXmsIzkJaASqsJRb7/cd/iy/fjEJlJx81EISj3d+BnWDAulJR2z75lpJHmBwm
xxvsVKkIqSwQdM2TnIr+vVmDRU40I4kbLjX4gLJ5SviFDO3h0kNXgUwcrSbm2pp/
qjvJPuAuPZc5a9jjp7Xn1kEp4xc6UEwTErn4nhdedQut27lXHHzl8EtWAu3wqKcD
BN8jvVwP3B9f4bXk1mJduPWFSpSSXLwf+Xg9uFFJi18vnygyDcKbFQWabk51VqM2
RC5JJy89kswuwDbBKz/8HR+XfWV93iaiVfEnWbmVTq2DPy6FHuFOPc5MBMQ8FH5j
ok6XLs9k497lv9GI9rylaqA6y9N+aFVwhKFDKJzT/J9A+4Zyk4qssjRrXltMizg7
aQ58Rya17RQfHafR5+ATbkWkawaIdY/dtMqIIOMuf2p8MmPLsMo4FBgH0JAAZoAf
g63Hy1DRrrRodPNMCdSOkXSDP/kJUNeMs3gmQP5MNH0RqNVbMuJheKJAnJKzeHFk
oUSaToWb0NDW12FXnIXs8Nyv+PrWU2SfXkggB93HUOcJ/e5J1zsF+lGlJvWWDRmo
G+aAHhkMl33GR7ZZIwuPL+5iMg/I9gyLudd9MUbze2qXxTQ0yHclgt1hkRyeXWCE
ucAx7Biny4Zc5GpGu+Zj1HYMkneqspsx8+HJ7kNGZAfKU3XjllUf19kju62Epo+B
FwjmDW+jiweZRgTTkGQ92sdUfyvMpG+NUF29euHyCWzD8PVOY5Vbs2sHVWhOVNTu
cZ7i7PVF0AHtC42xK4r9oWFEO7/0UzjTphLkM3cAz3NgLI/d7R+u3asRPvcuy+bS
+Uv4jkYiIicg1gy6N6mwlGZMQFlz0BhnCIQ/teEr61mb6MS1amO3X6uNOmLez0W2
u/RckRCsCCUYuAWJyXnOFJDb8hQUodsrQRqld1eAoNIxVxuMzJyAfAO9v0IE87Nl
rwwcW79ki1jRxqz97wL7A4VZuTxdhpVIAki5GwYN0U+EL2dmboBBn5ZIDwXqTziW
kVPr/wXEWCsnPCbQgW8sLHHhjihV0olCLNUkuKmsv4hPljXqxeA07xRAbmRUUww4
jY4bDYo6LKMjeAFV1TbXkjDzsLB2hpAsGzcV4dZLx7LPj9eTfIiqOC8JJSS9Cpg2
q/Wp0D9+Ntw9l/4dGVM3SHhsJikDmCLSvYXEOavfVHOcKYBus4gOjJ0Lfjd6LfLi
6AxOr1hPlUq9A9UODOfOHYIubNM9rT33htw/U1FP8lToSQ+GEd3NkN2d1eC7ykRq
cc6MP6j5MhucZqJ/EgfwRO5CxeWyJHtcV1HJRD6rx9JZlVQLm2wITGVCj+cA2B2z
kaILD6ZCkgMF+ogJx6IJXqg4dpaQoEIAH3vmPV7jpqkSiOttr4yA79DmkJFMXXT8
dqyiHIlq9VXy8TyI+1/Ee50B9LJZHkTFo94luXKuOKF6Grck+InSa0PAbn6oX8jM
/xsKNSfkDdjKsEfsTVyqvrd+cSsETD1RLupfEPw09exZYYpejQw5eOOvsemmzqIT
fbXlBfJPbtS0JA099qBEctnnBARt6Bjxf5Clcd0Ryc3846gCC7u3CqiamnY1ZWAk
xsuS6Ic1lF7LUkZT8DLJB+GtN1qKlsrgE2BNxolmcdThe4r7tRnfEIWEuIuuGWZ/
9HPoYiVdEFUnQ5Ix1OtMDrcMESKu8wfJall6c4M5ldQK6j35d4s6Bpvw8zfcWlzs
EWNcc47X0nJPQqHEGANTjwncWN9YOyaFYJcJ3gR7C2JG+F0gfe5/57qYaWc+/DLd
EKauMR2Jvh49WK0jWeBI37MAxOPE96nNMj1SQrk7vAVm610YWNA7kqDQx3QrLVaK
jHkCuBkCWupIMldaZLPWVMFnoz7RmHEb+JJHT4yZFVHOqVpRF994On03WEMbaIh0
N1DhUXGDL1wyGGGO5+F/L4Gq/7ERajSi0p/RgsIC25hBTN6jUf+73CHjmRi6+vbD
snNPmPq1hyot+B8N/CzwDohCOwJz2pYSX3eIXOupcPTfhN71rZYCdhBSMhU3y68K
BxDrP3N1vYCJLdfcI1t4c15L7Jo93FohjTx4x6hWUbUJFpDPRiIlOcZHktthaUEE
qxaMVZLsfT2yO/rDZWE0/txK1PCrW1NI8ZehFx60/REmwbNX6/04UCoQabmwE7Sq
Mito2n3u7VE3k8nPmfGbV2BmQw4yoqRQhlZp70cQDfFnqdD0WvD+KWjwya0xjld4
Bvd0Ttt4e/S9EsPvY+EBUnEx9tuk5wawrbIkRDhDi+VcmWhnIHmAZLKhJ+m/tZ7t
c0aV3l76mxSoSpNWHWF6vmC1aeBUW6G97DD4ZLh6Pv6yqYHm1qaNCsr5R2APF9lQ
A8h9gR37a0aTo5sNRopPXNS26FSgso2MdjR4H1ANCJylwuDh36kFGbk8OsB810Nh
EiedeljgzVHEa2ZcraUlcb0Ve6pcrAJBU1fC1epGw4G7MchFgyovT65md3bPSmCE
6egkSLygwVdNEvCGTMlmSHaZ7M4+9AFxMjP8EMZnkOfeZzGNroPjsDViiKZKjb12
wfPHM5AlQpCHzZPX7dP19dJG1Z8YV5SJTRnKhgOyWC+5DHwPBXjOflpNNzB6Qfqw
yG1RwYPnsJdHkm1D9OxhugbnOJMB2Q0jIgIbJCYf1nLDGgeWk0Uj4dAedTbbbpFH
95FgMBY0xI51+vw4TwZ70pCq99w1GdeSejR5M+7qxEqejVBxP02i6u/MxKVoXpMc
Wq52R2DFR3haT23lgcL89gU/HIMdz0AWVgq97M+uMFSrksD6UJ3/ulBVpGYtpvP1
pekHhp2azuVJYU+UWcsldQDXdldXcaypJ8wXzXxg0jWUSzV8/wm2DQnl6BaJTp+M
SAjuSYyVt4O7aP7A97h0GgoMDwh1vxAF4AIkFvcPfonBtE0gbjGzOR/6jRZmInu8
OIWdPMMLJ9DKk+l7efOFoEmbK+7Ov+I+U9bdGA7lRwbt+5yJq1QtgPwdjqTW2QMk
baCliy1r3bspDhkapwBtPMWveAFCQFLM3SLHdVk51iAaqFsn7agEwOBtjREqxVEF
qyXnlZJL3iN5PB857Fe6IAP+KsYVeLjojzPf9Hy3sJy0BTwO0/5qicFGhFB4MdWy
MrFIXB7PRbSEhhiBx6sx7aaEiXeE4tK19JMTQTbrUwSpGtFeIeF9XI3mRemOfBs/
IctVHIaJb8a92yjP7dutBnUjSWePufIE7LxFFBnlzR5KqFZuXUqgHLyZrMRmbX64
uDNQkWM+KHEjRpUIeamNmrJHdfwkVEWAYl+G5y60EiujwdajP+ZoVXdON0r+bNBO
+pHgqoOm0zE7+MwSHS4f4m4NyH4CG8S9WLiFffPzwvbYLnXQpJN84ux3pPjvbT7o
fq9UfPgICxUIZwZ7BdFL5IZaC+CGWHueb8szkXgl4KKKSYCtGPIke06swpm6dcV8
vI20fydxrwGajOIfWzQb50hVrKcqXQTffQMhtOHGKooU62XOmC3WIBL+IWuSJBXB
CG0qqGcn4KjkGdP0gKEO9p0bAB9SOsRWACrjiBuC7N8z4bAfQd3UDV1mQPhkoz8i
Loy+K8qAmKwh4OpY4xfcSfeZXsZQD1f5sXp3eDpLg1R0ketzLqX7vZ2eoK+bkyfU
uuBHXwC9+hk97jwK+SlyA6Y0nTLIwwFgtbEymobEa4umtDJF+Cl115v/ZTTbshys
GlN8YlFVl2c2KEUDnpECyADHdgTA8c+35xOJFONMXLjWgN7UNwIju5POw0tcheK1
8AWDF9udKt7TEU7z9SJsxEqGS6pUtgx6O5kxhBVXyvK4nhJXd1jFs5WQ/VetCMO7
coqh5siqBKp6aAeIZ4Rg+yztObOPUbFp78HE6fhzRm7jFTM+zNbb4qoFMrr+zcSC
kuWiQke21tlBYUQ1QBaqShjcpU3BUw7c82Xm7n1sH3Mp1Chk7/Ck8FcKUJY10rbu
sS41aP6ZB6kYHxeTRL/OxmjhQfaTSypmk8CjSBljJwsQ15ihoeJDraKf+/iqdu7m
WP3a+uIunEmMf14LKIVJBKI2jqAh+20aYXGx9FIhmlYBn7wd+UwPyHv8nu95uAS3
QpH1nF2xJUMlR9gU5jvGiL/S/6iEg32Tb/LPXIa7Yp8sLNRMr0agLfdC+g1RTASS
EDx8OfO08kpb0mVNHDOtIMdCYWIVplgyR6QimPIc/n6fuQQhc6p77eMsa8vR5JNf
a6vHNB4dGKT9LRApqm9/PgyYzfVofxEo7poXHHWXMw/Qb8U/Z1HalqI06GGO9sqa
xKnWhgQVhHcTI2nARpSZMd5b1f+TUneuHv2TRKOlaNH3p2VxaVXu41X6xdPbISFU
GLVYvtdKcqAgHUDzWJFUN0jW5l7YywKuxDq/PmihSxeSDMHKDaTJ3uoWp7U7zqPB
Oq9WOm2QxAgYtU0+HYkn2uY+s9FDJAjgq8/NsGAFurVJk1LQorvVooQMP79FEUjR
72TQsacLCmwES99Z/m9fZ2K95FQKPhZmXiq4OvKHBwThZmYVY85glYH0O2xdm50q
AQjXzUsIhFviqscJINATGwn9/fpwxINHNFzl60ve5LSGUSF9u8xng8d7sCTH+UEz
lyyXalaq378Dl46KeJkeKtCerS4Lrgy7DfyhDohI5K9FWrzS3qIL2u4SHOS0mB2K
LOGtSCtVGUYSOH/YwmYvXxkHfETGiJmbbOP2mYj3TZgT4IVNvBMi2s5B9kyBpRhp
460mB9U4LwnFgBH3GvrIeVZQQ8r2B8Bdsh3vFMdJeB34qDqGQWEYqkIffbssGVZl
lijmbpSZX3TAtyhRSAimr4VwU6RKgZu7eav9f7cLXF5BAfel0wUYDCpOHF8LRXjK
Lldnq58BzoxstRopbEvOr/G/P6BH4LqpbcKbIXsrvfK3mNKgw7chK+Lrw8UQG7TA
3KPj489mnxohoFJft5iVkXN2ykQSHvPoMWISUE3CsBqrMuF6qTMMzx44Zwep8XbP
QEgdhA6+Fn6HKGqwkliqnmRFOBoAon+zyNP7sNq8RzSUpDvskxuGcSt/FHIJrjPf
+NI2FEZ++FHrXBYTYWTEhG5b8HqlZRsREelfe6Cq3ta9if8pP0LzNZpyE+MAUkyk
I+WesXUfo+WrfQ6/bHzM9MMCBlkhnwcnY8XleAVP6CYYeqR9i4r9V7Rb9tAeFpQd
18P31ppAlafnF46OgeUHknLrNLWp8lDqbKOO8nnTfv0WAmiCIx7eX0fqQff+/3bi
CfFO3KOdBtIkA1QxarV7v3/vnBhaicXfNV8KnSZNSe/ARCizrqRTGLpYW+z6t79+
+a8ixQRE3VndivamklxxnXqhAtm+thSSGpzNCNuUYb9vz7Es7llNq9LFP0+qr6ge
s8gRycVhtb2nY445NWG5UBbWX4vxKQz1mdFl8yJ8VP0pVF/TWGwHWFXY5EXxtBUN
wdtAuFeDOsKDxfWhnCT0zg+bNYTgsCmIdCWnKbh3LRJIH3Vi1h9oWxeqbt2XIjPj
lq114kyqu9qPzxdttR6IvgQrveotXtzmcdMeqrlhzyM8UkmnIwl4ZchsT6Gw3hBo
JR5LxPu5XQWNqnk90SZlX4mNQ3GACH47jmbOVnkh4Y57nIkG/QAzHZq4PPB0d6WB
9Q/Md6+TNE0d8Bgj1t5kBOllXet/txAY4KffbJFnPLgva6mVcLkHCOBSAyEE4mlB
LJ1Gq/I4VsPovC+zllAkZZlG6crgFuH1xeUkxwLtVdlitbmTfq33m8q7Ss6KR/zK
m/VMWANoG2RdhPoE077/fBLzfVGYVHS+oprsLORI4M05ncJMj1KMaBDNS2LVsaID
zPe7epnjKAv0b9YdiuUdmJAlGjIVVZ7II+7ReSViNzpKq3rwbrkyX2Qpir7Z8u5N
QkAMmGLYAvDeIijGBj/xqf731Tb5FDcskmSZwrLLpvyHJPulmqZb/z7HQrmkpmqE
H1+BgLDgKSgrKu1c3T9SzZM0LfDiv8evC/i+oVgSRwPrC9pSYCFP3n1t/Fr3Ni7u
bo32ie2oSGHUn27UY/arjqUUWQ5LTcvdaQxpIN1U8b6VZAd7hW8lzApGORGGItZf
1sxMoDj5AxtO2EV5Pl1c2tCmmVYtuHsP/Q/CseXTT0zIyTdli6/X2H8BmUePb1G5
hynx/3/pNOBbLVx8aWfpp3dM7g0juq37i4/0dg53si9TgiHEGoAdf5kzgc+9OrCK
UMRba2w8zYqCA4RQ6MurfUMvIsL1SoNdntVODCC8N5ct+GF2J9NzZhPY+PiMoxHN
Fp+rQAPzJwyC3yqmC5fnX8pi0ZR8CrnamyNamFzFM3xDbYUy57UiJyRDvAB+x3Qw
z6K6lum5bHuNrgZyWJIp5So0O9v2VaFh7PPr9zUHdSXRhXgNx7Bk60sFchk1eG1/
+dTaRQzdvF6T/RMsJSObm0pNEI487VpcEOmAE/McgQjiHehzM65tRl/A4ccIpNzg
uhnIyzEwp8RTgbg/07VFqIbAXCMpImFSEFVOVxX2MSav6LqfEOKsOy2J5MBxjDDa
rIjDbwiVMzTczZxjCVlFyYPDYs8zt/1K3uBE6OXQkeCp9LQeGl/sg7jDw8Yn7wtz
Gys0r7DWg5xhw8m+hYL1GyEcXoFPWs4BrfpZ5vSX4pjR1c/WqjlvA/Pbjx8Xu2qa
XpVM5x2SIrFM5zIJe5Em9Nf64BA3c1lBnUDNmeoMIph5J6jIKwH2nhNiQgppoVIO
O2k5TGAmRB2b4lhhSxUI5deHZlCQBN8lvDTOwvXLkrsIIIjeNkYUSHamXmps9+wi
8/4OOpBAz3AwmW8Xs+/1C3fik9Z9CovFy/IBSwGLnvOIYBxN0sHxuRK1OVVyXdi0
tDR5K5zhPmp1x7NzFLDmIkHsgu3xSnuLgsoSSmEfHSk0yIdO0OILwKx2cv5cXANQ
pmjUWG7Z2Qyh1zE0iMqMlfGdGA0dcXjTTLXmSjjBQPs6Rh4JRb4xugf3NVzr6tia
0G1zrETQnfcVGouVteT/Ljz5m2Q/M10+5yyxsE8BR4Eq7kkySd8Ppmw7+k74F7en
UoTgR2X4WrtVpwmYqjp9qinwdqZkD0onTsvYfXfAzddSLaYB5NfZ5nlqdu6ic8si
M46IvImI3Dj3keZiW6Za1qK4j2sLhwuZaOUgKFGInJn0bgobs8NWTyc3WUwd840e
oxkkay9ez6S/6vXX0w13vkBXjLHJwaG8KhPKWzw49qurZnmfGgM+5buA79m1uqyX
WAkMg+h1UNrNUKx6aiAfcDac+BTQakufpWPtsc8QuK9eTuAr9VMJsetw8VVafnik
WFIAKXE+S4Wr+3SVj76RFbeCulRd6I4SMLMXfynTaYkTAg9ey8mf0kkms/4VqRBB
plj0i6gDDz6rqMg8VDt18d+NWEPEO37RXJjRHn/9zHcDjrAmDkNNlK4hccJ1Io7K
obxMGIXRnvk8597Y3zLI1i5sDXpvNU7rkPYrzwpQVpBK8/JtNlcaqXYKhTuAuYZJ
zIxFsdLwsYIHgCTzxidabs+FM2QmFPzMQV6zd/OmEhSswqB/5GZeq2H7zOLEXNxC
/ldJigIT4Az8mmA2OssJ1CORfO5gaJePsZRwaGvUgZOkGh7alArvLe5RW0//hUu9
QrgmQBRC/8/vWvp0OgSRA9nSC1sFRGiIj6GZUhhLweaOpRKuaKzwTlXoIqhlvgiE
ZEX0AyOuVLyGVS2UogLeNx6/g8WtywuNg548Lj6jN8u+ghFUJfjgOodGdE9fSb2w
W0Z9n/ngIH9CrJFkwRpvznNb900X9hl8TOp3zNo1NW9qOAxWG5sCzu9LctuymUOh
DQF7Ivdra/jpecPvO7yLkadWJihwks7p0EuJ1oS69BQoqz897rfOI+MqxMum73zd
O39KMhjGtAk7uLIGiIYcra4ZFUUlvs5MB34Sq+OvSvXWDoCoSVgmLHGspSQSqAqe
Y6MbRAwtaqWlPjj/5iYYSGoEuYt0x8ulZDK4i7iQbgAm5Ptc1wCbJ9Xl5kE/z/2y
Cg5I6tFxqd0Vo1UP6AGJCKG1EXPVVb0E6ZMPdpRJ4mfeL/m1fTDkWx8yIRn/lHli
0esCfSRMyDqOCdB8VrYhLbujFWXw5fqhv8k1v1GxgDGZPcOd3sFv8tBj5e+dGboc
crLHBVV9J4GSLpq1p9TvgLV3TmoWiSpfkgbtP2ANYi+5I++oLyv9zKYxOMlvIs4y
VH1VG/yJqe6TXmAWkSQCckivm1KfnnI6EC1wvNECbLmmNJte5rBignx4kL3KcVDe
R1+YFV8aBFY6DKkzZq0YSCBKKZvQ5VxcYoeFhFgLdQaIlrlEcanecI3AXV+hMIcf
aIbbFgqIm7pw66f7Bip/Njc2XRQgCDfZYA1ZBEu5temSj+hZPvnW9p9+P6OECZrj
paE2RcmDk/m0bt6K0oe7CzGgP3iVfHmTW8KFdbW1JKMRs3GsVa2obLDzV6HawefL
oEBILhQgpROZYzbgRk5w17wWFqRAO66MiBnAcfhtoFciCX3LTHrYK2ejVLp3Ax4P
VJIIA3VbedQZ74TqxJRXv/GPx4txZMJeUePrmVE2gaPcrXDk1/3qh8gJS+Xuj6vz
AiIGgZOgexnyjjyDC3PERNwjSXpZFWr8PvTtn8G4VBvk4reCkc5jbAnBDuObHKqG
cCxbjuUy7qt33nhVikxQn2cHfgoC2l5dA3K0AUtkyvwSW09OLZmo2BeS2s72L9Lf
vObdHBJGHCOgE1Bru+yq/4Z8dGRn5R/pSiAnoeQzXlYPnZ5/neQdOM9RPtBY2u4M
TrdMLRM8vRgjJSiojmI1N1qBxR8XUZIm/HRf8w2Qr/ELkRu6y18hCQceCXj84EtO
Q1aJz5ib6Hii72wOj0L9z7OlQS4YDuPaqgbTWZTFL2GP9cVTWzVdrDgeJiELXrkk
XuQzjohF/hUy50D04mBOcwoXmmYHAdPSOOvmbBsadIDkf0vxou+RwHt8yRqozQrJ
9cRWQqkPG60y3/KbpOO5Mjqy9uyeASg+jWT+YfJllr9JZwQDPuzUlmpWzz5jUbVF
LQmK574vxe8vNgzt457MnSHwwCW4WGmfyCWMK9Tk2fOzV6NfAQzzt2APEWAg74kc
GIkvWhg3cLxgTZZFDOzYr6efqyyPxtJKZejwAg6ZVT4v3iuOQvPLgM9RRgKrHBTU
5ZqsZOaAsaUd/OtCdo2kDiMrJ/YXDLPzRZK+T0vh7xafMQjyfaySFXtCkgRMw3WI
X9DuUb7LJj9nwpklRZsgKKqP7HGBzQ5anTNOX9Po4WYEtzk5GiVoWXSscS/Nwzbk
hC5rn5TZ1wLdvdoxXZEZDN40qpVlBzKzNoNwZ8oZim0/T9/9tRehLln7E3K4HhCK
TruIsyiCOQOxoRsn5TEfUeGSqJ0JH2hgvpkQ/RpWEZbkcKiOn0oDWSh67UJIwmPd
ww7AmlQleMg64SdWeysEo9PrnJd7keOhmYfEzWLPSud9IeNfotXc2eYCd324eqnl
Qhqu5KeEoQBVOEVIRkPKxSwQHxOaI0a3xYOwbZ8fFSJ+BLOgdwSSkppEQZs9AWec
+EVZruqi6hQcC5SPONW52JvvN0eSLFwNHrfa1UL8Kv0+6Pv4uyzOmwE1Png83EqP
+hIr0jIGeIXYD9DQ55T/03DYbU7tQD2uTuqpvpokS/dTZk8q3IguXt54PoLIUWCh
u4r21xAX7cB3v9RYYLCLQQYyhAb+vC9XJLPGX7ARn9QHKYFZjpVkLfOf8Hy8pK0t
THdY5HTAi23YFgIIg+KgqoaNZXl/fyOLDI98GfMk4nOSgC5R59IvTQ+diKUPeq+s
eCGXyYMfpZAHVI2P3fyLE9AtYLAhEAIRimUFp0155f64rOFWJbSxqQl1MEQcgLUN
EmFQWhz3MspOlGe8xfAYvv93hF3dQDlCLQibnOnC8kGi9sVhPTcYNSu0mvT9mHoN
rjUUKKAc1l6zApFa2kg7Ssf3ALzovRZWcSYDLCd2Ln/UUmTp+0yG6DdL875JTVYA
KECqvPpFspifiv9TKr09h7/RB293PEyttc8e6F8riwlcmHcsyFfRm1kjdwner5ao
lKFLmUOUpypi4YMNZDEpxpnmUXVk+c+UnZrWG84EPqgbSGYAEFTDRnPFcMQiiewa
f0/sZoGX7j9dssOIcpmiCFYFnSl5PR8Kkv1EmX06iPkiOso7545HiPG9J7Hd+BKf
YzAyocx1To0UvZbmA1ahNW/vZbYlx9yoYW7v7TGg3ynWNVJwX0HkaAbxnvRj56LA
7QfsD9KA6Bn4f76AH+cNOP4zmqTyp4X9D2tExIxmjQio/MwObq2ELyULlQq//AnD
YzVkXbRPPpRbtkhiF+F5bxlaZrOm/Sea2gMJkoDsYz3qaBRxYi/2n4sZ0kRTzlGk
eS4G9drRZtTJyAZ1MEnsVpIoT1zT680e3H97UH34RFW5ApplgAN5HkZDe2Va/NmW
ZXgmSYv3xIFA5Rng2t+fnI3plkMvPnHi5wz1xc1fIDbYK+tQCVIQf7b0axeza7eQ
/2ZPHcepb2502hvNvfwRceVbI5ZWlZXDMuwYrgyOvaXtvObwVMgc4Kd3Rvd6h2EF
WrgvkMPkXAOFrvjUxINBz3CtAsG+Y0EP4zXAyMHhWV2V7PTZy0QRiFjNkCtk5Y7Z
kSNs9ctGUG3jLfIcp1aPwal8DwoPSV2cim1VEti7Yvv1HdonYdoIKaCt+GVz82Ou
tar2YuK7W9fW+qMF+qxxfoobAGdVjuAF+xSJ9xZQAVEaeDkiHMpZlc84R9GZzHvh
eoTpFzfG6+uBAQJlR3eo7DuobCtIVpl1sHIoTji7rfTki5Xj9VEqrCYsKh4MyKGT
GyXRj+OeP/RLVmTmkK6fs5+su4sOOppH+O9RE5slVS9VM5WHdlmATfQLcDuP0WO1
ot2mG7pspHRfrPbZPSmsjnMc8ZSZSD1ZG59o7lxkAQi5drh2/pKFUsRJ15y9dJ6R
GTLpd54EMTiGrpgbxgaAaoh8ltn+9CKs9KaxjE2AxS82+t1bYJBZDPW0f9VJMBOH
EE0YVhAzF1VQB3vYYJftZTiBqu0idadcLOkAnJnWslC1o1A1Xh/uK5z3+4ju5tCH
U6407fTbfFNyxdrhtuhNd28NaAtXbBOl4y2BWjDiS9af/IQGnE7KYH3HejXG6U9H
WrEumLgAXllpGH7JLDpkkKzkA/tRWPBJEE2n7OsHjN4l0Lg8Ggj9TfiL86cJTtJY
RiULGGQJxeyEggxD0qpHiKEaeau146v4ouSemuzkkREvUoejDDmCG5QMTlBhmUkG
EBFsOwx+z+6Ni8pOXFCbnXIO91gTNRf7Nrkq8CakXdwKPOF8qlnE5i0vb4tYoPgl
BQkJonox5c71xoj3C2LnL0+1oz6PQDjODNeK4xu2ZBlxWYagUwjPhLopLMKv3wtn
/WuiwcUWRd/rGfkB4840kuFdPp/uekEzKz/JFo5R/P1UH2mPdTfJQsSmMyQarwmv
aG19EnxQyGYTO/fXwc7CKSkKN2n/S4S1TsGz2cNhs9Ewqm/xY6wn7QkKgbcWPG8M
ljFr4TCwwwRUU/eB3FEp9KZUQi13CNUwCOjC+r+MsAlmPLLxWWwRMJFMZXNG/fdH
2wP33UUTkUpmL9UIGYTGHEKRbGMdl/BAC8QYKeTU1FY8qfq4pLrM3zVKXy/7ojtC
Svxc7bXbs5J6WuntROR1ROa2tura31QWx3XUjBW6fIoeuIlG2L1f+izThpfaeIGP
dEULlPhNd5RRarLyCg1HF4B9AY0Q8ncD37SwC93enLQiGycHZEaco5Lbxo1FDPSP
hukYwWvs39LPt5jhHvszTaQOlNmSTUAmqyDPFNm7hnHCtE/gUyIPopEDaLM5DTR3
7AI9i81oCpXQ8pjj/+tgcRufVAV04MDKhdeK5fpUzBORv/qg5Ug0seb0gawIkfoQ
r2ncyEHOZ2jN2GGxqHxak0M0uWCOnwW5B3u1k9fRSaxn7aYOEYCJGo1fq7++Es7/
atF+AF3xrA/AlvgSZuE4I3WBip5d7mIndG7Nu446JeW38kKexzX4LysC+ycRF0mF
HqQ2sHI07RUF9rUR0PyrqN6R0+RAkhmPLtCnBkL/03cHE92IiScKOR4eZ6I/4tGf
1fguEfuYr3RzPfodOyymRaXh0uR782Mpdbe8cLhM2p2NsDmRA8HgjZVqq8d8QJSR
qKtkKrmnN6nDD/9dkKMThoOSpUWXxIkV7wGokhKT7zkQIKddJPW46tJ3846JC09m
CjNkYzUfhBRVOupQsqJSzVLEbHciPMWyjxv83FFEQlI8sjYrL1iGQqnqBOj8Ti01
qTfkRvDym9fXUDQYCuM7CQn8TDrA7AG3KOJgumqv/QWvsDI6VzCy4H9YbGVYs4Fa
c0yfHbmZRTb2BxJ68EmbTChzLFwszVTG0NKEBsvl95uJ2wPkpmCjeqtWRA0oVgF5
PrKnq2FHO3rZ4JbmAh6smZ1UwAQ6teihjuwl9904GNtCE19GR/gCPJJHwbYlsjiB
6YhImkfdrDUyzSJBatY4GHkdmCjHALjdraCq8tZ1d68rTSiZw52svb9vsPMi7VOj
+67CCE1vuJp5VAd3Xdka53KNrJvkNN5eShKZtWCXJiAcBO1kRLCVr5N9O3d4VViN
aSAzLKSNYpjdD9AwppkFFUOBJSf+XH6pzEcELq1ow+Z3NxyhGdCO7zZzn7QNlHxz
64CcqaNntKDoc4Npdbecm4crCOXuTWm7sa4Cb4U0Z/JKZQwn81+CXiB2yvvh7fr9
G8gfKI3dJEcwRGE8XhJ/9M3oz5I2KbYNAmy06J4SWl3jd0+tIt2LWUHhFAR6ncvN
wT02gwfQBHQmrraW3bb9YGAlU/kglTdIgq6bU0XU37x+2AcCxXjpKxY8N9oz0lac
W6x8g2gHGfYii7C4CXOlMOLUzbSAEqDlhoXQvYDorUPn6C0wmIKX+bHaPR4BWzHO
O/LNxn5oEGEyXlbehSuoSli3fGtNl8ZSgGfDl1YHh5aCAFqENt9w1tSJAxOOmD48
ENvpKPSGZK/v3agZyZVFx2klohWbLRkbU1o61nIntjC0Z+8OQAHK1zHhZy2irCbv
RyLOKvH5OZ3lCxMaGs2p3jIrxJqflNHAJ6R5+YVpLb56AuElyUNyqZpFfHcDee4O
eZ6Usfsz7FtaNeMKlpXZOmH2rKoArwEGyNccvHarxJ404pWsxHZrJwfQ/mlX7plH
psFWDVLG0ZDDMztGlAnHfFgEl1gm5DWx+z/hkbUxRBnI+bWA4j9o/NmZzUngKpT3
UEC8B0c/BqzMtqLHpnEUY6QsVvkr0OtdS5be+QjCHO9xoMd3CRiWQ3dwH82Jd8R7
MKShbVg2cW1x86P4Syf+wgi54TIR6tTAcmhT8jnftrolZV3t7LpNbBVMMoEt027J
oDiil+JxX0/GlV9nBbrAE/kn3RN0lWU00HLngZBS+EjkASW6/i8Jwc53mE3Ukubr
gz2VGcdPrcLH8YwWx7wJbLNURfNr3Jj2i6ILSLBdxDue7I0HZlRaIe0mgB4WdSF1
Bc37jVWmlWB8VxJxd2sOnZLpyN5qRa+KsLwO6jpoS9mbVnLfZmLr+8qanJ3yQTKS
6r+6rEBU69cQPIveuuaU4WCXggohgKkDMJJYsa1gqBPD2u+VESsiLW7ErfUayseR
43D4DCscEbK7g9git1+Y8wKkuKpvFvDBgReirffJ6Tq/0BBszL+2ivR1izHUNjcP
WYvuNWZtDODMXuVd2xZwrzKp980HB0TSIlWG2llBo9UYi8wTXmzaVnLmyF2dzirF
1Od6VUO566VJvkWEHuuOf0ZrjvEHQGYGvI0RFY5HvAuhMCzemnKiUI7wOALFqHHA
Hzgkap8a6hdQtp81H5n5+dxF7YU/zaac4pZj0Pfhm5F/8bidQFkUbQIVXn+jmSkV
Txyh3Fo0+A5lu0DN1tJbdlqA5VUOklfTzqQ7jFHv7u+oeWQoaZK8O2ubbj5s1MFs
FejYvrwg+Xgiu0jUOHQouiT37VgC2Fccp5WNia0RJls1ECHYLIPbyWYstPja1KOs
IraZAaViwM5q3ekqnlmcljvJXOIfsR5Nc3EG8oypeV/U2dMEEKM9SYbw3CEoCfyH
DLF2/trzR787H7kY6vaN44Dm5GNN2p9BG5pZwINL9yY7s7YdXLMBUkOMhfsKct33
dAnPy+VQQOwKK0DGvYV3Sd+Rvbc3l+7CCzjlnKQfHlTftTO2BOT8yKLhgRgZsiAn
13hjfh/cPEVO8hIv8524MxjUUCTDfP41+ZxNDKerwG2bbSokvdq/CN3VZ1r0NgvK
qelC9vuheNKrQqdlEOzyajhr+oXEyGM+XamjViCIf1r4y6MTMsvD82WcgBRZ1I6d
9wSHDxZNW5479a0mLmpVwC6BczbbMmo1zBeVwLVQsnwrvzhSuW6C8WaCFeNQod2H
stnt8OyHFUQ4ZZuJrEPa3amIQvT3pTdDOVqVb9QAcTNHgNM8+/xZTo1ChV34H0of
IRYCbzQgqeErx48hA4ke0QKOnuLPQXAcpOiHBO1klvCozGqiJxVf6c+9IdcY3suE
xrsCb+LGrXCXXKYCXgqNZjaqjTVl4DoK8POtAWRU3Q8b3EieUmooTcs6gK0rxy6h
mSgDUFaQo2cSDAHfFVtW3ybwWOZMNO+x0sRBVjcQEySZVsWN1aVqVueN/fOEoMYy
GDCiHWfDYwWluP5DCNTZqeLvesBPAxBub1XGdkHKbfb63WoN9tvipeDCm1eygBV6
2Y7Gon1iW/R56DN5PiUkEqSlpXjTIwvDTXZuTTbrWpbHYvEbzhEygC37nTY+s+4F
LLPsLDRze8MT/wJ8fDPXXoSm6zXJ+9qwIoCaotQL9xD51Tv/BaI/QNVzKKOYOuzD
6ziGkFQyrRMyGpMpbUzA4m8t4VflkpfuDmkQ5IM6NA73++cGmSoUipfmtPL4Wzc/
CNkwhjSMTsxzFU1fqyELKDj9QgAZnkxygEFPeqoaQ7UfRzzDoD6VQK+r+iQxlHll
SymDsH5bWrwlD/TfJcI6LlYRGMeZSe2Ocl0TzkiXt5dw6ngztOJTeSC8LhBlAjqU
ju0r06gwYpUWXy5d/jACtiwEXPgnKehz//xn4ETEzyyaEdsWe3zrCVuTf9hJMmFf
QKFv7gkCkS3qWrWEPaB3wgAPhbw6ZMB8hYU/lM0v3F+zhNO1ZbpaOINk4WhTUcq3
DucL5zMAVZ7jxRPg/oa6cQ1V/chGeb9rWpHyyz5lPmnzVL8/aCIS1DBhDaPEAv2f
VmRc8DgF0qqk3TFhAgXSV87nhHmVk5lqFGL0rbtsEPjMInrdNgVnZ7WvAkT3QuJn
UZSIPd33MeAdldWa0aW1uiOYmOib0LTuXRzM+QhuU27DGLAnxOtanN7GUh4njhtB
cw8TNecWFNiYQBfj6zauASAv2lZYYh7sgcStoAXXKVJHnBqhUrySCmKYyh2pP1Hu
wKSxm85vxKEXkCgKlZAuh8+BCGjSCEL8xtkI1H74uiJc7WKCaGmUVGAbds2vcsPq
FdpcbzoENxu5U7cMJjzf66dWmOjRbA4Cd/97FBFz0Y0FXVbYKzLbptqAtmcnycYx
NC9V7K6TaoIMFSamCw1djkVUpq37O1FMgWL6msDbdQ50oZmYEhkAszkb1RpQpusg
URJw2H/PYkSd65/v9xGnCJResJFNmOk1SKfrn4rIh4ezvwtAShsT5FLiB4q/WtJj
jmATHunNjxjlsJygA7fFIPSxF9i5mKVpRH1wvEdNgJGkOdcVXYh5Td6ubGjqwu5k
9aqQrCjt0GjAYOi+fKNgVVFTcJJsKLvg4BtT4pMPba4mNqQC7x/BeKRVnpcas0M9
JCYcE9Jirl1fOLMwzM4MP8MJg3TCCDla++MfWhrTRq6Bm8FDJUnjhgQqqRyjpJ69
q2FtKXblMel8+kqU12iioRF4E57Hgc11JAu5c+wFAdSPmlgEkOJWmdEEoTiN3LrN
MNH/P6kS/+B4byT/9WDkRC0EP/NKH9DPiORGilqAHbCsnWjFQFmeaqmiOe682zmy
SqMp9YTOvLxAPuT+NHl1qHZ3FRNET2xahIN+rxmL0rfRh7+f/ScHLvYOSKZlcO44
hN6ZX9ThTwQmZB9vJ6kJLZhBPih+AhXbTGTsS+TWSSDyyEUJq/qjmbKiSiMYwsAa
tvbo6odYZKRXL0iTPRiR10GbZV5tRyh6CqpiwP+PzOai9/NSkxB5ZZr4GZCvm94G
eKdHGT0DHPNMa556q3qkdt+S8VrNJzasaDzwZXUIMJ+rjX8rWOt35uN/60CZLuy3
Si6icS0qH7My3sRTbDYnqUTVB+8ejccf3Zr5GTvMy2tbbqWgcSU+VNWP3+vlZWyp
/SW4JucXa1JLKGVlFPCgicJuECirTSqbvRHsJsjksTnTx4zw00g3yF/HUEBTcUis
t8XXKH7hQTBCt4Ybo2qrmRDFe4WrcGzM71wJt1e91qVozvmycjaElhAgly9ssd4z
4b+ryEGTrO+CD1mD+bGqK5oPMvrLRZ8LV/IJHIAT899FR53XPKXfkC8iTPM86NXU
YxG/kfLJRIDPDbgBhUqnnrJlGCv195/OnZZ0JevCuzSje1QXjrvzc0R5w4LBJ5pJ
xEqTFN9YtgfPBcqNIOQvZP8nijQX7eRIZHu+P0JFZlCPB/KPKQ7QLmTv0NZpDjzj
fiJgTmhmJnZRewiNiA5kpbx7cInaA3q4IeLGCOjuDp7NFASwTXmSSas9qcakOOfD
f+7BzN/zKXnTNpFRU7RscPr6k2hu3hdMlSSz9lECjCfFuCdqxb7OpH8026SZBdjM
3xi5EInd/CmHZCVcQxZqLLqcBeZw5C314O3GL6PmAkNmXXcPm7WViEwCe6OIyxP8
ZGnnfAn5UC207IcG7+y5G6MjnH+xu5AxVztW/T9fqHMAFtB3GOUzT/EXtuSTPoqW
OiQQlrhZU9pOz9wL4OE+MLoaSpQVbKbg8pf9/iF3Mz3pe2AXXeWZEQnqxtfeX6PY
vxDVYpZYzTf9BmiWLGoPBFbZc+l69tJclBsQ5fJ4lFfDTVtv8STdmHJpg8e03Elt
ppY1yPlim4Oji09/nhdLbOxmF/2nCvWSGlx49V0LxKMr/8+iNrXtVy1DrHyFpk8k
ZZ6Gx68PYnOovU2F7N3yXAzmwBQLcZRnzKUk4O+wUm6Mn2JhSkDBz/9r9BhggBgO
hG0Vf6dxxBdnCRLt2WS9BHFxnquJiP4tn82OwvDSbKmgCXQVxrjML23cbmdfVi6X
Tg9v8zlWArSlqLUGRJcsw8tSWowcmGbN6V3Rb1WJAP4svFpW8edzSw1f2qagbQxN
u52VZ2/9HxQsB4qqM8A/wDMuGC8GajEJr/8msc2lH0bDIjPwqQcvV33lzEEUuAF4
8W3/8QUqpeXUD9EcEAuMAPRs32lEvb4FAkUGXz0oyzlIMGnzl+G1GNEydhb00WDq
tPBr+WUJFlrN4+7Z9r8EzRgMz8z/sJ940CkFdcvpH54W8/ENoaRWfzZvjV0sdI+a
KsFYvaLhfWLk2SJKSIRo2uG+EkI08aRPGqmCO4D7XCdF47wCPYZn28QIsIn949mS
7OkgGHB0jLLyrltQBVXUZD/L57TRQb+1RjhR42UUmuXawirUMWH/AgV4Yv3eGp05
N67w+josKyoXerHQudqFFdcrR1j6Ow0G2N3f02U8CjtW2ExkO+mo9fR/BwX0yeQO
LTl5o9ykTONCwwMwNd8rwYVNYSak+ym4yy35aJ6N8IDBseeIiJp61Tfh/thcXvw9
qUEx6FkFe+vDElxJOZ9NjsJVd762KNcrFXTzmk6cRz3JZD6+wJ30Xb4jcUmks1xT
9lXWLsC6m6YqTRZR6IfdO+OvEJfzkH8wu40f9PKzrFyduTjapVVL4YqsBpafp/Aj
zcn9sgruL2tl0qTKi4RmA7KgFq8Tmtz2ZGRxcdRmdg4qH0DY5icRhvhf//zG0kR7
h8pks2aZ5oCdy6URgInMmyOHllawQcAeIkV8eHkSum+lg2Kf4Bw9JQ4lx+Pw7Mbv
oLzqJcKrcc52waaEwERDMi7YijDAiXcFnsBdDA0A/M9Q7pVqmaDmzcUewLaJI2mu
l7lLmHMvSOTOLbQtLm1OmdBOlKyW1pB/A8QitEKjPk3v2qZQTD733Ol9QvfxtSb+
dUQQD6DO1jjJtlKVbm7yu5JzA4pQpNYrMkkhpolOm6IhtmGhsF1sGl+HRgzLjNFD
RBxQmkrarke20SUwztsVEKN8JMLegQaHPthbD/Xvftjsap4A85AKXLL62J0a3KpS
G9+8ll4fgUnMT8mBDFnr7u29YKeuKAKi42plktnxppo+uZT8IWMsxX8um/+v0cJV
VEbVYEmgJeUV0NIYcsy/XCGhZPCmhPwRXMbqpAyHizUlPJOA2jbePFVjynEdro3H
GaQe+K6r/s/okokBlQteih9CYtwbZHKUOxwtTVLWIXuHHfAh4mo/BKH7s5jdvSq8
QIFLXauilprD7xlLx2vfetHmdlC1nlY4WSRqEnwqVwkykKY+Ni/dTK3V+5TBNGFi
7vlwc6TUZsy4H/OC5ZCEL6h7cWcZWdxbrWPyTmekYJT5vrkhZSoqIwaQjT/qeURv
9M/1LNAWCQs8Rd/f7gzOqTCKZzxBf15H9+q81OXOWXtuV+VzRuZY7Tqzi8xc6r/u
r45jmBYqAcOfsXcqklps30tZspjEMxYy0kCIXGELazAShaWMugLBBBVfTY6QI0A1
Yb7UGimSJU2uLZlUxfzE5Lpqnao5C4X2BMR3HMDLwxXym6PMuOIjFVun2Cu2heDK
IlD/GlIFH/qJML3e4ziwH5gksaVEwBWESB7aJ+wmwjlM2nOUViGGmG+92JfLlemC
iP2xhnzC9Gtv2bmgiQvYtO3WD+0V+PeyqbuA0yV/gu1p9XX2PFgrT1w5bTZonfke
SPAe6NUe/xuFnyeyLwDhtcocA9JCaAD0UZUpUzTmdGrjtcEffuOfhxheaVMW27DO
fwlR+VhCXM9I7YsO7TLkTOy6GVnttke9Bxs+wlyV0zNlSMNaHt/H8MNE83Fw3/CI
EPI4lSllgWBSfLF7Xir7V2NW3vCwDLLK7yJuimsLIMeoTmr9reK+yhqdxrWH/GQ/
+jLl6gQXJ0bXp5G+rM9rYteASQWjvVwh+s+MJZ5QHXQfoe1POrCSyONvyzO8axV4
Tnk0ogWAfvk+GOV1zVPmx8ftLnwOO8uGtxvM1nIyg3e4rktT2D7Ys/K0SVIHWpB5
6MQ+HW/XMcWq0k4OU59AmGaTFVJbWV4GLgY4/3xbj3drl9LMfZofljBZ+pilLzID
heqA16k/YV7fDuZZZ7Hu5l7QrZiB3mIUx9pm7UKib4JMSuYG6bEH2G4FXGaXJaV0
JMSbUNIRybdUiX5RO9oWtFIFtM0ssVMXaYWRLA5WzF14ApFqOiEbJ9IAb5tGv1Lk
pqP443mIJh/dSk/g/0sm1lsg8mHquiubUTwjpShe1ty3Bko9YpOC4PgJXkJ7vqTX
FLRu/jXj0LNVP3mC7h5xSpeRa59999WDCSEx3cIAaa3MzYzdd5cWwNBolNMQ2hJ5
75Q6OuM6bFFdGtPt8g31h/IigUg2WJ8J62XWqyKhYTE6IbNFzGUDL++vK/a+7Nzy
PCaaY4cdxU+YVHYUydMKENP95qxbAOE+VMK43Ce1CW3C4jRcFiqWq372hfkQwGWG
JLFKRGqbBHlmXUxHpcVX9+/8BLLJq1VjYKIeGAlxSI9B7BQk4rKQe5qkZJP3bVZD
oZW8/34iiMCZ+wD/gSVspVoPWoVRKMi7PFJ5DSnPSQNBZm8zGn0y0vCD5kdsZhv6
hHRxdj34gDahu17ot/15ws2o98DrBGeWX1i5wRoebNrSKg2y//2tqCEKe6W/Ur9l
Ru8I0W8NzT8iJiejLDbtOygoMqin8VXxod5uUy0SkJRYHpHJyCPfGAaJ6KgMYqzv
gVUQKZvjD/+BaBJs0N8voI0I9xXl8FEW5mK8pISkEU8bVoY/rZgw8DjAQsRPotyj
tl1cHuVJI9nea1MCmpOOQF8Ivoh7oz7OyK1gZA6VqJCDT3gYVt28cUSe/Phj5SMj
/eopsI3aemRUoMFH1CxGYH1DWu1gTYuSmE2CccCSA/4gU2KguVJIxsVmYsov/knz
4fQjXDS53YRKkRQvQI4mAjvXwlwMaSu3ZGOi3g+jzoNclYnOZqzyjPWnl7NQd4iw
/2GBZAwg8Bqscf2j0EChrUH9gWihEMpHwgnRxuiHpp3sdX+2fZaA35hUXovG+cd7
yXn51hO/4WqKN5KNIK5OJQOcZYJA9pBJNzgSV7DjfIx51dcU7PcBgNOZiXrCUNs7
XjMzQH3qzfYvsxtzCcYlM/gc0gnpTQe+VpKBwhthTIRwLxTsPi+b3IJyPrDDOAZz
hZVSAWZ08XtUk4U+8ViSoYCpBi+IjR9J1gAZicEGcsO3Y0r9GLHkbabFfCG3D6+b
KcADQdSR+LoIP/Hx3dANao2D6bcX2/3y8+4CJ08yAE88FqZEx8Tu9K+DenadDHkX
2LdDkyZ0venKSVV6hbODZlXZ6PdyyptfaCPbXFyWsRXomtQy3Ys1F+dDSikvGXZm
2nkP+iroDe3iqDgoixImd9MrlNmsFAbgJU5z3dmw8fwCgT0HelzG0/cLlGXnIPGz
JDk+EJVlDVMlL4plb3J+a1DlQNqtqxvuxqvCpuQqJRdEWgn44nsuvmtV8a7Uws1q
AvIZa/QghAMsToYbEHpwKh9UvENvdFLpLtJqo2NEcITTwZ/S/hIQ4HAcwEtnKIBi
Q5GS/GObfPop/besGmOzwp1bA6fiiQHWfMRaEFTQrobRrQnP5vN+xcaStxw7LEpf
IGYH/E6vcbt26Tu3SzYnas/Y8n/dFDS9ggriEhGtxMtKJcqdRhOeKBfz9yML0laG
2fvKNXLjOjQYkkUZ31Kc65gjxpBVvHN90Tr23Uz93cGLzdCBjFDG8IckwWjsIYFd
RpKbaR6d/wQS3YiqUi+mN5sI42DzfGOH3PK+mmESuo9C01ZBrAXul6vzdmD0Hi9Z
FbqQLwExsZ+VUuptQQj9uqo8NMahyokCXVqtNkvn4WykS4gApTynJ9bwcc6ll8Da
s+g5CH1GPSt1e4JYuqyqxAJPSoQC1qfs8o/18WslqgeDdSnNCeVLgj33+osFP8LI
21/bpG+tC+bG/BPeA7khA6/IF2H+lqraacpznPOiVQjHEPcr7BZiHt8sonFCRWvD
be+eGmqoL06xPUIBwrv91+hRHpC9I/RXyzAVAmNq5hl8UJasZgq78CPUZC68A/iF
LD9PQxr5njsTLNc4cLsabF2dKO4tKbmgdll1WBDiNXF71x4hdKm7vlQk8rae9r0a
kkk8M1XacsHi8H0i81ef0W34Fog2Pv0PKdLxnUMpRv6COIs7JsFG4zIx5tJtjf8e
acHE1F3+pR9vNKDxg3rF6Nyra0GPbnVPu4mUb1Wqs1dfxgXhKbKxbDKDdWyXHjuw
BMDlS8HZ2NoUwEEztcsd+y9BhIWQi/0cKAT3KcPboOdRJmxYlLiYo6V2tKo4BCGy
OCRbEn0qIBVRAwSJrOTJcV1s/is3sUjcqq8/BScbFLDyGuAMcnWWCYkY+P7cBUBd
Egn7UPJhalnEVRd/4KDBPqZUM0rEVpa3xhACPvU8RmEHHu+0DkCVjFRjKIG82D2C
Yeu/2+YuYVf4t1mkscBppKt7gnPnBW9bcmwAwddp2QOwvtXtoBcoYCZYgy5Skh91
pKZFFUr4HYEndJyP2yiIl3hhmCNqGMZyQOBIFkun3l7C345mBgxYf6Mp1ZfsCVmj
7vVygWxPzH/+Hxdyn7Std1K00SZ9LikCcAqkKVaL8Une6n4ElceeVXYHyXzytLxe
vd2rLczlStYslKN8SL6TB2Q+8bMs9OYcsSBpBJvettZVjTtbKlfheTbj43kh2cqH
aVoYQjgZn2lztfxLDtIbc0erRqv/GjlAcRpU/n6B3uYhSTNfZ9XI4e5Q0TsO2G28
fYqzt6RdJ1xlrSfEKBq5uKTQzFd5f+B/VqJIh1HVHMpKOVWClkeJRFq2yek6OxKa
GgviyBIClX/IOgq5Rp2ChhBvdSmNtucYR1ePj6nOU1VJ9NdoX0yOeKxvlGISdMuY
p0VY8RQnTyKzLB7ptMC93uqH7LWVeVJdeu/2gQH+SHPvV8140kRovT9PaV3pd/tZ
Vrmx2I41KCdD7NbVh/5gi9kfi2NlYXXmlWThv+5GGTXTINJzGCxkVVVn8XKaxcni
fDDC7bypjkmTsJCZ052e7+N7oZbzAR6CiRA5V0CDt/w9MjPWBYSo2wB/27koCtsH
btHdodaf6vemBKbkDxU8ZTnfYzUyRUb/1yegYRF7iUNDZqvCD1zQHBcnLOFOYxw6
YGJz4abyB7msG4AkQP7KW3BnLfJHHU2QVcAcUeSCxQ8RE9dm/IeJvzrMDeaNHQEI
nTkMmOV/SZcdblYa+MwNrqco/NM4yf3zrgkwhh2Xbeu0zLukyraF4O97hv40loyv
6PmcUsr38XTgarJd658tt40IA+Y7aQTXs9jx8R1uX60FgMjI932rrZCnMrc/CKl4
T5B+1G5qvxABFnIEBtSRr319jk2LuXeAkhbwhZEh0w93phgzBCu7jmTjzVPKQU6h
csahHH6jP1Wo2Au3NajFQSWPAPFaQ4lI1SrPyB2g1vTx0Lia7V1tfwb0pP696Scz
bRhQ/zDrBlo7qrAkGVKVbHEZJer1JY1p0qSyIIvMXCE1G2sm4odg4s9V5kIxDHlU
vXL5LBTFMlP5F6DGQvXEXWPJH/evg83j2sKF2pmNbkzFbmzyPwquAo2GUFOE4Yzh
LiQad/tSeo4NKmIHXOGfb7eS0JrY53ZaHx07a4eWBg4X0o40gGOE/fMwMQ8iPVSM
Yp7daCjwHGa3UG6bYXOyY01ijadlCduQW4uTLjjhR7ifmz8VfJPirrAorAYLQVOV
k0j6NUUsK6mrWBUHeGjlq9ukMcgFQT+WQOzBdSQkPjJem+SVng+11kQKsAJnPN7G
p+sJ6DkPQWjP4iuZ5D7AMKabsrU21FOgTa8jSc7ZQOnNo599TknkNRWj5snRuzhE
xZxkOHQNtMxoP/zuPXboC6hRw0hi5G7TNumYp0BU9aJmHoutDZP9LMrq35c6T4Rb
oYqGF28H5lhEjQfdIyC+15rQ8xmb+FzpofprCc8qAxVrHSMswRKlevdXEkUgGhCs
qolLVPEcauskxn6TIKfisrty5UYKRx8xz5VWym5wpGYqOWeR0JHOdJMUoIzzd0yx
THpcfZG73fubeYtgPw6zXmmDLz+C47OgdYj/oR5JmlQYKmU8FLM3j5XMOgl2/Tx7
2Wk4OmhYkPo8IoeJZSbwtlKMpBAgIaLBwO2mPaJBDnT6J+1DlWKMsTryNKrKNKj0
kFlB6LHdrJy7lTceYeiCMED0QvsY9WwkOqtKQJ3BPIYdAd4bkMQrASAtf6zq5uLl
1vQN3tD/CBBmsVoIijbsDPc+fUYkpI8iOCjVQYGR3z9VD7N7gJjYrTmE/kOAxqah
qnlvUiFtwYhdQU3CDxcKZ7qIKJ2LCKqwcflyfDuP3mNABEbr4TiPCWZzNZMntrma
N/vCdQqmptIPKKGNeigI18dX3lvyrpYCkXiCkFwYzGdYPD9BqZkHdynwcT8zO/fE
OAI+4tKvVP4NFjCSlTipHzoEG1aYhZouv/UJv0xWZ77yReShMPfqvtYzDcEpbgGN
beWhiB+YaEWYH8QoRpB0T+0gw8A9nkh0vIrK3tnsU0zNLr/jgrIasTbpIyX37zWh
jVfK0VdIcqlvjkW/52ZE1h7QmpbZ5ug6hBNIDjE9XyXaIj7cHsF4+n6HrMICZJqn
X4xgOqI53u8Sldnbf12RfU+jU5q5A9kMGjs5b+uwgHB3UJfX1CULb84xhmOmhs9p
UHZwn1ERJwHsBT5pzrQ+R6eBnkHn6GxSpFbz8QxMd91dbbOqULbi2miHdz5p3ygB
ZeAIjQCi5egALAOhcg8DV8VeKN7UCfa6c7tFaLxHUXa3Eay7uzeuEMZDLRhtqhlX
Pk5XaxYDKFMjZIHmf2AyG/bNIuteJex+tc1fzRIKYEahar8a2DF5kc3rlYYgZfnT
Zg8OnwdJhhKSkXN00wX8OZgK533l1XrRw7fouba33yefU3idzFYfVAH8NmxvBpVs
+9MyEgWAJgQovPFWnoYdlkZXSNYfmnKIEkZVq7ni7n6SfOa7U2pljOmKNazWzL4t
FCq+LBe9W6endpYsZlaOX2kJt+PetfbOFZdMO5bQ7yfFJvyj/TPqktI88VSFbvGV
pcyN1c9zGONnyUiDUSYWRtuOySMdvluPG1OwRKnxIxJVNtDhkYcbXNsqVamFJGGQ
f01+UU2dRFo+cu1rCp1QUA5sKIsOFhsObAYNL2jyeS22E194e+j+b0Ran33Z85PU
Dhj5YdYnLEqPJqWYcuHeF8cvUOgzNfIfxxGNBGzP8/2y3JjcRcF3WpSp2qM9lHkX
0wURGx5tEntioT0pKrdpBRMn/5BJCEpsa727uCChhJk40JXG/feOu0PdPCXahf9l
Qvt3s+EMDPSGZVTezMS8GymWGGEZbxTDyZCWPKlXqJO2GMfn0gYj6VWI+IHwvoEZ
8Hu9i/MQ4ZiEt8rqw8rgeREtuzh62lcM3a5bkWuJxCkUs/9V8KEFsLvLXJkxZF45
kX5xvQmPf+YQjF40/GZu6USqEZWo7+3CUMSnIjw5jUaoYqt4ZupJZxaZVKO1f2nH
7SifrUGITE3S22AtrD7s6lmbBO1BZ/wOw2ANE+jvVGhB0INqO4KIkaFkZVYu/PIX
E8WCvKR85XM2i7VboSavbbVS9v7BmNv+IidMBwguYhdOBvCCCjMR68rmrBvo6Iqp
M/lXTb+X8mvPFPFrjQJBM48FB7E7Cl/8V0kOoc/dIkh/p+A+skcsIykts4WxRzS/
rUiBa03xxj6ztXbxQOdI6uWbf1D+q21cOATX7FJ6mqpN9PG/R63EIoefikazu3RW
IVLUxRrNYP88J00PMi5qAkNZ0nrfJsBUcxVHL5xwNEFni984JO8N5ZYcdWX3uHWw
4ME13US6fEK62t1O96nUyOH2SmYK6d1JK+voDkuWrcP+sQyDK9gX66pf4xD4218F
w7B1t557TYIeSwL19lYie8RLcXxpFRBFPyg4+4pA0SrOTIhpExVvPmvHNUyJ4SYX
SIbMkmf0liAJgEYw5ozG6IQOy0bZdc1sgglrc7jBw39NF1j62hr+4B4yfUoKuM2L
Q7/iTepyozr11LFi+GDp3j0PylwImvYEmdoVe9VsbDQ2HQGxWUJVV3nMOln8tOyW
CK4Bhep3M5rimyxxuFTwGtBqLxSJAoMneyupY7dcDhYv4QID8+JVMYyXCNLNYdhm
TPYHvcovkUFZS8Ra/x5hybTgns72Cl6sUVU92Z6UrtrtuHrL93c2dtns6Uutwazj
JWchpvB8UxLUPEpYn1AiNTYBDAkvBbOBiSb0uXI+tPugAxh1GLUKKS4X0tN47CH6
2kPTWZAJDJT+p8MVEIOvYR8xvKImiBS9JEoWe9aeooCUFQTjj0ZAAazRPU8+bW3k
iDZyXNsWVQIu+4Ieb+04qVlPod8UHv8Juqz5Er6NzgTyQEO/xZR5DhIK+sn69Dnn
1Ex90PeCsWQ/7W4LE8DH1bmx41QqWaGOcUTit16LoSk2FC0oMNUcQ0BNcNcUP+KJ
w8jz3/R2q0ES2nWUsCZR4YbxyUskSexA+u+Rf0D4IUzJYiPzGwS9IilQvivm9C8M
UU0itt5lmVFL2iMFsj2GU+41thpzx1+AFrNe6pbkqkLG2yIl0S7NvKSt4JVSFFSe
ZL1dEqXgy3tQW6Pdm0gqiagUSwtnh+Xw4CCVApRXgKJotP4hxRJIB8FJO4VsA4En
5+V6APDn68sJRLkVZegOGVEaN/YOQOPHPGNw82X4GoEPAYPHyj9WFqQ2GYD5w6X8
IvzyTlPiSGyozAjYYKTK8dj1QrGEO5Teu1mJj2450qsb31DW1nRygHF4LsyT8P5S
eKEyBlBmkCens2wC/nNm5dn6U8Pj5P9Vxks4s+UvDv9eWWGn6Sx/TMMlA9bY4FUt
W3a8cnP+gWEVoHGCxkB+EbPjKoCe4Mf2zqBAj/LY+DrijsUm8XoKO/wmbM4zjNDf
Lf8WMSOuRmjMnOYdk2HXpueXsWhV/nayDROKhOU7uV0ogfv26PJXaYzTKf2TywIq
1oUazSrBR+Ut9OrS6kOKVM3f5TwHq0uRETD3V0MMvIeEHiIyLZ0/emfmK/BJ18Al
0aPaCrYbQM5wUWv4bzwvFcQBNuf7gbVPdHa8w1DxfvGLyH3/3nHbyliCnvlBpaGP
wAlLdsvcioTws6YRdQJvg4e+Owc9dkxJwCzuhI06S8GuKW+KSL1H2GM3c07ZxURz
j+NbvgNm/x2OqqOrdcqogAMnSCereghgP19zyuDU+EXVo2e4Sw1gcdFGSFw+I4VX
FxiaaKfjQzD96ogfm8PpLROdnUUYlVmPVPMX056RzHafz/sZYKZZXiJioVGN75z3
S3MG+R5OGF5ptVZvygn8bR/Izwc+l3Bl+fIjiWx8IsL2+YgHPylAYTM+aK8PkxEx
tXbBRBZgkYni+IyuJoWIck3DeUn2M96DfNzIeBgfqM6xVEan0C0kqp95cYimxEdB
r0Tiq/sWAnkUN4x3iHOzbJv1XeZcPukCPFj7g5wZA21BQfOR9ng2j5wgYc7W4OTT
YdH5uGo+8KcGBjR1q7V7kU/Tc9wE2VDuGpQba6JMoKa7nsrgWZOemQy1FSmZ/hNv
fy9dxvhb3Lup2wnj0k9pazOtcz8jU2eK2hlEwhNAoGATp/DV1cviM9YKW1U253cL
9tWGtDLQ1+KwRWQqB+izWrc9VAjl1AGa3ZP3pV8ztQREN01r8tM9zogfLGqhycip
8n0pUcTKP4BAUmGVp+qoHGYT1s6oGIvldwY7X/oYoj5CRphL7N+IHcaGP34JLK9+
OBhIqURPwnbeqUJ7zM0B/qpTbujAlGK09/iStxbEvpJxLoXv0TcqoW+wxog9YM+i
kekWtsd5f0JRyt7VkyDQYHY9Noa5aANbXw6XkHBIQlxcGKBgT1+N7KygCgNNObsV
8uIAPaIUeyok+5sS8FhjMhU2M7210+dzAGeP4boyvUydc0WOaiIkzHx7vxOqGpjR
qfkoVbu3Vt/x/MgosRijZlsSwBZlYar6nwUKJqCYGiZrgBJHo7eISzm7XPvq6LRT
54mvYhIMVBC8ukSFIXUrvQ==
`protect end_protected