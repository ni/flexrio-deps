`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzltuEBGe4K5uPEdMunCWo0h1G7JJfIh1iLr4zXdO/Rhz
AveWe+kAzLRv+HP8y3qzctpKO1CV/g3M5M9jEJhfwvf+NG62DSHN+vlO1XgG/zs5
ruTNUwbgsQ8JFyag+F0rH9JmSO1IFyfd6EG3We8uS56WHIZoGiOauQWC9AjOFSGY
tFi95e+qXS1uOoOlskvmRP1ShEzkwaTuu8bRPOgXzmr8KMEXCvB58j2j+iT0YMaW
6idyAWo2XoUsmksP1ZaYQ+0B0GTVAzhJpqs2wKnOTkfkG+W9xrGqqwNICJ75S/Ni
vHDTdg7vEPeiowTA/4SrLZIkpTx/2f1t+S+9OJE4efv9j+5cnEMtp9x//DLLxRts
FVV3FmTrUyOP0BXtBLu9ckNOL7qf1S+8czK6ax0/o+axlluZV3lATBddTzhGQgDC
dZWGhw4F4STH5R/s6hjt5Oe4X9kJA+xjqyoZc9KSN+P2+NCFGKJEiuFxK38GdRHM
hR9IG4QUQFK5hXdmX7cKP9NAzNjFYp6j9QVFRoWtJAATggzScAPA+sKbXEsCfNn/
2uNe/1pLH4pmMDMS1lusZ8CnximTY9/coA9q29B/ZiUNYwxIsX0koRPaPmVX70p+
YPHJXIWi537AZ9At/PDM2ZgoP9LAr0+3P7T+C0r81E9nftFXPXdNtYKlTrP1rR5v
hFNnxkdlSCb32CD9lXh9vNUQ8Lz6PU0m1tbcW/dUispLEg2AbmVLd/ukGFNzjykv
TH+xvPzuOBrv1SEfOiuueqlXO4JYhjcjQvHpduZZ9RtTEe4i4+5igjpk0zfsugDF
JUkRRl9ic7jCRZ2e4nnwa2Kk2o3VdA0gmd9t9LjUN6C6sn34JZi4pFlokEUuZfgA
rhn298mLueIA1q2MHALmtwOE2saGYG3+iAdamYFe+iT8ftg+/ZtlweVQJvJzPXEs
h2xQ1vyWgUwu3nqLLxOjQbBOsj6MjZ1g2t5uAJ1JVrLzpqRW9OcySh3AZH24DuXe
jXid9cyLeMeSisHNF2SQ5tsuEI8r2jtWAqxcv7aB3/z+hLy9ViioegEy3ONzdrSt
wQA9UA+QKM7Igelt53pLS7f2sEq+dU4Re7KikETzXeWJ9uftvHZ+zdKniyLL8hqa
2SZbVsTWEHFqhNsQPV1NU9mr/oNzxcW/tk/su2QNrCSiUVQzxzDAi6vc0elieNT+
h2wuL+ymMKuAfw7qOf6ES+X1kSDPBlM5rm06iWF6hIWGl0Y9gcCR9JZfep8HQiaF
lIRvT6jCIdOFc11Rt/Ffj1RpuwKmlpQ+1qFXpMJhk0Ttfx/zGSGaVGVB8q+UfTGy
hM9IV+1RohCa2GhEw9aBFakvZa+CTeWsmBHOvM3pPXJsCFTTNttd/fxhioQ4UEKY
umb0eYWWRA1BEWsoVEGF67rMjrAjhtP738zvwynZ0Y2fnbkDBlpW9R3D16Gp5NOK
4OJ7jYlvop/tg1dOJOM/arQ64NKmiFO5TWOhkxQZnIxCVcaUim5c7yILyDIt/eSb
oF5/nrMfwaxpebT33WXGGIOdZh+wB74yHtaQ4YJmXOUFmTeqkD71ILWdAygaY3XY
MRoGc9Gjrui0Y+YkvFuCiMOHs5cTDPmimPf5JeNmDwUz7kPlusiXXg4J1ypmNk95
hmDo2F+KPRe6vo/9ICqhoPjwXvCQXAu+jdQVLPYvgTn3/1agdscWEAJCvqRFo+mD
QFWZ+dWwi30PUK/ctbNPLqIlTxWATUCcJ/pYxGiamnP4SP3BNrGwYk1LI4nw9aZU
sMdpx7rke8WONx0REM8dm/0HrHAT8ui619X/VHa5J+2FCRrdAhKfAkgV4riiJcI1
4gIRtIF17x37Z7mPXvE4fpV3f/DrsE0SnWCh6REczZmkQ7BmaY1liy5z2Eq4b7ec
ceYhDHPNyDfOQH4xbcp7EO7n5G0smhsT+rKvZrg4KrOcEZxYfZ7eC7gf3uqvdfnB
Jj65V/fy+d5COLU8E8X9l1l20sQBWahtkV5ghUqGidGug77BHzJVhbU78vEV2X37
nqddBP9J4YtBuL3yydik7rhpYrvj4uTRQrMCYMQnEsX5XqgWELqDZSrBbF9GpSsO
SoaNExyK3Kt57/wJ8m7naJYYhapUwMkRJ2dDyK3bpIUJDZr29IwM1kBypTyRNpfh
2aBGawpH63X9fKAuTcmPHDk2V5V2mg0rZHEvJUsTYL2WZL1LchLCc5LvEMIW9i+u
JWESGShKH/wBQyMohswtRB9V1sgWfd9yZk1h9H+/WMoxm3nXmsLIv/SOWTU1E6MM
rG49UggIn8ZevweiDyP5ZzJA/yFIFbCZ4n270l+6PFXV79A5BQiVNtcp9P/B9mjZ
bfPpiA7Q51yNgNikxlzIwhmkoA8bNJkhNvnRXe4nBICXW63nBfLFv4E0hPJqL4Lm
wj78zILp9KSMEq6Z+Ai/Pn4kjPUbircyYB8GFHyNU00AIV8yzD9qi/EllIcg2+O3
CCNWLk9NXyhijk5/kTen8bnleHipyIE2pN5ifzRW3tnbgTNoXVgFWxLv+Hf3P5Id
eUBQUpIDLRiA1t2HxgF39YZdfPMv4lQuLGTjt5XWCorlNghg199OVfh8/60Lj3yc
h3yIxwkq+fPET5Yv4tN7RsolTT3CB5kFABrRu7owTxLMLCGD4S8BB6Qd9BORRBrs
s/UTanmmCcnUOnVOMKPo9h2Kc8tBeezPXz22SpeR2J85XvIAIHJODdTI5BPiSkDZ
hTeNqlkMny/gcAdFJVttRFjGvxEBORl3LrufgI2MMw9ZyY33UXsn5cYKvkl6sxzI
3uCAPpTBzeNA2yfdRmvjBrD8883h8WxLfF4Z+j/WYyXutJszkVt39Gs6yqGQP9ot
hU4onpnY2vu2Akz9Fo2uJXKU7H+EvLy451nqZaEY+oQ4c1I4blNprmQbQSbfCBMg
sDjEP3A3BdGLGAverbz6fws0O8oTiwKpeHVbzhZCS+1lbGy+zR7AfIxxmufto+NW
UlxA3AY8fjAJVCcePO883ZWGbIebGnkVDyv8n7jtfiCkvEHb+P4mhIR1QwAJi8Ux
yChrRQozFcikDhnzohVZGu1v5+WgBL3pol0ay8WCEYMjvhYVanQhs0QjKTgIlavt
0P04uTdZX5gqV8g6r9uTVOQqF+Zt08HrK1BD2iF42u/uBorPtVjZwMTs31YhTmPZ
piqDcgnNKtp4TR8dR0AaBYKRtphYKlf5jB0tYGJb11aTyMagYAvpBgNBdTvBjYc3
/e5Cj/olV4wFdbKzg+PaHu7JVkaBo6MZGxh2cLTP2U769YG9nFdHsqhDCRGJdZgX
1NTWqzgocRYvEmeefucT0Twj3yTQ0AoY6FrN7BaCFtnB2OOWfLjrFlz+FDbWHfOU
vMxVwW8740okdLCKCkJeUqwc0Oi1PYebAiIjYBf5LI8bLflWm5l/O4gHVBkbXS1u
l3iLnls9iCRXi6SI2FKAOyp2FZf/OIOv0dmyG0LIKzMHWEjM+ZcP2CPVGyeIOR+W
qy0V02ReX7iLVF0DTp8hJC/n7qL9zASRu3odlDaS2880nOKFcEnoybUadYC0UP0j
pZ1atB6+PR7xl9HZIM7fPTnqS4pPaWfKPjNUz+dEMzYTAHQCb0xanhT5gQnUrrDw
OqdOGNw+BH2FN+DxjpTUEwHOnBi+kikgfMuKUHufzybKmxryRPBB25ayQJ1Sdqt/
TxjJvXDtKXwCKDdswpW+oJM0TBOqAFlkPOXJHyAQjZgUmF1HU7jY2UhtYlwdUvdS
Z4n0Sq1UoVtY0JbscwYUiK4fRzVis1bxhA9aGzCtvIpi8UBxjQWrfDSZB9IIibkr
TvByhSTrF6+zwmWttfzHpjmwu7BzLUfClG5DD8xcV+AbtOxYL0+ZW93VJSq+2ld/
95TxospTy+/CYg/L6QzON12oLS+giJ+duYupoXWx6YoeP+sD2zAEFYKmgHr5z6jo
rQMt1w4aGVQWGWwt1IPuH+0dcTn5REHG1+uLcqktVNB/AbLevRywOI/emJaS9UGE
YmeRxHo1U4DXMvDIAF5/AKhIbty3yE0QQKN5pjQehRW8DRkT7KJtTkggIMFWi+JD
YTnspT/1mPXsvqHBhXmUocmFwv6fpjoHqWgsphGaqSTCk+Xkp/0rSZJeTcbWM4/5
gsvOt9+yANAly1t9qIhEp6QsSBJFIUcd0WAUDBZU/MOXwULhkCv8xAQu4zG4tXqy
ixIGHA8oerMdh3wjELW7GKRDFnvFnrb96hDf4p5H5XT3J8N0xuspDrghg9uMkOQ3
X7J19NAOXuvvX/yJcC/n5I3N4HImocV9AGuJCVDVsuMeEbmduXDO/1xGFuAu+5T0
VS/VRopv5Rl/skU9Sa1DEaH2XT+zLHePoh/G8+zqWiBrKgoRujO9Qh6w7crBhNru
FqiArikpDbf6SqnPE0+y55E0bmD/20/uVWPg51GWOZAufHhJx+t7Zb7A350DH3fd
UPGQIWzxEyKEvw9ZSfA0lcp87RWIqLvFmXX6VUm3+xsu5ffmOvZpCNKxZ4Wy+HDq
/VjYxg5fZNbhMG1NMF8oB8JIRbO1AdQpoakwlFOPHGDko1CyCWj8VdYGkY97fmpq
trtwwrFelWdCTC+ZoN5JsSX3nCLO23HWzdUcyraSR1JO94TFyAhysNxo7smVNIV1
m1da7fujwFYhw99iIXxMkwXLcr7KK9yskWNl5B+s3Nw3avq1NE9+VdfFooCr5TJp
jblz2IfhKyw0RVToyKrKUOfHnZeqrT/oD/+ZGfXUQEClXv/UCSRhzZpQlv2f6rmD
jkGLvGFWZoUqW7dYy27S+JVD4e0TB9rrS8ASLel4J4eSegq9rqRARMu40hQnGw4G
E0GBKwi7Sdl5Wyvo8Syl5yXTS8bg5+6LN5YzA1T4KaxR5n9rQBeAlhB2ckHiV2WD
r+Q2bbzSI5NtOg/eV6Z6dXb1o4loSx290nVVt6r24Cm9JKMWhdA2S5P/9hd7NcGo
ePSSpjIzm4P019O+4XOF3QWAkaM5CyAwJV8fI9dpjsqKbysNs+xOQ4S/llcxf5yg
yzqgGMNpsIl9vJuitDRgRH7k9sXoku3njgIn2lkl9gGWwPsVbvVy+vI7HCIQrM1D
GcTGZbr1P0HKhglCo8CYJ8Bjs6QclVF8P0YMo5Wavm0eoHSGu7zhU+XvFkb8/M8R
7QWWPm/j0nT/pHQOhbc0zctC4AyvFCsUYmO+S9qXUW50Fr6qfhqAhiWR7YQqVMxd
JJjnj/1yaFYjxzx8P4YISyloQ7Da6l7H0KLm5AHCgVIcMfADEhnbN0KcsEQbX7hk
F/XORrDUJTnv1H6qZFbQ1K4TEYgcFbb6On3v7UY03TBleLGcjl5abWdJwO3u6sHz
u50ZvhffZKr07wk/aTu67dZoWd4RX0cZoARL9iB5F6wH+VL/+v6ntlLK/7hyux+0
pDzi/cI1iAf7siVvHwaBJlprZ+/7qeWwmbByoYKmMJwZNlYqDVjOG7bkDuaBbv8L
IJPiW/uzLoKOTaJdLBGyPTt1soZIPe/hrLvFFRn64uFkM8QYZ7Hg7i1q2I2y6Yof
0Hr41eKH3wz2xi99Bt3MIM4mjP7nkk2/Q7hbBpVOE/5sw//HWJSfMrlAi4nMjLrP
PANp4sOOATaVa11WWwqS1OOHaGZf89S/+k8spIkv+BGgvsObMgCKd8h233QP0n/G
s1V5dz/AimfVIoo5SOVXIDhpomB6ePlr8J0pO0nfPz+/DfyXUwBFIuuVLMerGMje
lkjVP3eg2/bZddzfcnnHr7VQegnrt7umiLFsBYxolk/cR3LQ20rJZNhGM1+4kbpy
EHJAB0QB1l5edh5GWuLtWwvIzr3fujBh8oPIWn/RGrKM/H6OXkAIGmHZaKG+u6I3
tLvE5/tcKY3MpmNtDSlPvjOORPgXapFORhBHOqgOJcGtyyXYLdPB/8gGZTIkLT+z
KSRdkIfALFiSrnsJVJFqWtWaxzAJwnMp9Br0Za/ltIfbiJGuqPJ57S9wE6L+plrx
VkurQiS2KTIUBWjhWoVhQlPyRzxXfaW43mstdpya71RF6cEsy+Qhi0lQ6P+5t557
HNlhETRZeLvaAhh4e63BnCSHJdskpA5GFxpcEUO3fMj23oyoy6USN6VWp9J60VxF
Ai1dWtXoVl90A8Lao0qJyC/jzDOJfCKNI6J7g2aPNgcVCu91B5/dWDUHfBOP000M
fYTgEc5kCxHc038bKOecasBavMlnn105NYK+8gN8uaP1pyB2JEYd/0T1avjEsUXM
IgQoQeFxC5U2zT2z40s2qNSBZrnXKBPf29HPt1TyN9fD14gvlTuQQX6d/wwuJitW
yxXABO8x/TrGWLObCw454lwqnjY54NxdNauIRnJeTFyohSaZa+mGz0dRe6xXfQdJ
h8RV/LFY2mEmv1CDSQWAQdLQy1WGwyS7FbZ4Ws0NtuBcTDCeljvNRCE3GIGyKNor
LgqxgYVWO0a+6XFeDjF5P9qFck9r3O5y1zrHwuEvB71iZPxevRbOf47MGPiZp8UJ
KZRDxkWYUHLyFJmMeDvT/iW9LKSMnPNkpYTX7XTl5RHI9QzP61AEsKym3aUw2OD6
qG9KuDHci7z+fT1HiXWO4/F7OkkfH9apq/OdlTURDF5Vl9lHD7zbO+FxwVFXLHIf
X30hPKpSh/fheZ1WbpOTQX6TztdtOnlWdv4DKlSJE1c0tQeWoU0CcyTxnu9BxYgi
ydqBdZWBYiTEeq1aIZpDWEzm/unj3jzLD+dEwcxxlnehNIgcjblso+5W6Q/Bh43s
XIGxaLW5BL+iRFiGAAOXJvtB+QyxftB2tGYVN5JRCoG9pB4bw9Zntzg3oi05Qtnb
NS5ESC1BgLXdPp26QQOyWuETDN2PfkTtczNoscMrqoZWqFNCzvUoKp/de4TbGd4a
F1JN7jd+0PL8JPuGqng0aiZ5xCWsVa6U+vfMGKqjDj4VefEohpbJwNaBUWC9hFeC
V1G7Ts+njB3oYK2QZ22Ctdq9Umtc70qQ1N8BWbax/3dJAAsWLy7hfAL27I9iacbw
/zt997Xz5e/2p3qGLoVX/KfWlbVwZjBYMg3MhqRzEYhpW79l/rf5FRxoPpzlEC6b
AcAycnODGb8W/A5syi3k02O2wrlx79/wgt+GU0/nYgxwLz4THYyCwu0xiM0ZHugB
nAP2QTXM0bqJKc97wmg8CQASxID5zF7AR7pLnX88heyCGCfJXa1hRKdIRAnYGgEG
gFbx3PV2qU6qQGOXX6F4PQZCAtGAdwTa6GCehhXiITb9ThZiBgSZqPKlVtU8RUi/
gac+6yRfHKXQL3zgfAZBAshKFxCqwt/6Ec3e7fdyghaDuVacK/3B1sodIVbFM2Us
4lZPF5shu0jtT8YlDcKV50cFjA+DDfpZWmHJfvS5z5k2t63CygLmn2iVTCzXM8mz
aa0FRn7OaTYGziDqT/vKWKZFVaw40YgKXsxDzUJUxC82tITjFWvgMUpu0yNStrYI
NiJruxqVRJj0Pk3qdu7fpbJC0OzrCWfie0pA8LegM4T6BimU+pZAjgWHiWMpiknn
3AkrY+ozfLoCTPBcUonp5ow8aXYgLZUtL4gDech2KKl3vTUHGsUYkhQ9+ng+/lmQ
C7cUWW6xhV4rX+FZNxqu/FEMl3E/fjg/0wXbDbvX039KvKF8R63iVJBrhS0JA531
V3jtgckwiUqa0JigRPuTH1R+AKtWLZi+E0GykGvqs7bKz89eJFPjTT6Lahp1tBz+
+7hBt05UhyDKLtt0qQgtXfGtjLjZC/c4e84WSqucxyUqqyQobcFnBC2avsxYCH0h
jFDHQ7u7JUdUwwpZBggbIWYul8Ee5WawHcPWS45rB6cdC8RNsPG7mZOmV1q04Bux
HyG818esS4Xpiosnd054W60BTKU2i4HI/O3mPzORFpufeAk5C0TT7VRtn0unZYhc
qrTydj2NqmIR+8aGX42poLoCc61rfjd/G3X+Ttcn0mSgbbzfybIguZzVMIZZqIo+
m8j545GvAX4XxHiCgOcArL+9nupe3p1ekE1w09yDJyNMkuxTjrtbua6r+8O73Q7U
+zEfsKci2HZD2s7H/o+dqMO40qfEiFNF1prycgAjOlmR8TPtXkiThYplfKO6VWTI
D+Styy4D6DKtSNlSUSwTY+VSU5P83upide7G7x7Kr1XZp0uSuE0elf2AIp+pe/hP
EHyt2cPMUdoLHxsqVfRqBilQXJQZLtIrIjqnsIamT5EUMFHp4Sb/eON+mRFdTL4+
EZ/kU9MSd5q82TcFdkD3aRYUPMcrEyGo31MWJBs3jJnlix35teSkix/P//Yh/8iZ
ytahfguWP5GtZ+l9iR2yr/aKuyiwWhReX/qFWJsESeL2dZqqD72ix2eJzOMJckS2
mq3jm9dcVYVBV5IeyqA9rqp0ndBekt19Mm6D0E46TfUGQwb3e3TD4oZtxx53KjOh
QhvoupC8RS+wgrX+c4ZtKRIqRzM5KrofTKnyX6WXfSDBl690qu0Ht5s6rEtrVnFq
h8Kpw1iQhMtlDeDkXG6+e6p93HM1JgMzv41iX6RlFI9V+MTSgVZ//19v2HD5ZMIE
kX8ik1eOw6goagbBewbB3IHRbJnKDjp3nd7yqBzGef+lkd0xHPwQmiY8HVCZ+ja4
l/cUPGR3mwOUGit9I9HKEKE2AWDVVtsX+ITDg43KMLmeTYj1hQtifyltK/GITwpp
ncZ+cNtBL0N4ZREAGwH6KH8a7yh13pDR1xoJlyAdMYvzXxLPU/2a4io3kaabEGtA
2uB2s6i3xrjduxXiLVhRLP6pMPzy0Cc//dpfDa4ETk6O5PilaJLDAt7qvxCHkGQf
6YOkCXzfOQMUNBE3OkcW0+Fz3Re6pN3Vxz2C3CeZab8YUmY0HRkdGCUAXVRew0za
iP+vCTDsVGh9ANbVhAwGSFUbPSPIyqNvoJ0bjx5eJp6PZMDSC1xancIKl3rV+7Ze
XtOxhx2n4KVvcsitFd6wy4C/2hRGV4w9Xn50K6rR2RhaF+pkLlBPSqLlnKApqKc3
+AvES65DKDTH+SHn++lafb4pazCRaO3/OjX09IOrV80WZ1TjGEH1TWwsnt0lclrb
MluHAImDb4UIqYw7LMJ1RiYXUKJnSaTuY1/1gMPoVBiypdhnxIlz2D82CDAcZQYJ
f4SOO0q2w9mkMAARSfmDrdpKrtLu/YVvcGy6c4p6sBiGKk4jQ7D7gyhPLwAZc6Zr
/hVNAMXMgYD+KrcrQJ5Y3nqmaMQTXlAIBy4Zbb5duKh2G5bbHzCMEIuqA4MRtdRb
bEg1xcZaw79yFiqFPIuhuZ1JQF+dCiSvzFb1Piiwnq68fTvRbbgI2V8u6T+XhY7I
4UJbqjNJII8pebYBxnLYJp7O1VrHFILTisWlmd2gv63sllyaT6lTRlMfHWoLbOyI
8thrRaWVd76t+anVJ6cr10ObCqJ/H/v8ByQkbGHvP9nElhU2/iZQK54c7Wca9/zT
qNa5iOT1b+QrHcOOP85rv+GUQYG9zKK/DItvPts76oD3OeNj0xSL7CxocmZVg9qo
3DQqBnTIB2ry6B3dghLmePiHJ/9zE0aouD7hPVgKZTlTm4CE4YRPEiSADLC+NsAY
ISrY5p62JMREPWI7FesU61AexLEm5bMeQ2Uzy+Q13fpnq/fLodWzoEOppjqtvCNj
/qqINyfyW+Qsv2zraJSo+7bYnh366w9iIThcVqiucoXw1WLV5u7pdRdM+8xsqfme
/AmzHOA17MnuyRoywZ5093uYkHrJAVSFjny9oq58Ov7uTeHUlckF72lNlRDgo2VZ
Gz1R1s1InOSe5CbaGleBra7XgPAGZgaOqU6Z7aVfsGahYLXARVN29bdFY4nAjQTC
rem9ZwrT3sVNfiuthtuyqTDKr30BXwVbuxg51qJgnhdCTwQqH7/XDEmkgnPNSUSK
PdtFZIX2pI2cuZQ8jWYswmrakpDjcb5/R7JA1B5ctqdYc/A/S1KeLBu+0BhQ0dbf
XIE28v8vZKzseTOsvTuQ709n7n4KuEdx1vXwd7JeUmvCDidPJtIARS73nZXN4SKW
Y3WWSMF8yt3EUB4s8mJ5b7rWwzQZt1/mpmCfw4Ssb4Yeq5VFG+Jrz4DuoGIFCTgt
RU5PekYnhlsZstktPqObZBgYzVt1BbJTvZHtpG//Gw5IIgdPV2Du8/AArMN6fqzR
Y1dGRHNoZcOJ3CyPwIzlmbfJVoVHk4uGfXYj0zhzpfXJfq7SctLXiAGCT7iEC7T/
RR3PXRzJA0ymxMwx5zxTUcGOpCeWFmaIDlLTmPnMi3ZpbqxL8ojkA9XauBN8dsA9
OH20xspLprd9WXAKp4PvLxsQeCGuH2VQZXph400gHYBqXoP7shkaYRBGHgukCe4/
3+vHMdtEVSco14A98LtdVkS6csO9ZiU9wQ5fMNj7xJm4+N0iT3x83VfnvIV9BNrM
8Y7DQoI+D09thVREpw5GrhvSUPSoWyArDUDbDSR5vTq9EVve+BHAwnf1WRhMW7oa
hi/RZN8YJTVq5bVrcQvbasAcaSGhHR/yYWlv5IiPQBI2NL608E9qL5YOwfZGi9/I
wEvjqZFYrdjeL4uBxg5IwXsJeV4M6xMHEgaLtuXU6kjabEOJr1s93EdMOhaNSgPO
zpY/Tjbpgu99V8S5K7XQTifL/fIMpDBe+GDp77GGRjvamBT9jOZXeMgrrmyZCiHD
ifFzCMcUrbF22HzNKA4kL2ebzJzUthHA8emr2GbMh37B8rY0O89BRqD+o5v/Wo0C
5yHVrryPUCRY9FFvYk34c0PY7bvomhZeU3a9Sf66RByBvERqdph4OUoL0LEe9DNM
eq58/LW/EuVcYHJcJzQ5uM5QRvrLthdhVlBh/t2VYnbAIPOCWTaERb5ot6DJ+fBV
VqMoPzbM1eeEkMVYilH7X7W7mFqM3OXjUF8J7Ky0cgSUnypapsxyb8gCuJ756tap
2JRKi/hq8L2oGdYN19VDrNGjMhq/QDc1zJrWef6DSXffTz6Eu2gyPuXIA9zUj81y
hxfwEu/Nrk5cGL6vCKXGueAxwCp6ezZoyDGjyR7LvHLtatNkPMqS5C+9diojVLnB
Iiiki9xQclTmL2RlNCTiMx+f5bzsAQbCtqattGFrVSXBZ2qxhE2WyuIIngl90twz
ZBzzXyiYVpAn82pfXKPbJ3BCFKrZnrL7Z9neH23VNmXQwJR1IsUAvWaashKJU74Y
60z9ToAWCWOH+1k20zVrrFEhfYL3mXxJ32ISqUzTvIa60qzGy88EVbX7wwvUKWx4
kybgFDMcVvPbYJ+6G8wFjxSKkaGa7hPhSzZ90ubvY2l51i0+AF0eGU2vUqLsL06i
wttQdr1UNZ1cDr6WboaqmQkHvKEHqTqWvaPKe84s/aw2LPTWQUnmCXpVFyAzyGlh
RXp4mcdmMnvxewDjzLnxBIKE7tQPORpQi2/sSOsrj49SSQLYhxhfz8JJH4rseDBe
7jFPbi7O+PTDWPL91xMaH+khJOa9BBFaya8TYIS1QwIfsxfnPFm6zFWLfvQR9Ul5
BPx4GOp8mNBQ1zvBZqVxLKLWLCRIRU0tWPrDQQ7jJhEknIjcze8CpUE8V9FIfG79
DAPC/r08czwY5bmpeLrNXP1cEZPLzB37by/voVanGcAzFrWS2oSbYN4NEJ4RvvuD
ZKxfpkATm7uP26b2TOgahzlTvLz60JigZXU2SphZ2L4XFsDHnmTqu7Gd39Vq2Kpv
MgmBplj0CwwroKJUzr9yt1S0e5uJMHiALg0ycWtJCz8ahhvrVTMGo47edeRhPpCQ
lhglg13UHbEea7uEVwbd2MGx37Fw0990ivGSHbZ71wHrXJYOqReIG5yhr6eS4UWq
/RLuDxtJD2l3B0RhXIzBcSv8Y+L6Ni/i6D+9tPTOtaBO3Mt7VOLwlxwUkSYUkdai
66XYiLLFEhYLq3XiUp3gJn1+rlwe2IT9BwlyVmglIYK+ZY94mqB+X0XRpKahZq0j
kXk9Iog+za6v7kYNZQFesF0420arWDdjZnOHEq0HkNO2LqVyu2CFp41uHyBH56+F
eVMgse8Xxx0Vojx7d8tTljG8ONjlRv0OUVbL2LO/w9LgTPcXIFE/n6oTGz2OCQKe
TLIC5eTqViVQsfXeh1hO3x3TV3Lc8r24vQt+yNDK54MAvKtPo/ghwuDHW2I2oDW9
Os9tIBw29OU9nx0SnMQsfFsqSctutQA/VqQe5HYuDvpk7luP6mUTD2RWSaF0DY70
rxL7CqKE1Zg3uYREOqloBcRuebR2B2kh4I5nkz3aG3IRcvc8GWMEXYFmVV3Pxcxm
3D99cwa4ykENxX/tZvKZICSz4K1M1CryA+i9xGoWD8htBc/I4o+PA5vnuD8lrBZG
9Mkehw3lnmls+1RtaODeYP7lQtrdLOdfLq3StBYuhGR9Hw9a67es1VanPYQXibk2
G5Gz9Q8QHxZ32NuzUcjufa/eALMV7zmsoBs9WMh91ZJwcIFQuUfLqBDihcsZGX3V
LodrfBN0eI0fxChfDJ2mxJJ6NT3ise41oMGvzvbVCD7R+OnZeOpYlwMKg7CRJ9ma
QUi8wP5gSKkM3fUC24MeXPFd5ydKzPr660beRjKfFfW9NjI9TPx7a2reDmvidBS4
gq3g58i74Kfs8tJNb5IoXpsxbk0MvR4Vyq6NbdyN9mDSMUl1tiIQsjflpHNsD5ZD
cPnK+VRvfz+g91i2SjpPmqy4vimRQsSZtkrdeMURT9dEIT1WGTZsSCcbNkWwSCUH
NnirXmgmkxCg08mqfl8OvdZNLrCJLdYLcxuzAHC9xZ9zJxhqPolblDokD7ixQY/c
Y52Y92GrX3mE+C88zlkyCyEDqgv54oNNKNqfLoj/eivYQIIvvX6Mge7ozMfyvj+Q
jDRr5mgnHrliMT3m5UxQsqzb5mklz4mwguHVrAAyN9Dv4RfoCxnYkK/JGcC5vaTI
FlCY9PDZf6HGyqiRB/u+BaEOEP5aOPdlihKVDqn2UqO8LaR4awMlDJjeJ18EekCV
t+RKFOUKXFUgo+UZgIamsdsltPUPUtspFVF2eAeFORKbWUmQhhzYJ1vscq63F1Ao
ZYwlNsveUER4wKQ82xVeOFqNh8NbsxErN0W63rH8KOTBJ8H3sBFuQ+gz6LuoRHGI
KxHTZA891ub/3972VE/PHjUjM6r3SUqQ3EhpndXZMxlHJcm92S1WcuIk5CmB4evn
6waItpQRb1E5FTLZodUixIczTRQQvjroLyVHMiSfbbLAMJJZpW/mKA6lq1pE9+de
kHc1o1e8TPywfU+YgVP06V9HZH7yAtLn0UR1JmggwxqAY1md0cLNr873dnRfjEcU
VxAOB/BQgppF/G1D4blLlwBzt9u5t+k6mDY7B93RZYx3rmhejS5WGjla33QcBfG2
RxV2j3jlIYFp2k0Poab0to8AZueBC9s2BaP2+lczGpGAVDi37mQ0CUqodA9+n56G
JWM2iLJL0kYkO/faDD1Mc1rnUM1jv5TyahHFWO5ThqP9wGuwgaYg2vxT52Rz3qS7
sEYIZYAQVVX401AMcdwZVVWf9RPeuCIxq/c/tPh+nuHBWoMLDyqIkDfLvF7lDwT2
00NHJahL1W83XYLhUz4rSF29WMZBv8wpS/pLI8TZ6GUpAIJlG7Wdjyo2hP4rzPpi
RSqT+MxtCOHbRl8d3dvBnSK3OSkEz2zPi3drSsQq0iiY+XBFkUdAY3h6a9bBd6w9
3OsjDBaoGJaydLDMc/I/ERD3jHHBUkN2JWcwO5Qvn+nlVSvINqPE0hlTXmBYJP1c
eKJD2yFwOl8aLQQIyzTFbRybKTumSZAbQx7mJx9+14xrP8EnI+oCSaF7aaGEi/MV
PMTK1+xn389ge4kYnHyHOwiHQ90hdto0nQG6BZ5Cxfe/HwnqjFL2ER8FMwEss6BO
8dMrPhgxe6X8B7qaEI97/GUuv7c5YPGfc4C3MIg3Smpjjda4gPTdMgtg6jipkw1q
iR6mjUsL5JbbZ8iCHN81b6+HgXTOFYGL6eA4Rq0nNwgEWkQEvM4jjasPCSuA2sv0
w+tHC8oDK6/Y5ZrzJdS/YXDtMl1Jm3aZ+8zPfbrdvQOKpoWUp05blPuQHomu+5/t
hnYWj1XtFoadSFoFc0hP2/2Q4JdF0DJGx3/3OFgXz3wP9802fQHwzf44806a5nuC
6vmzSUX1vpgfLWxtuTl6hWGYGRUcDP2LBJvtRz5z2TUr3J/8VLWLPHWw5P4CtmU2
3PQ+7Hl/NRDwgMqZmFCN75QryCOJBhg1RLSeMZpOMBQ8wt3h2Z18Fmn/FWybirrz
IdIj+/MD6bXdlbznEbgUhjB+aoZD5Jr3JcARxp29zJsQVuQu7Rvhmuz64rNZCWf3
/JbEGHu+14NzIjQWzzicRsg1Vbu6SCvkKFJ30qHDE9Tk51s/7Jx4jgJIRWgZXba4
BZiI7SdkLjghyUb1BzV47UuGGbwQuBKwtPl0s7Hm1e8acmbialLsTSWw33rRqGYE
t2j38I+ru7ceXek1pG62bN1IA8hEHPcLUvQtgc7JaTEGaHtu8Jl2R+MVkAmGIfQP
m2RxcsauGxTbdswdbhgD2Us61SCRtH9RFZ/tbaHyIQfmBE1D+xpo4xXgp7us8WmJ
MQHGYXjzpMRnIuBjHRzVvfAwphTuHuoe/NRheXz6YrslKfmvraThb5rzrRH9AQi8
ijjb3vNqrTKnx645w1QT3eerML//WgOPZWYetowehYKCN3+67YiKo/NqA3Sy70Wl
b0A1t/zIrCcgamLKb0PCG3uOCBEmKLVVkRIf4XGR15H8Bf4S3riroFBZvHiTa2P/
3C6wRla+lfd5KQcYhTqBKQVm942Br5IKNj7DbuoN7tOgV6mBfAnnjStT8vJME9zb
LYbqzVnQ8h6NyeeTjTbttgj/H8PecjIafqcjRc5PNGH0O1owS6mx9LxuKsfrUB4X
HEL9QBsWO0omJKH8trmDfc+U+B9ROOsWChglDNLHDl14qWuI2VlporyY3DfaXstW
v95VsZi3B+/Qe6735EQYCcMuS7rv+1C1D7H6o5CpOry7QleelXoInsvvKFIhJBdc
6DEQ2NvNEc+MCo1bfUBYNoRfNQMsO6irA7p8RHHBSLzGg78vld7SScff3DnJdQrz
75peN8P7nxxsLCHQkkvZeQssSFXqZep1DoeGjv9uLjsqIqQo5TjY6KY0rgUkI8KY
M0eSCCAFg2tV+wy3E/sBrELq54vpEtlnYHKdRF6CvrGtjuMAVjPvqXu05qzePoxp
6/Say1LRkFD+h/kgkHjuYs2lNxvTQYasV5eBUaZJRXIobzXOIx1NnMTcXvts/lid
hqLizPGdf25cOOMMaDILggA5sunUbngMggQ87pyONzORhCKaWwowkmjDEi5nW+tF
5BDZf1k6euxLEN2lNLf8629QvfYgmuPJfOb6EuoOCUhHb+oQyWK2I5r15w1pibZE
JtukfRsWwZKPWH79/GOE1MBB+IJhV1CVX97tAUJkIwBpgE1KyhiYGkDZS6iaftUN
OMuHHlm+yUdySGR4mc+tH8NwT4WB4pKf3SvN0/3jG6Yl8Y3eqH1HNzBVqEdZHQCh
ankNRi07+XTvGj8o703iJiwKZMQuzI1CLEteaELcKenQxXpQEhnSWhcE5dHbKUiY
pRxY/ZVXH1f863YZrAESIGKOI4FKYVmK64xSiXDDeYyvxUX+wrAEh23vfPd9qoXO
3PdXp93rmLT9SiSMUCVp3UPxX0h7OjNn5LdBMnZsC1q+I6zUJWXPskQzt0OHx0RA
JLFZ6MQJr6bR0AV1jpxHXO22EhpOQJ0u7eNjPFeWvW9gOIDi0e8iOqYJqz+fknBJ
immoBxvb1/ujynbh4B2tcw+6Gh9O8oV5oywhtVyb4dRMTU8NDP3zdO9boJT9bNl4
WJ7rhSbWewQJrn8yjqsvA87WQdfqZBypXvFe4XxmH0ifevbNXH13CFfAksqEbnGi
csUAcvaStTRwum1geMxMyINaWP0QnieXVQpJJ7JoAKVVz2/ozHRE4Mr+bOdIZoZE
/ZH5j8LGCMRL49ooZdzXB0kWP9HaJ/JTlb9VZpM1KFZb0/IJWgS1sm9WuDp41j+j
I+plg+IL7i8tkTMDSZxV2tr3ZAstl2VQ+8Qo9fkFEuFfyKQZ7gdDXZ6eA9OoWSe5
f4nV4TKE2hRsvgNRqsDVbjwqtErZSWkkJuod5wDpW+qnljk6POpReZHTho6NWAvS
lyua7ZPW88FtiT5x9xRrBenpslIyz5mI8s73Yki8DZiwAq2IuAP4VX41OLpwuG4C
K/3anEk3Ei4cDSFqxbEvwbKZ3O61mFlbwq+ydqQX+p4DDhObdH9BKDb5mtqKkKLq
3/dzYEi8Zk++VbYycXWqMzuNwE+ZPmkWKj5zcKNDjJ1UkJl+wx/kXeL55TM5EEot
tKzROuGGShmk9k5fwzD5PUynWvm/8+mAQLnKcS4wKIS2HFbjPOgyxvTaqbg881dn
c7RBUWHw0azn7ZrhNEVQ782uKRvl84i2f3GOHqkkGFc+haO30Ha82zooO6x/nZRm
132NVHFJze5DnKJQJdOby/66vqfoJaKYnhHRyo6GFAXvJVU+03WYSvxl5ELxf2pU
WnrJfCP/HLcr9mMWH2Gbea9FeKaME1lTyop5+0joRzxN+s+rY2GdWWBqhJB7Nf+Y
1T8HKJP7YtN5tjZlr7Tr7OYqsr5KvjooteFtQy36jL6v0G5E4zQDyaX+PKMpMzQU
uE8Qa9xeXHP8u3iLFUfSCnhMcAkKek/P5NYmEjAoNEfP8z14h9aCzqUyHV+wb3Le
+w8IfDI9nzXiE2LkNiKbK82I4yicggTphiDOEmwLYHR1l0WKLLtQQaJU/bIQVByy
W885F7S8r7z4l5/lz5gdXlpjDqPjrRAY0MgZCqFZQZr2clCDm9An21/atnYJ/q7l
WDbjVugzb8o4EV9IKpnytGYxgbueElDpWNjAvI+02YIkU6yUya9Zpa5es0Et70Px
nr1dwmn9od/749kO/b2xEq18NB3RqLJd6gsK8nUmTLNAd7y8jBbEx4Kjufvmw1T9
LuyqwlO4ACrzQCSC6DA8N/z8PmDJpvoRnrj/tIDHMO/vZsff/tBax6IsC4gK2IRL
glKJc5UVYg95vbU/czDrvMv+shXfc2UrpbKJhHbFh6XrtnqgVTPRLmFySkXfEF2l
wdDPdkAJESbAzjGjOdgqe4sZN7BXZT8SZcK2234i3k4Pzk5eN7bavfFeYg4ecOLP
nvkYzpHc6nESzVVF1OA0oPWki93nwOFblfZZerbPmtDnHY4wmWosfr5krzBxAuHa
UoMSqAVPLvIh2Xl9PnLSbAKzAeNhf09YS/Z+sKt+9BeEp8KoAztPCMjx9S+InOkD
7D46sjv4W34mmDOc9n4Udhhw7VJQTrfLSp1SWFm9W540NTv+JFehfxarZIzwXjEJ
wTJ1JmCqdisIDZEg07GBo/r9O5ihSm20A8xo+Dvs5+TsmjJ1SCsN9b+pDGHyXiLH
4SuEOaT3ORARFwS/cedTx2e2FNOTA6HpYdVk/b5LrjICVxRWYaOtIT4Lb0bbV+T0
R5hSSPzTJ4cjK24TSjLVcnwoxQ3q9s2YPZicPucBxPEUWwkkaGyId5tB/awtXxT8
cryVEYQGwMy0yRmeO9NbMym/4yVbqu7g+r9sfbol/UqeIoqd3ZCOFHZ/Rv0ZBYc5
TWT31Hq9VaZCiNweEd3nsCEKvr1nsv2nRWgQYHNVtuURuW+IX8yNUjDbMN7FOeD9
3NHPZS+TMSll4ePhLb1Fsu1sk1IbWLVgts2aPCiQgEAmlRYYkCGzVlQL0fJJNllG
qB6P8WY5oayJHYy8avrW5YLAebFRZCuq7VsBQELfP5QafH5JGuLVfEefare+wsKc
Gw7Oun5BK1VBOJlJuO6vnA2A6OgAKkwYymTOrBcpm/PVEhFNuo6k+CnEttxNgXN3
fnB7qqXx1z+F4u07LWexcZAlur9Gpb4LcngtkYCDtUd0hInKf9CszvoLcAjcrQvO
3RmAgq+w5H+23Hp0hQuj3iVZerJOxNswhQEhIGlJ77ukg5P9Yb3ZqlI7Se+h6ZWM
C8EvXvgEkK+7QKnEkvEUkO36eAhGf4/jAthxIQC9Lp4AiVklRDbQGJ6brnpm0cQS
Es0YxfEGspWugFela+B5ip2gdVQbRirWC5yipmFQjIThapr6qNnmWCTxjqiGB+wR
DEjBaEin8iNlVgvc6/lsQNMhawcvEKRlWYUTd17UsYStb15YMFQn7BiHO8vEH8ys
qO3yubC0c4OWt5OkN0PruISmrbv9Bnls9f1lni+zvixYt84e93cGdHgUKjLnBgNq
/hk7Uz13y5uiEn+lDeXqCg6oO0+LhB/Uyg/+Dxpra4cHC+bXB7jywOmvYpkGOm0e
gQ+zzb0L9gc2go+OST4cftIYgUTa/g75Dfo3OUTKjODQ/WpVVQbSgRIUyFJaKKnA
x0dCboAYpCQPThL5stxzJUYXgEjJhfazvI1n165mkuSLmowxra3lcgs2hsREqfor
e4IL8FVJaz+0bKO8+PXLhsXj07B5zgxRJqn9Q9VsNABpN/U9nk0DWBAAD5vHCZ8c
BfyTPN2n2PeT49S/Amwy4LmL/fBW0sMmKF7sKXRyuFE9DLy8mjhyMexWJkJxItGy
QAMp0rBqPfE/GPGGKQy9zvLvs4/8T08Wct/dGMeiOSIcPPqe/t6lqIoEgPZ/O7JT
HJNFVWl436JwIOxyv24WR7TENP8L3ESZKXUdBO534OUtJ+a3KsUumH+3Yf6nqEkG
yeMkILL3xnYSIATQz+qjSeMf8pPixlxpu+6ovDOKem8wXWQH7pYUD6S39Wk4fQ0U
HBpy8dP2ujC5v7HqReKqfAXE/pAP1kfQSQznP1rBsJcIYtVRZ4n2p9M4zNX8jnB5
r0dZnbkwqVi+8dw39hMabQV4cyMMir0mOElizAxDmUx86IPAKZgJD/aiUSjMzFJv
0GKjicW+Ij/5X1c6brDccwgIldv9LWvcnYicLGNxWVayt/D5/Wnp5eQ7p8SM3nIL
imkH3z7HaPa4LOG5kYNqvGG3GRI+9Ybfr6hag9DUDgIlWHVMNChjO2450DXHZ8DJ
FbC2XGTeAY6aCrwHKSwU5GFXu7zqP0sEbErhIC5qPzrcuPP6ZcGYohBYtXJLaoqD
xzeevOhcM7iUTH7TunHTrrdGfQIWxXsIQAB7Zzw+7TaKoxEI1sDWi6Q1Dr5FrSND
qMK+GJrb5aBjP/AaZ6HCvxjck1XrdrtL2iEtIwHx0wfSNLG487gk8JDYZFbyxeiU
0+BN9Y1YFYZ2kVFP3HANoa4xuMXozxZPh2dC5/WHpBgBSZjyzp8DFXgSwSz94IfP
Pi3pBY8YZYhpIDFsbUs/ii3b9H5CKCBwMt0CaCjzZZh89RA6avoEleIMQNzu1Unl
EAvpNH2VluhP/krtaCXNxCTwvpvvzoaE9aEnf+RQWY+5bzFeX0ZP4PSaA4Xc10cW
0MLi921Du6JEp6sryzqb9NAvt3NF8XMOXBo1LrzZkqllWFR/66gvZG+8fKNVHl2y
gVVhz/A24CdRdmBdWJgu8EBSbuctsP8kPWrCPGzYhUN2xpHNtx+d4tAnIrtJ/owf
a24quH3YxK/XrfFe6LoNoVWViQ61Lrpji7PVKy0VPH18Cn88e9YEbsIoUrGxc0mT
GhCBbmqczr1Xengv80RmCRgy3mGnhHmBfVF+KIRq/3HzRUeaCS5ug9wy14TU7MhX
3by1rZVnHti87Skmmvq/DmkXImPve6lRFP6CkJvquW+wfSoKjk63HizOnlxgUPlM
wK4uA5Vmy0qq3JfG9A6kvTXUW6BQry27AgPsQ1EyVYtgt1Ko0J7PXpDkJzDBYdSR
BboIfQCE3ho4Kc2BO2f72EgMh/P7thVLim69qpfy8Q6Upahbkp6Vv11EQb4l2E3x
ymUQU2QOLE1iiYwjhgGXrxi48MisdqeG5ILDZ62RxYgtzq+PzzX+a5ltGYJFjoA3
l7P1Nfjhog80vF+T2WjJsANugixyxoeIN4uaxoLYk23UOPo5ZgvbonTREyYxkBbG
wY6scPmBQviLbT9LBrQoo940+2YVKqYwVIvBCBmi1rWwKmeHQyPWx9nk8Wd+81G6
aI+mYo4F4UVW0w7WiLMwrvI0zj1pgkc2F8dlSIwx0bbINrhU610fKdvJ9EyJ6u7E
iRE2vwkCksRXqje8PqiJZdDoUvtRAsoVpDDTLUXCy2iPACH9zpH0VkyqYxnF6L6B
CAVO01UqvYsFJO61qdP3aqpbdPJEkua6M/e8yzhc+F38FRBWIn7k6Pn/uGd71GeM
yOICgOduMNbutiVDEaFKGOwSiVm1+pI1+9zvCfLmKXwr0Sj6T/R1hBk7qv/4Bw8C
JzSaJ1T5Xz0xA+tQhMw1M7BooU1Nro54VKSOVMs0BawoVydJli6FEfSCZaLZhxEX
hs/0JzYEMAJ5yaBtkXKWZcR5qnWMIT23v3UEhijiK8DEF0pmP4vM0kR3vbyVnXm+
J3NVlJ4nTAjGuiCuh78e0hXAFOnRG+mMWPrseKT5DINuHp5choGxkdZWdZYoNjLl
02N5hovdMiBOJ4Cly72PnrDdCKjKttSP75yGfMazztVDwynkRxIGBvqyY2vNI9LP
Qg5+8jtevLsJ71uKJf0Zhj6JZoSxIxyOWDAwmMS8/Caeo9tY7iuBnPLuDBSG1Kwt
4b1oKEhTcCbTnycjHQmc07ocNJ/oR+/t4/BN+a3Ph6+itBEPsq5ew1rkwDhva+K/
eUsaTKDf9ZaJJBNIA+9mbdcigs5+aE7skbNoH/ToSfPFqwg6khSesoqVv0mqSNyh
VPCPUxJ84gc7L2pwVF5kgTij6xb6a9U9VIBOzWQO+DwhHwZiawxgx0f3vxJrr7K5
4dPfoXTFXQYefWZtOI9c90A7SVrZpsu/W8Dwo6Ftuir0Ry27YaOWiJQvxN9UqTNE
f0lCQG6rOV2II9/aYZ5tbZ+04GFKksEhs371dJCDIuo9DEieMVhPicVRHRi2zvCH
/A9pabFoA+i+ekLZRXwyARUpnBQyGn9sCzL55kFsScQtPi9cynhOy4C+gGF5PcUM
bMTxcDieY8xbqNPMeRHKEVJ4UhgOgu5S5cE4+qyXONM05ybS9jUXzE+4bvY5OtB1
Ekccv9Eu8z33HutmLyV6ZTgdp+Qmjr9EPuTpZBc9If/MJywyO7klCCr7HVEc5NQK
YQMIt1m6b/gC0cytr6tYcSzH+GK4l5+7XQqBzeoux2iPt2xNA/vcPKRAtNnWvExL
evdMU+FZohYMTlQD5xF7DOuNEoqfmsXETbqspWXsiiHen0E5bzDfB1F5rhbhs4jm
XUfhhiGPEr2q0aePAuhpzX2P6p/7AUQkBdCcSuULaN+Rl6JyuGmSYpREfJ3264Jq
BI5+ZkVsZ/x7le/NyaUte9mJ0fgkv3/umIBslvuEGgu4tK1nQuvTqanyJUo6XR5v
EscgimtXMG2Wv937ga4qBKSnCxYrDPupRNCwBA6z1WUkyjt9/3CThebnC6pbsRTZ
ig3JiqlocOasu2Wf1p8KoVFv7SjSEI2DGp7z5UYJJOv2+26EpgDSdN5B925+OnmD
WUHvob+YfbacKkHQDwlVkYFoup2URNXR4YyBKMcftmDnRc2yMFQu+nWVlYR81CqC
GGVeeDovu0SGyXUsmpgbDJgfn3F3ZCB1B3ezizimiW/prbnXeoMin2dZ51vkH8Rp
zQ3T70HDQOELLl8tiCw3/16zcNPidJgrTzkbCCyDPfr7rLsjdgvY16rE419kcleC
dE572zQLzUtkEZdhOihrSF0HWCjLCykVdotMiYi+mvFnRUXod7K2/9HXoYxxxyny
KepocQnweeskAxa/lKKfGsfm+Bbi8C0hQiBU54+Ed4fVCAwGrKvzzDD0g8uSJ772
a+EbULr3NuoB7ekHBNfGIhnah80lAPkyTITow8Hqn/+OttvnJHvwfA17Ju3Gd4ng
yoapsLzWHBJt2vCXe7UKFRykkIQ7sKR5UMbtStswgxrQN40g0/hmv2znVkdRiGvp
AyntmbT1AfcuqYF1ro0LYvzAnk620NbBbKxr3diP4y1sBDj7pGvau4oqePRnoGtl
mwrpzQIgK1CYa73vQqnBiPFxV5BrJPZL4u+zMFNjYZtsscFPR8CEjOvnAhfYdw6f
wfSQKoFkxbmdjvX9nym9BMTI7avxrfFzBXDswHuA9QYIevmB1adP72mRfIvi6ch8
sAycP+aUpb3zMs3cCDSU0CWuOJTpAi1D08vTU5prC+JYlHaV8fQAc73OdY5kO4gA
SuSEk2H9jMknwDvELMc3bGI1s4mmP2Z7ZjBDblza/6ksvunZcNZ/ssMv1evsnfjP
eh3pmvhGdLiYhgig+xt/HkbWqLIxaIun+9DcIBFR+1jfH4FXkUp/1k8n6XamCt9V
fimY2QPvXlG9O6WQKHIAFl6XqxdUz69kfEZQpgVdasnteSsrkXDV1Z5Kv7AKKEa6
SfspUdqEwB9IGhEe7LdtAE2i8RlZz5E95j24k2AKHfhiD6CiVeYPHj9t0lo6D316
n0YKjHLLJvFEd+fX8co5JtaLpemy3jg+m+EGari6Q9OgbakgxNxEYe8S1qQy/f32
MvPuOZX/AbW5rc7X5eWvzXLbMjK+cx//p2qt0pCjy1eNSJA2odHP8rjcILBpUu5M
A1fh+00RIDgph1rA3nefcXDWbtqN0VZIPJmVwqXT809QIThbY0K3NvfTDpaSp9zi
8dWFi9+soZMd5ORozCNBHKkR85nOUq7exWXHN/gfMqA0m6yvNU8K8S33O3sqy0q1
uHaPBTRQQGQqpwJGKElFItZctyQAy/iWFNzPVBGaa08sciOROV73XXv8yS0gdDFt
Qo/msn4RcJwqNPHdfNGzV89hULN0hSYe2runVE4h3s51IvHEOvoOP9fJTaiUduNp
o340DivP3SryHOaZL+lNPJEvRTx2WylgNUEC7PgnpGd6in/iMZosQN+iPklzlViy
DEvFoTOpA+po4XZpEf3fP6ZscAx9JXfMn+g5BSjcFhA+WEnBa1ga+GYCp1G1/HN0
7FYha7+Yygi38TXx+Q9LX6UVscotrBiw0+AA17OFJwOVyAInlQPfJk6woV1O4QJS
mROlK/hbn7KWwGj3PQETy1Y1+YW2E/e8tbq9VDrORiwfRiN7khTGrIcHr6QXl2Ww
iEtd+O+49hmnbs+jlL909fMQMS+uUfTuCKTgw7ffZouJNQcmXjHEPzJQIc0x3Pcp
ZQTBhBXX8st+iH9i1ns6VRDfYonEi3Tp0QqFuiOzfv1jfhExOVnSLXr5KnwNjEyA
mkf/DKR/ivyc25uNcTeEJx7NSFurE201hOcyjkvunbFToolFhzT0TPFjWVv8j1Vt
0NNXgxW44Uohjled18N+mT2O8rX9IZd3xhpW0wsDy7+hUqF/tBkL63SWhyO/a4Bj
bjtXxJnitKH6zFyn1mb0xX9EDQAJNTqDdnDf0tFqMPA62ug2nPj9oogaWcss71eY
VFy3XtzzB7WuInMXjRC+Rj+LVzkdQhPFiPHbbgj3DQt3c0MgE3W4KRsWMRvpEAua
7ZTBfGrm1VIfS3877doZFT7QuRA++uqA4Y2lUggqSOmKXX6x9mtuFUOrZhcWGuSo
bIuRS0fIl3mOCV1XQD6cMNmgBfmOvIxo9dBJeGm9k2zsfQwd7VloSXP4gKByP4W8
POXR4o5nLOiBp/onP3zXSzoik1gZtDX/ddoq+R8pO0zD+Ss5/l4ZG2hassSuzxb0
nWtfzAWrEYVqKaJuKpadKiBB3aFZHMZORXEqo+uA4HlIuRZijndXRCtTDbF7ZUbV
+ZEBCxoc54tdpyAPy2tjOUoka8M4sjX+wNYHKsDMph3JQ/WQbOUxxSC8S++gkVIo
ekzajnb5U5vn6xCWXy23wUnI0AZnuEB6iIvuzKooDevlAZb6/XSOzrlbHfxjjzPE
y8j2fbFoUrvNVjy3mRkc400LZtWvjaKNqqRxiEySfaEcNPT1FC9fV+/oHmKdcNXf
Rw0hsPlUgn11q7W/KcyWwvpkKcdRYWyZnSmP2F5w5KeQsOxLOLLwhEO9+KL+dxG7
ixYwPMpkOYIpf8QxB7rxyjcoLKEkPXPuUWuv4Wd8RmdAEjpoVNy+aRiDTan6MJ2Q
1e4mKqEpOzIwXgEzM2D0LTHNGLjQTQTsmFim8f5bSLrWAA0M0MHOy99daXto1NZe
TacoAHS8RxLhBjjkXm6+7D2BhqIAUGNiLQo/L6m3IgKYq4FKf1NsFNDEx5w+C6qI
yKljYvtnkciVZjm2H5VdtctT951krrYxk7wvOx3vFya6Mj3iKzyANiD+fZZDyNaI
ZdD4mfWJWd721IzyMhE86bU3A07yfkJuJWyQQdgxE6vJefhBCPTN+c5+ImOi9/PX
jsBD8Rkz25hO8puKO7F5jAIn4qGxjiyIwRzQaat+NlpLHM4emVHqsHU9LgyPS8Jj
WnpFfmwu80LYvAcx3HOGiehqmhj33I1/RpAiXot4XgO2KJScp0qZyI+kQPX3Bhty
UakC5mPs7tQFubT2Y2LB3IXWxeqKhSxeCV6/AYmpy0qyfPI2Jso3zrmuAk9hnhDE
TupJzdqzIkiKEi3mvdxaY1OxjQtb9SWUTUqLY328HqtTvjels2R9Ha4Ku20jvAVh
mYOt3HrcDCIGQSeEM1DsRCpH58vnVSL+Jlhy/fYJdDdQn1LtGazgbBlUCfpTmIws
/URAqsQ1J/o1fr2PTBCkjDOPoMATZcQWFhC/YA8/CY4U6sD61QnP/N1PE1As33nb
eIgH4w4F9jKzMnGyrVBtkShSafU4tbprGpKkApVP5P0fe23efR6i7JfjPWVZn4i8
+Iw2BMqFuPSWoKSYWxtxXDlSEQKewRX+EHk4+6VP5dWif9qiljhwA2R2G7wBy4PB
H4HoA68yvIgQGk/VMw3a2UEgb8bEfrTtkgWRf+iCEklk102Xssvt7ACcIVZmF2bd
bu5gFNHAvHzijzvCWyGnu1bHozIdx9viZieLU+D06kc3ubyuEI1gOOAmbZtUxYD9
nOdM7C9dXWkbQmw3TYWO/QXifOOpnonJh4R27WS6uRlHdpfcKT12Miu+9mDT17oh
FhiYWGhfiPZlksm3LWt3e60nEKoH4BJ1ihvAYXrkZ4W1nEltwE/ImQHfSGDfKMLf
SwlbPxE0pRM39o1l6iZpT9inRFviEfwj/b404x7ivjw2SYO1/3EWm2BH8lZbvB2H
qfiddiab8deyUHj6gBV9UuEWuim9ZEJ9aguFLsMXXEw+6QacF3MxmEIADdciENPz
kA9MzrXS+KNHyv+xgzOns/r0LyXSlDe88hsnV5PBTm9L826E2LwNoQ+PGusxUaFs
8cb65NFKTBkkojTNDd8of/0qFRcKWfMj6vaJPZL6bk9yHAPdEhv621FAtdgPGIPH
OSRYojLvhUIswC62U+OgPB8s4x4sh1xJfRwee1pq6mQGng1AOCFjaK8ZR07bNyPP
dgiFRq8y9LGrrfgGifFkLVBqQUJRUnpA5rrtBY2wGfXmXC7AWGXd4N14uK6zKHVl
MxB/kwEKrZf+ghceZKLejbBPQ1d6JzpvrHRiUadA/DyHjjHRGv8nnlAv5HIzI36R
SPxnVB68w47bRDZH5T8lXyR2xq36vw5CsO+9SS8wEjqAQP97FfTTQMJ4wR7w8yiG
T5elWXgLi+eX8/VpXM8zmunPKUlTZjMI2wHnBkkblGgMD/gEUfKZQCCqBMb6xa1i
viSj6LTuRSH5h0T2u+3gpz0qwW+m9Q+kWGTuUT9m0KjUB6aj9yBIWrqpd8xhfOuW
MCbqPoikW2iKwBKyF/R6fHtdch+dD7H4Rt+h0FuMSLDtl/QHswrQIxQgkJxxtH/t
2UoRBns6OWZZpI0pz0ngaN0jKrvAFPvfwO9QzWxs66DzRdiwMzEvZCZiBP6j8hyC
sh+FPT7odB+o3tWsxnjVppZXcp9GIFaKvt6pMBfxIS/MhIh6zbI83BuZYBND6RYt
iZP/UGdHu8OE8XhyGx/YYzPVCQTBk7+9fElB2Q2Q5o5wyvGfcnD1Xk10iqVndrOX
vRaFCL3W8M0YcOUt55AzWQ0kpDILtmtjbQm83gYv1+JNx3JInALFLEJmzzXWlrwP
g9emMMboFJCgN/yOYLbbPunA1ESaITk1gVGbPQYh8LrKywhfA11E5RST1BFHJGn6
lVisP/V1PYk2a4920XR+jaHlXFwxBOvVl9ayL9OKe3niGbu+CUWRGXhAfSiFmVnq
wiqVlPBqYeDcLSg3NookDcpTYVklw77H2hmzl04kFkB1T6j5hAXTam4XDtJ/ZRJt
Rc/tRcjRT7q3ZxQYmoxEBTLTrCFPc+iPXBgaY41F8wLB+yPnaFYRJiRBFZx3EZ5N
uHL/zxLECFot7S4LS6cGzJheFqgnWtggEPDkeeFmH1TLSgs/XcQGsDqm7jRYo6VB
SSw+zCw/5rcH2QHA1ON1knNKqafgDY/kRaED6cCoha+2OvlYtkClAyFd2S+y2Tc/
lATrZE/H5iUSDwLD20Y0zyLnnO4U6Ge0s2hWzgsICJhO7RAwWGwCEGi1xkj0Qy8L
0eUcnWGgFOGHIaJT9UR9ZJ/QyY+nLFZHfCI66kYgIBIBOC9r5I8qT54Zul1iTFza
XumcEo+Dp7d6u5EO2e163T7st0u9rTjwlELGSTu3fcIj0R98nxQiSM9K2MGk0vdH
CdTAIVn1T8eJ1KajB3VsnxxTuh4myJSpFyTE6t8sJTKTASbJi6ZmQ5NMc0aHRHXf
HJxn231V619sWhPdXSKodt7z5ybuYpmySViBdsvpMmstcy9Bbokde8WGV6Dzm2VE
MiXnJgs5fEaq2zxncnKtx9npwPnpvwfu2NcaQ/q+DW3yyltYer3oxJwurPicQ/Zv
h3zlphoOQP/JzMxVJXhYE79nJiI/dUmJMcY8yC16WLIoitfUXzrerbCd7EHjic82
ky/p8E4zAerARuwvZuKiLMK5lNyhw16ES/kQ7snI7PbsUrCVXylJCjwlt0Y95il7
ZpZygQDwTcEP1ZS2HEnHHtN/yqFr68nsRdxucY5XLyoxXQQN3KtBzixJ5+/dgY6m
2qvc9p4nUgwBODIfzHtIt5kBsgjCe0hbLMdhOHbod9lf7PDADHrT2ZoMOmQ86nw0
kwdb2z6cbDMkioEofT/qkmoWGy07bu4oLxed6ZSveZ0RvVL1tMMaWGOm8EItSs4A
VnuX9rCwjsNv+eoXMZOVG7IkgLPdce1E5gv9YioFa/mGTWJHQt8ILTRpn3oJubHQ
70qqZW3p+ci0aHa/A6/POEBe7Rznu6ie0QogPR6NVcupEurhWspHC99PvQeqroOY
jaxWQKLD0UaAuO0rK3YKS1WKErxP8NP/8DXXdLHYm7uyy5IwYd2rXAcIt3/rVkkt
ayA9ttxX4eqTX0i031qLoEuc88qwdmYPUe+5VF1aw3KPVFWUOu7Rsx1FZ5HMuwlR
BB/LNjb1sVwLToiBiHvxIwR6Qn4ZtFjLHpN2HTv7P2Gq3Das6WN6ECdNHJsyDNpE
xcfujaFV3hsO+m80uG4yknjVnBAmGwbRspFHRi5e+BH5AebC5uPx7pLelueuPiSW
L+GmEHhWf1AgaLxtM4VSLnk1JUi37YdPPQqO8GbSoPaGjsKy82RiXXM5tfmW+fN3
mFQAHu40EQXi9vZrqOCIV5TKvPg4G6wOG1aaZeKhK3lunUFxlaB/RDgCVAchFTnR
6+zDm02ENOEk+GcOiGtL/iaXTugR4alcbHUOkXJy1X56n6aX0JFLan7pJ9Dw4ep5
4zWMqYisqbwA5pkX1UDzYshr1gNuuDCzF7UgLXSKBltAo/6m6ZdH+T5gNno6jtre
NWsM1g77kMx7Qz+F/8CkUauR9ikx1FF9+lNpM83C1A2O8LEgwnWb5YYU7+FpH9Np
/QLLz/0QJImMgGlx1mANNDEJ9hVuvgL73vKrRKzIg6EF8PVUuOh+TfHf/dRQ38s4
f0YN1kcUtuzNYKYvcekoYLwu7oK5mmS2/CZYIWq73wtPc3MrzimrP31El1BINqcu
JP9jWe1LcDQTdl0gW+LsPeFB/5M7PMq+vp4FIL2VxaRo4cZVSVYxyela8i0Xs4me
We4NO/PCxtSQnajBd0ziegde8asfWZcqnVJASgjl9MuaRcLpBTN25DKKnFLTGnTU
qTe4Qtiwxp2pin+IpMi4/7FcZcyI9aVnib2ZaBQdlW5OLXf0IINNtUjXgQgnkL8r
mkwrzeS0BYMj/4PlQoMDw/KXu3gI8zvlbWFI/f3em9JYludTDb9PDE60nb1zuORp
qW6z9vbaQW4RsUfhH1+zYzBURztQ1IQiSbgzPCqmO1dauOjPPcANPgpNBmQcerTs
rlL3LXl+SKpdnFqgqXYoUhEIln/bLS2Kyt/rq5lzs2LTuyY26VYwqqcPa3NaodW7
SfQdfN9w8vhYkttWOu96hUE2i87JX/9Z2zG9UwKxshG5/rIEovM48eYrJTIC+Rc2
oxVaJ/tyDqw5ezgxhgbMiETYcc8ueWXbaUqS7VnxmRGp94YpDesXB6f+tPgq3n8O
mkBHae2q1HX7Pzq6XmyjsBQ94a65YNUWyQZOl5x/3Fo2DVQ7w59TB47Vi/OZ4wJH
URh7rs50ZzaUR002zIGvPJf70ivX3qMaghxcP+dq9tngHf546bUuOE+TjL1ELijj
wyVKnFSmh2II9C2kK+0YzNpXQ8UG/jQdOE/fUgZgfbRaQzF5AtxVPt7h8YgEQdJX
zTNKhhZqn46ATsd7p2znykXf1MrjIvHX1gasDESj/l8sIRr9ObvM4M0xJgiwcqAc
mb0gScoBaXdaChuavoHmMHDM7rP3+nL4MkKm8iVrqMddXi4CqJ3eBAd2G/6bqgGr
QbMORCgGxtu3w4+TVCZKjMBzsBQ7SxCQggE7hootT+QHZ6oJAg74cuMLNpXvoU/D
SMsoqSXKZcTycbJ+GkwqxS93PXDuHfFBPzjYjV0uHpqZ8Cj5wD/CX3WtwLlsv2nA
02V3WOp4dXWAV8OAsoX0UU9g1ZyamKJRp3UT0rpc6uHszeCyjh2FCJBqrCCDIhX3
bWjELkH+LWgP7LgI1iu++0NP0/l0zg8UrckSMiX6ga+dxjKyGGqbPiLy5PoC8xe7
uCiLkhqyEQtfJjnGyA05dsjEv3WdoxRrAWdMjlh+z3AHh55BmaUFlauwelqEoYvW
UjR5/Qh776T9/3UNnrVLqJK+zj04qIHlI3EOtxsBgnBSF+XwnoeFx1C1FdChtFjf
IM7n3WK18ei+U5ClvzZat7Rg/jxTl5L2zoe4+tmN3fNUxgzQUY7AJR772aW8azDm
yUk2ttdeThTOQ0VVFbhU6BwNenrw3pSjCSdt+g1yqFpfvLeqcFdu2Ze2jFDiLaXY
8bKd1Rv9Ha8cSobnsIIUkyp+i797F/ZU8IET7fbKp0g8gyzMcHcNiaGkB372aV78
Gv4Luo8YPrfhROxOMD0IGWOi+YsjPg1xguPlYg6iG56IVUAtN97DqSBccmYmI5RT
lv7uWpvaPUuEtzxzoHd/rFOaMIwTcFeGIxfLeEc9lTWD9EdVkzpawSl0sUBZTohf
9Z+7ol57CpmVLUpRvEpqK/zc9NivKKTa5nTtbLF4s5fncwle6DbEnMLS5cy4k734
ipJ7HqkKkWv3G+uZ/8lztpZYmkcqbFtiXz3cr0SrlgOYRvp89iwVJmOIBbh2ttwS
8UKeFQby1p4C1xHXAAk/oizjw83EBpFAEPpB5mi6BY4I4HNkBkF6AAA+bBZV4/Tu
5r9c0Ay2NIC0Wypdx/tOb/DoUNDm1d+xSIqOIvRNeTkeKTC6PuamtykPzkt4LkUa
Tp8ZmFwIVz/Y6TDzRm9B2Xy4VYyZ1i/nquaBow2fP7XjvAh3KCYNyFcrMuxc+I5o
HxO2YeYecb0IxtgAWnPllOHVD/X/DbZBPL3ao0PJtYV/pEs6HG9PhINxC02mrrD1
lYYl+rT+gM9nGjPrF1Yh4OOBG9j5jcFpayJKPCdM8iXMLpoRBItTX6rPni8Ug4HQ
TzlWNk2HTLqNlGFQAbhR1pxYkUrPTXV7CVr2ePw/d/xkW4blNPD7o90sDo8Qpccn
fmAtk+jc51QSIDxd6DoCt0D9ebWLgVGEPWdN34+2bJaXYj42OOKAnWlgBfyyTmOW
AKhfncA6+zUfltnl6G7YpLlQywHE4WGld32q7Q2NtILYyFm7NHQQmNWeJt8WBq07
uYJHATVC6oFL10h+AyWgpdTQgSRfrfbwjxu8GrtQuIK9r4HAtBc4nSAhPHyqydBJ
ZABH7OGa3QA7KecUs3qETNrEnRpgr19tQqWstZpi7KW6AdyXm7IWaPeIi46b/fiC
2bmLCmbrPxr8ZmodrCLSMce/SL6n+4XDTn1Q9DPVicYlIBfSG7pzUdikw4swZNOG
mekEI/IZqS1/V7oHegc6f3gQcHBtnd9aTfiTs+Rn9SrXAodNMHifKcBbK6px8tiG
4TirpR48xcRw2Wi8B8nQUL+sxPpWnwH3KRoF+2UE+c7wAYwylb/3NaNEKiuhMFid
UCGXWN/nkwzTxIIXb9MS1xJbHECZX/zCZmkCFo2QgKkb8JC6xmT/LOqjaQ5Xwvm5
jSGzs6OXjo0Z2hI/KFJ+6Q+ZhqB4t3S3aqt/nNaHpaiWxAZS01dsdqHJy77crZtc
Q6J40Ep/L2ksdosWiPGnVyZSVwtsX4jm+HMeJOLma8Od665PalV23CSH0bbmPJvS
0i1+X8Jm0xBKqWk62f/BoUtPAsTSkUaX5zr2MMtu6LvsurTkNAasu3oN8kCbIm9Y
EAqz1DvCcexniK0TObGerDMivDQKL6MUg+4aQBUc4hxrV1U9LcXBYtM1pXoz/TGP
ovngEO8YmhQv8bT9AoJ8kKRVqsgUei3/HvOcQP3KI/PsbiM/Gzh1d0VI7E1hkSWd
lWWCIVndqTCPqx7qnbdMOmMeVFebk2LGFdwvdn5Rb8HTpJ00/sOQIm0eXFesgwVW
d2mX6reVP/x07KzOVWTtg7JOBBrKHqxMo9xGA9xDdHdhZVtV1+RsvF/NtsPQRYTh
DbZ93LlZL9yaGXTj9IkqyYjj0CJ2zhrO+zWExIcDsec9xy1qMtb9Bneo+r37Mp2a
m8AxNJmr3882mq1/EUkfXUQG+vybqOmSAHIIqbKeDKud36b5wnV833aR4EVya4pV
+zz52LkznuP9GsRm67Zq2zrIAp7jt/CZhbPYfQHtfDc8AouNAM5VjB8jlDRBteRD
H8dhwoy3dWaDdp5HMKsRjzBZc5emHNMBqxpExGI7KG4JebGMibAJnIuNYkjO5gEu
4NHuVZoY8NRy5Co6UACoun9xV775c1O8uw3HZurd3uGHvSCTs1iuUeeCfikJqnr/
A33gHBhxM9donjqYDEpgnSWQyo3wE0vhK/B7GXLAwVLHf2qEjeTMdFVgU/5NQEi5
WYZ3Ex0IDi8y1w6m8nP0tZSHYPziPT2I2XwIqNQjAX6A2aM+20L9/u8hOI/B9p0H
mYP/RDCbTwTrHXqtlx7JRvkrOd3YeopyuevXYNut/TvMdjZrcTNN507pDImVaCsl
TFj+a/Je8TCeMg8m86JKwtHGveNzq8Vq56tYR0HygfyCM1S/Lgv7OyQnkEs+BUkI
qIE1taD9Q7E0xgogvljMCEvk8VXO0Fbr4fevnjrmJjiGmDIXIkjcZlWrKT83HnG8
sHtAIQ0mOiKeZC9G35tadv9Ms+ChSVqGwOQDOu0uZ7PxLdzCd2Mp8/x0HlgSzCR+
w8WlpHxfw0CGwVXKiodGVpy3HqvvoAKDN/3BioZR0xf4S92G0U+m6KTazR1CLvqP
lSsPey/FHx0enkuqRQ0tDDOfQdZueJCjNrEn3HXKCcthKH4zvOFTdujsN593ogwh
gweH7rp84OhduJ8G5PDMn+GPtPigWt1FnRp5gjCKB0Mccwb/et/XHa1OsU8D6KVC
RAFrHPRec/Nqy3jQwzzin2UhrD74D9qpQlJlFiH0I5bQbiZW+iA/IKhqjwZcn9lQ
oywrzOWmmDPVKfyPjZlvtuR5IYdwjsnxWLzyZykqGx1hadbjgw8plnT75jEI60ZL
bwXEInuxA9f/fSGVaRM4lm2C1hzrbFPlT5yT1+LpxX55jGHhJbAtg8Gg14qDb7ix
R/ZzjpMZUzTyEytXcAHLcUwI0xLVi2PJbqmKTyOHtijlQSWRiu5Oorzimb5etf3g
YEtqDEx2KXgtCCb95Mbd4OH6soWpoYJMf4KGPvNfK+bYNegHBQhC7bZhWm8eujlC
AuQsnlwASFcFiGAlw5CHeKC+k3MGU3iyXzreU5jNsTlXPeH0+//PI6hPr6bFJEmI
Y/1q8HxDc40Hz2oJOKlfFZUuLKGVnFJXYdnzJmYJIEr9YfExifYRurJpoGzPE5YV
14+xKRe9ljzhuNzoBM37Mgjmgne4Ggz4nj9wESvPs67u7wt+MuOR1RRHJxtGCa2u
jOSoSPonUpMbyj7U8wtYGW24Z5n0GSQrOHXuAC50yasZtZQf7Rpga65qq5D5Oo9z
n3DyZp0FNE0LdKXBki0K1u9eV6V42HJNbIDMRiunO/BAJQuR9L4o5dF5BuLgfMLZ
bjaBikpSpabCWlKXJpziiQPDYD0QYG4cXzCKPDmZoZniMzOim6f1tGwyeqKJsnQd
TE5rC9ZPYqkDw9bYMxu4wywMZg6FhlEN7tUmMlFRQERW4QZee2xgwGobp8cjZ1Ev
EbgWcku6jrxwLQVVLxC9BOOxksNO2NElkQon+8n0OjsYRutg7AMPCZPUUl5ZjS46
O5bOPfcHuzFL8RN9AKhUAWVmAytj573+CelBKN9TBvXkD9zILVWMSmci3QtmFOU4
kn9ps483Ue7yLbBYeei0rzejYSrmgb/FK4At1LRnEf4lzrf4iVift+Xj/cgUmEak
1Kv/sMl4F+6B0SdZj7+pC1algDyoa+9C2pOQVmHgZwopDPrWcmPcou8mjWzX0iC0
06M42ArlAyA/J3eb9dXKzwiBpe1fE1Tc1eJmNoHwPWxyUELQwp2wF8vKCrss2cZP
jcBwiV/sm+wWCU6KcB/IwKxA+lPy9ZE6P47GMaaCcmtjqRQjcoHPY3sJUJ6cAm8u
z9aj3nORfkyGSVU4YIst1o5os/6+0gR835STwCN490hSeRFMqdwXVckGsvmkc3Je
Rvczpx0LeEuFTMWbsGVNubRXt1Hf5yODbg9R7sXZ4Z76kjN994keEJ482U94WPVG
igsBmye1mAO1YAcfrGA6bwpl4KcpFbF3rBn8JQinaxfAX/IcAS+5Vvnpc7YE8bzK
v/G/etLsPWlHrXTq3npmLi9CjUkYHlHQr1IjbHLXrE6OANE1knZV2xOcCJ5oxUEw
x+8SQjsxexlFD74TuuwrwPqFH+SNZkXTytIFFncZlCrTta29HCQplWeMDP0PA8x7
vJ/Am6YEIb5Zq/W9ALKi07XJqpdOEnaGhnb174PyzytwV8B5mke8PUKARdw+kIAF
ryUBdTlWAAm5OfpG/VIqBPxn38CMUG9CGSOo6xHjHPgpPtok1o22wjdH2PhyDKBf
dG8A9dVpRw8aHEH7JRpURQnV4O1IObmnvx9zRLsVtNvgRzIt+KJwc8lRxhBFC/aA
k5zBuC9JDE9mi4MVu+Af4pWp3ADDDzkwQS7lp2FOTc7Tr0NBmUq9jUzPZjPLGzat
NrOWLPpofQUvADjljjhROJ6JrtO2hZ5Y83QaR1ApKniBfobChfoNsWehkVGs+EGj
QZ9Ekn4XX+HbJlrpJ/a73/gJzwdhVQ5f6qjaJYpuJMi1ha8CteBDwt4rYOqr/2kO
aufHWq0cMRs4OFiTNOIhg9an8ONf7DjRVy5Qfnu5HSyzY8d0MLgBnEsU5bQtzfS3
WxX3mMMJFEXiggeXrZ0Sx3oGdsC0zLOL7xRLA+NJfB1Vi+DFQadShx3PIH2aECnu
jrrVYQU9qrf1panXqI+OFKr4aVcaZ5DPKtadBhUldParXVWeQb7jE27ExCDpqwws
KxCUcBhQ+T8LULOfJWmBygcJu346Uqp22U7B6bPd7evmav+ZV0b6dj0np0B2EKu8
bEf7dv2D5ouD7A2tU7uNw29JZ1mAZHNYgyrz3n7yDs5o1Tblwe44UNU9tdJcDRKq
sSyikYGuiq0Q85oPH95tUu3UXQBl3tYu5r9Lv+sg03VOEzxyWQT1UZEdopFezk/W
SOgHCAriYL/aWHTNGA8lzkqdp15GMTCPgS1asddVA2lTObfiqvSC9hmlLieiKZTt
TTDSQRL+/H/fn3EjpsKoZsSJFGWzSEDWpgeNYvt0aqJJvy5o1gHHDAECmfyEKVih
kqezE3GFdeRCiIZH/pyvC8DAB2M8Y8Dl2meUkerLiXvuumJmKdaa/56HzvEVrEnf
SS7nhqxvAJHwYyy9wfxB8Tv5+cnyhrNAibUehcTEztHWv4zCyITLJN88ncEjwmLl
Dt9DoWiKa6seH2rg6y6QJEaVEU+9kZqdVK7lqi/UGo+FClV9ZEKUHWlISP5ioiKR
sNojNpjI5vbW5zTARTviI63bUSOSOQr53vion8J19npgJ/LaPjG6wwvLp0qnZXLt
Qk6RYux5QGW7D+HOnPrMjSH5Gqwu4XZNMz5vHMhVofcwU1DIOuku/cX9XuuYxF31
5mM1NUATJREWT0fDrfdzVnwIVhMPPJ3Y/Smf1UzTzREr4YhhamMAvuHuBxEP9Jb8
wfmb0tq21InfDbbvHlfVNFazvdJ7DWt29dECON6TSmout5bx0leTGeJK1+Tk2ZEW
TLBKMthmuz6BaDKHit6KZD/Kxm/k5hkcTqD4ffuYGJ8uuxP0yJWTDOsSbAVXjfX+
yXnGE9kAu54lnIbZVHc6Oz+9muk8hiCz3kJG4dZDVaJ52NI7x0b6h6imyu48/NHJ
W9vfxlTDFDRfvnr9zCbDnscEqCMOWuvei5DnTKI3LADKIxkGyMpbpALaycN/FnMJ
Nnpp9gefVPlhcevBiK81cV0hmiTXbUlgtYNx7w9aGkNEM2EbLicC9Pq4uCTpQ8ih
mXvHxKnbtZxdvSDPHiuOUi3zxJhirhpBHIlVkksZ1VvjvbUyPL6KkbwG1NdEBDfG
isopRdSucrGnpoUBWKwzcAA8eSY6Ceq24aII59OFYlRnO9vBIOxzTEB5LQsdCruY
/RXir7ubZEGE5L8i4wc2ovxXhLgHDa+KtYxvLvhDeDgZl+HZr25LFQ/mXMEY2ul8
vwxU4nH6qpqek1ZRKqxbZcymdHActoef1As8sw9CHLpTwpmNCcZgMfwTAuiWu/Dy
r8guAfq3suBT9yO+rZdbgBCykhXFSkowzMARUlUgibvp62dZCXXYScex/76+3gV8
z18PmSblYmKi9Cc0nrrwkkvmElZEJ0SecM8gN3XREggHV2H24E7RtSj56gXwSpZ8
IpGSPuJ0aqBHl0CTLYH0xNJEK3Wa9x9Q3omRUZ+rr9hhvZmBh2BArt2MQ9HhjurE
9UD7wk6sYD1gHztplLHZkbi1jZpAVIdjydYanHfxBsEuQzn7iQfu2z3poT4FEh+W
wOiE4M8X0nil43hlPnMV1xSgHwja9nNTYV1Qx7ONApPGbtggMOcMdIpc/NMj3SVg
57PnpeLBpZ6WvXYGWLV6ECwneP+wEsfOsjoWELHj1I9CMQ0DKWuYsodU1Wbs1KFT
M4pvwLNQ3RQF08+NBjVimTeCSlDkGCZ5My1x870XQwA=
`protect end_protected