`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTF5eD4vnEDgRfA8fED2ppvPpWrRC7EzAw5tmm03bCsJk
pTsfJgVTJbGLnaoD3Bjb4hMJ/prSwpAyenEFsJ7hcB7vkE1jMkaE7A0fFgauCane
au8hUHiNZ3lV3s8Ia4ihxN16RjHR8H15/jtTugXorVYMWSJrfNkZQhDmp/ttMd3J
yKT0sWDbPok1ehAMzV6XvgalYpdI2XwCmT8tHlXZITaqqP/X0KfjCCVZa1Pit61O
cKkTYDFab+xySrmbEStamj+Jl6AVZPP4MpqZxPEFTTTDAtbxhxPRAolRjnbZZvHS
WGodJ7+gU87H0DUUf+HT6MwpREMunapJ4WslmkKjEuqGUhfL0YCPE8BvZgL6LBYl
kfBTsOgavauZBMPxL5oPMCD3KOeLn+83QaHd4ZdplaUY06lRUpo+QPJAMBT7t5Pb
BgYDfnTxSQ6K9vQYYRxCh9WRrjfc3eKGK4KZwIqkGGSgNLdMt30D8sEYdYudbngc
N/WNV9YTpj5ldPHbodh7zrBcCwxd0O+XtvUYDWrfGdLgtPddovGwHKr1cgzad9a6
GmJ7NHKPSW/7IE5SEmDDdVY43c9TAQNpao9DtEiQ/pZKnWnvQSMVr/7L15b0La5y
/sgzmcPMvR7GZsk8MTzUHk75uZijw4S6l7Wc8ps/TxcKpaNCctd97N9fLzqk6DmC
pUG/UPh2chZvugn3FeyLf9OO64QAFcRMAJDeFK1G3QmN9Lcax4a0n4i9WZwBaZUp
x+6ehUBGt0WDOCmWFkTLUTVJQlIYTIyA6/n72KtCMJzE7rQVdE78wktip5FdsxtE
G0B62ob5vJUmfx9RKr+Zd/y7tnw3S8mJCOO3IOl2dwCFN09fVG80TIGErUtj0R9R
Bb8jzZFXcNv4ceu4P2D7aLGeBdDOsMG12WU7jB6TiI0qMzR33ayxVS6UdUq8kHIx
FKcDZrJGBP2YJ4GV2Xw24j+XwpCPFcQgxFRDpfQ9Qbfn75EKvdjEb//Ydde5AIw1
uIKkBWOM/f2548Wr3ZOOw/C+YQyz7FJY75X9o4lsRwDJDTNDxv/SlxJE1YSX8fic
LXFK4yAiqar+WGLNRQpu7UmZd8MeBwzu9OH7iZciA8mhbQvEo+dmSQsmRCzfr8n/
h/u7YU0JiZZWMNU8WdOFq1H634yf1c+IB/ndqDpEOuemMAlXxCmr0S0ubOO+5Vt0
/B1sFdq94MrbMF7jwVSYuJh/I5Ep9G+SIiKyJ5hXN43ltEk3+VoHlhh+meZRut/Z
UkM5X9aw6nbhmjIV0GWvcZ5REspfm4e2+H2cEeuSXvb2E6qw/e2bu9N1bIO5ITt+
xo4M4GOpwCr4e2gUki4z+yWG6JTt3oizGUHFPJ6KBiyMTaHD0Ag0Ngx1Hpkbq3HQ
DBFAJuR7MZ15px1Ktf3G/vjMNfw0Y95en4/9VfCUpEnJcBi/8TrKR+Galun+NTNf
5V2LN+cZ8yOoNCOfwLzsqS6bau2lMTUha5mcFsaCmNQQu6Na4LIOVepG/iHlMfGn
jpfZPmxJGyn2/AK3CIQhnHgQU8m5vg5Moas9nIPWtO/ttBP086HetOPq75xDFUg8
FoXVJXsQM8Yvr9epa4MKIcwCsxH8txOxJ1cKdkVr1EH7vOjVEzlrzIpZMNx7v+oZ
hgXmWZatOoHyLGecIOPIti3KLT2sMpjxzfoTDCdJ0pYgAxdMZylKsxxrU0203TYt
OxcWK7REfB9rkv9YxWQlpHR26g+U93mNbfJ6ffyHtwPy7irs7JbFjPEFhJ21bxJb
Q6XOi7RQFKpL2HsN67VKGk2IP4vy2E579Fc06EFU38/noyecMrLegPsN9fE74IXm
HYFKjYi5erMUkxSyhigBXwnlWXjVEYI4nCPywk1Ul/hc2b9LrticVbY1Y4DyUo3u
YZzt7P1jJ6HRe+3o2DMONGHpDwWHto5jwoy601izGUEt0+8xryMMg8pAPFpgCIBf
G2wk9+8ERIh9qAD0NEoJbgCTq0Bhctqwk1bHjfsT2HbFg2+SDM313kwaLAP3VDFc
xq15nPXuOGE5WSmTWhGHHoKFhlZq+sgm85jmp0n/b7Jgtn2FStkXO3yw/QrssvY8
TdP6HYyd0bRAZZ7Kc3TuYsCxl+VBYRNGljmXGvKjDgjPW+j/Gzjq1hsxlwAGt1C+
18HC+sNQ5QhfnmEBrQHsfzeFi0gcz2FS1EuDuSO2c9ILPiuZ1WHeRrAJHmeTrJkF
i4kcx1XD619sLG+akfP9RBPgjr+Wc9jHBO4l0RJ9valxrmbuvrusnxkd7ZB7ClrN
7JjhqYysrSvJW6VroWAO8yzEIuhLTC7M8xw2o9R7ff78dOrgsg1X35k7y1K/EEX3
KBTktxYwU6KVUBypVlcae+79D+PWoRPm3z8SHvaMnm9OzXvSvOr3+/Zs8Gb53H7L
f3+Cm3RbgUA3m+6Ldh2tTJk9nFn/TWKyHioKX3R2EGDewDznn3Lhg0UD1YoPveuC
JFu+J7Cbfc7AYUrjbllIXw0o5FtoYxiMF+xbw9mo/Sme0FuzrqsX5XYOTjNA5lyU
OfITu4CaP3gARI7lmM8sjuK6JLYXAd48hQqXwWmwGzky5RcMRFqmCNFcHWQ4r0kF
5waGmx2nvFM8c7hAmlWJwA675wcGb/JzZ9KeAYfbbBfV3mL6EjxK/lEGpIEpVGp+
ZOksMKELvO9VQS635HexQdhiD+Uq9v4LMiVqzgL+qhZItaGyD2fIIgwMOSDBEOc5
fK2an7c8uwhTiwzxc4w+KLlewZaZrrVqP+oIH7tOh6SvhXwMGBhcpLDNfwk9/9yL
Eubps0/xcGQq06uHkS1v7L7o77NT1dOilx8NmAxTSpJNq0Ai2897Hcs8FV2VZeS6
8IDNbvbxGQrH9Nlv+1OQeTBBQonYi/s9l/TEsNU6kdYx45bt3jKDh9clDk2E3P+K
hd5zEYaGVtjR28BAjdmWasyH1egJZLEDx+zP1R9piMooxgCmAqLi0DMcYeTalmr+
g5VIvm64Q4+bFbIFEDioiVLz4YWHxK3txloPV+KAq1PyZwzxwknMsNlJQz2KffSb
89XGj6kRZDhSI3DPl6X5y7Cly5HHc2cHu1XlCzH+QeZcHOILdkocqxhZFbVuz973
dyU+T032SdNnSjEaCuZzGM8GuMhqlJ4RFflrxGvZ4P+Fuwgni8fHRKHrNrA6lh/+
cNTMBISCuQZLPgfiQWso3w04V9dVstLXszm1y/6dVjm2SlyhqRz/mPNwJGz6S8rX
Y2er9w3xqc/uKoQ2tbqChoStThFN1wyUpRr/xe7a++ve3pN/1X52K1q+zJ50oUZf
/VqrBSI6w4ypVi8+OTFSlN5mCGTzRTQw9+AkFGxaiKnUVYjA5JhI7f8z2e57NKFX
WfK+gBVeFy+j1ay6z+o0ihqg9DFFXVKs0gjrkkB1OqRe7TLFyuPA244XdJXJecsI
nBhnjKG3tvZcON/hPmvzR7CVir0QoWg53QvLPuYVFhSjBFu0C7g7G257/NF+ilTQ
YHzZyBzLRMlEO4yip4cTXF5di9HE7k2HJLF210vsfVaSYdNzNbdWXpcoRzWMR5Yb
ZiGeBsIfaPXAO66oIr00KLnvZVJ5mF5+WeQYZh5hFZSpbzviEc+UQEtn5FU8zhdy
p3U1ioeI9pJzQLuZ5+CCnSn+qtJcH8bVGeBaDiA5q5VLKyyYbdrP88a4lIwAT57A
Q8P0JmRm9ZM7XD7WJgt3QcozjAJqxWikfcYoZJG3ikjkGA7QyN3i5aDgh8Hw9uGg
9ukrcsbv4Bfw2qtMOFDxlFlo6WJhq8B8qMSTHxL8Z36wkzLhEIxBut6JpOvA735g
hAr013QvdxgXQmR4bjmE2ug6LvVnSwKrGATEvkm5bo3MuLNGSvg2NDHungm95TNA
VIyMrPCOEcGABks/2OZzyRzJL4cdhlEJ8SAaHtXEdEiZmvi6i3olno+Yct2wpP94
ioQS/ITi67yD4QCTs6COIxJXO8Ojzj0qtkzL7ru0qx/GSZxxOOlieyXHzhNwGZ/q
/ruEBbGd9Qe9sH80TqZciicMLrpwGAn34gPowvnjeWpu4I08qAKve3/usGw/c1EN
tP0vdUEh/sv18Jp3ALpvZ5glx0gCW78gx3ayGeQBuCw1GwEkjEADUzdyB6OTuxv8
2Enx27slzbJWRiPvLBozdQRm25MkO5zbqXssgVfZQW38+SG2N964hu6ncST3rgn0
wMtezPc7gANIkgYiS/7aFTfrrLDIYXcBes6c5+7fzXkZISGF3291Zo/2jlMcrtqg
u3Idh0v6SiY6wjUlawFErkFx4TeeRGKpWZ/vMSVuESrX8WPq1CvULeMwnJzzV3BE
i9vsHBpGHWTWac8X1WvyiKxdkut7IMVDbG34Qu2p1dnM7lcgbq4tsFipu6EW0jLJ
c7UE5luF2MjIunhO8iddoycgKkkvDOn+wzCEaDCiqLmPGGnXW68Ez03bpedjW8rE
pjO5aO1bck4LRiEJItI7Jzuk7OVInv5upueeRFL04ul+81p4e6DAAsBdQbQuwCNY
6uasEEv8Ir9u0v38sXojGRP5LzJ3n7rygjpfjt+j2Z7s+A5ouaANXBwD2I/OiMFY
v1zjfQUdKm7GpN54ds3h0C/lLZ91pTanRgXXQT3/s0iY3nv4HCabqWiTfewjpUjn
TjJ9M2GbOxdeD9bLA/f9bpSIoHSUKC26odBMhVZY2jha6bZkQijjuVyMXUNLSONe
MiR3ksdJ2eHPKz8zP+Hvu3NKs5Ci0xt5leIcH34HLxQW9djDEARKl6tuXbtBS0kJ
178kFPv57a/7ogJGk+SPVQ216FY/6CFTML6TroPY3ibSKsExFXBFh3U9EAHOp7Fi
nlnLajHKpVEQ/nOq/q0q5Y9FxCJ2cMeLpUJwMxViQjJIl3olXWjaLvUfnUjd8EUK
/6yKcjyqiCjxccHGkDCHXDsOVj+LvwoFTLai31j+eoVqSJ9Cj4m04XV4Y8Z4mt5d
4aDRFuXtvjLj5OfUs0aDFhsZJ3jSiRFifKaNbdKHBD8pf1KxLkhyBuxraIgKy02O
/LqaSrTEikT7sM4FkpKpjVqjKiDqHnjI9OwSCuASApIQpFoxJOcx0lccCaVAO99j
/kiicY7D3YHaUwnrfYEIKa5y8W8ZhxYMgKEiAXV2QJ6C8K07nGWj0POG51sckDsA
tAYJWK/tLdf8nPDoi0PCkPMZRnaZG1V5/Amzu5pP5u6uEK3mBK6BUqNhuBNEABjx
VHcibsH6J/LMMCOOJvcs3S8NgCv935N5+DtkM2Iwg6fiIwubpXIjgRSPWVabyh8s
6uevT2jqiEEpdqfXpmPb4cdIPiqo3IBZIpxQi/Sp6xFxnGOZkRqpSLBExMp7skBL
SGeFHrn51iJiZS9Cmu+ELJi1dPqrzKYfu3dfs2jl/r+bkhUjS0trEvuKunoX9E+K
Wxv8Z7kYSr14UkAnf9DVrpmZ6/XC1rlz9sqtyuhCcdwxUvn8vZgG35nCXESnuFox
OMIG4ffNS5U0NlunWmbxX8idAy35RQ4cXrsFCxemfYpLoYJV6isRFRsYBdi8VthY
+/TuP1UFh6ZLIt6pXl1HoQyfatCJteMuk456NsMSg4GoBSXRAH7EM02s88513Sh0
Jro0v2nUOAG8H2/g0xU9pJZlrjO81RBcSiRwh9nPCv5mlqDgdlv5e85MAhXkfggL
e4uV6qxQ04HAX00CMHuOUubjupQEhuQJKbDmxyRinftkYtu7Q3bdJDY7OgZNfOb7
qp1BEAs7NV/mtTzpFCSpFhdgBPEInK08kooqWssycMi2/9LGHPjgG7tbUE3MM8cN
7Dhmr0YB66W2btPsE/8uz2aZfHBAit9CGTa341yAmXnO1OevbGq6e/gvO+K643Kr
IaeoQ5VaaL09nzgHmH1H/D9L8onK0z6omDBAaq8MWm/03a5BbQhxcOFIUz7JdvWq
LubdrFSg6Gf7pFom0VyFvHZp33wkSvdbmemfwu/yrBC8OgmzacT4hKMAUfnsw2O0
cNP+a3+pQzzGS+ZDUf53+YezAdBFsA+AZ81U7XqKUSI0E0R8daOZ4Ucynilswrdp
m0Tco8mlt/1S3Adh1hnVnBejCL7/quTqzkE5H2WGsryOIOuaG2/bW98Ga9YoABLx
6Ttl0gwaUwPBz6O41l3rzXFdeITs+/rh395lD7q5rzan2clCNZrFlp8JOpWZhZ1T
+rTdGHE+jctxGo8EGJ8ZaXsxj62bXrFh9QJ8PcN0GklN8WX0usVzbByT8qTpInS8
TwlxSxzv/DYNRuCuHWVJiOswHdaYULhWAe2pNNrwoxo2rAZS/QxVE5SS6PPz1Xm4
u9YFOPvoVVhLjtvWL230YRjusLJr0vopkMPKGmvoPIrbIZZOPyzkoxwucQFgquhl
8n8ArTDIFbfjw/ozkJ9v8+EPWfeVlXDoziaeFV95xJXaeVLD4jMcF4p3BEHY+5wA
6Onc6WzGuk74eGB0cJha8hc3C+JCwoX5NNGcpRD0T+vo/6NI0uIcDzHk/nMUkXaU
iikUNvQYwJHrUnt+I5ni+GKTV4pOY9wskZRziMIqKTPGy4oyHeyrZts8vzBqs8lV
NrX3oUFNbVTecNg1AOri0svdwGVShOlOPx8IRyE+eiWod/neC3C60QZiO0zmOG9H
qg5AzyltvRaiLVFigCr/86MbJyBulxYh9+lOXiGftbPYiQxcrkjLfzVwP8eyD0vK
IuRz9OjfASyZpmUoXWYx9DzwKx6YH8bzeaUlJ8GFmfMbkAgEDXnDfPolAP5qkcm/
yLM8EDf+OxZ6p+nySVeT0VTrLyFgfGNAjSDaLLFyKzLTRhEs4T7A44Z8HbGoQl2O
/ES50aRCag0rnflMv/JXSAj06IDw7AKNYZnIhDNlNdbbL36gWeAEj2NM1beYnRFr
4tIAXzcg1wDUryFkuDq+gPqpY5aourqQIiy+SVYt/umE0NWghJOaMee9QQuqJWPO
PkuOoTVpb7Xs41IR0LiCmOgYm8pkUt7gHKsf9G+bZTOVjbKo4fZNpXUdi1EFfOtF
7GJvNFRQJGv7F0oBnCKNxHSFPAKRk6qdbpYF1kINgK4pWHmliXbvuYZFg92RmwuU
YLyqB6Z6n/75mkmst54OtjGCOXXd0QK4QEJYOE8vyiuCTtZsA+E4DMPqG4tYhzaQ
p/XVo4/EqAzI6qo5D2T5tERSa8mekXjCf+g/JOUioEleRLLyvnbnDsJdRTxaSpMq
Sq7ccyxNzvE4YzoWOTzvuoo+m1XRXxf7fAQZYAtgBXfE3xKL0xEbMS8g1OSGfkMh
5b49EtU5qQY8XBJUJvQ6+LmipvUN7vc/iFb6lqoet4ImNDlJ/MJ+1w8T391cH49r
xDC0GlGBTO8X6jegD/TNIKtD8cy1935PRBfldtz2959D2h+OT6+73R2ltvzfzlYd
b5sn1MrB+hTTBziRSNMbpbLbKGlAwz8j41IEyh5v5XsoXZ2TcHmvL66YU6reBvaY
FDBQFm4tDzgv6Njmtbg51mzr1m5origmqseuaNRVMXbJGqnXAYtcUn8/p7o7xB/2
SSpc2urGih1X85BE5UeqWy5ENH62llPQ9RaUc5GXUMvClfQG9IYrvlWvWlL0VMHO
VclgzmKq+Tt9zvouaCdf1lDz2NctuWclMCWLYe5TnaMIDQFE1ml/OqbrNEGCdSfm
zlU5f3fuRxjP4WeRYilPnG7/1cwIDFpbqveOFsfxjoPb4vcRbozmY+p/EZ1G+WYt
4R7Jnd9aYJVr09d9uv/oaaqZVi1B+mhal+ZcPRMU+XMTeG3WowQSkhMNw7Ynl1Jf
V7fQw9FBD12l/D6EpzYdNfXw0yveLqfRyeox7kyIXlN0tBr/JpqpSwrqB4OM848j
ZNpG0YQyHGKhBOxg/QDTxS0KW/gl6uXNQYy1qSFWzCLSiPMBGV230TEWcgkUt2E3
J7PPpj8QpfMvEBAON+WHk0kfIrnR1oRYG5zuH0GIX2V6vVJT1/4+uNOD3O5FqlIq
06hFNbO1a+3Todh0urVR4yfFujOCcBBCnF3NcWmbwMPnVstVfY+T2FNEk1U3/7qk
UzBm6y6nTpfPy5yYq8WGV3h+GjiSjBbb50ULjLUcE/zUBn0BrTfkeSuJvQT3N7/m
P6zrcxybaXAvaXoqfDxQQ5C/i6WyhrLu8RVS/hjpNnP0Z5ZSwnWNkx64z0jF1ICD
B150CWbbg63N+zqSZc10WRLCOMruUlidUivRIFj63hO6OGbUHGJWKVsNY8EBGq6I
4mmKkBD0mf98QoyZgF1LiigYpC6afqf269Nz2jQJEzA3aFXJAlmOrn2Tl/hj2Ajo
TszwWgEn+sWvuAm73uVKyGPHGIlAMg5OuV9PdaevmzSwDIP4aaWUsVDQ3ooMNNzS
nW6t31m2Jma0JxeGH6IHgrI1uROFKmRNGiJ36g3CaK+frzKRmUr5+Q4tF95Og89a
PYAdz3x40TSg16zwsqsTEG85PnmgakX1+5ToqVvJkgGNBiktxs06XFSfZEivu/Bp
HU+nbEXK6lCBwNeWyt8gKQ==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8pZkAFSqnBsdB4bulsx5j/MQKipSj/mjIP7wpaCLUahx
hoAzS5pTj5xU2d8dpqmwZKEioZTx+NnxoWulw2lG2Sde2ANRpalERd+ab7NoBhXX
F7NVBtFxVRZsekhBB7cavZ2MJWFP6L0mUjVZloiKU75M8VsovYsFz89H18Wc+oOy
EfuYW0BC1g0QQch0BZwn7cnKoEc/HucBc2fbHRPIxJErh1L4LLrXvNtdUX8bddkY
/LuNiNRytXhnIzDKrlQsELjPy4zf00IWmHhh6x5pjteIaTPvn+5IEyq87JoVE3+E
D3RhAl6KrtNtIg7Vme/7Z0+BAGScvsfSag4qgGOpW3wjJcxC93Rlgdwau9HYtTQm
tsCVMDnPJCrT6eWRb9vaBMf1gY1mBTHb7sUaw2akGPUpv0d90ruBmIrx78IkgpJT
w/p691v5KrPVg2JNG9AP8+KXISfyND9cPbjjLk+KuzIGsPfV4JHRQME9HBUzp4nA
1jIJg3+XBWm1MMcE9lo4E4zrxyWNVXu3fY1DInwnpAYzp567puTVloYcxyvSxN8x
vYKn7X8eAMAlE1RNkikfsbQ3Xc8AdP8cnplHfJ319C+bkZpZktP7oK3r97W9o4Ie
mF+SfDhJGkG1i7LgXuoR/2Dim6dE+rA4E5zvGav2Q24yefC3JM7TWMyfVIJJd8mq
ndCsLVatBvdxz7ezy40tTEtxoyyivCD8QFp3fsZwgIp7JZqUl9M3NPgZFbSRcERu
hYvPud0jFikhXBhlrUHdnnXmPBLgNyiWLH1SjAQe7U1GD0/wES4wfG00/L5p+45b
4PDrrsZeNgS4B4vyZGQjNewskFQvDSesJUVQ8LHoGvzXY1hU9cGTpWiDaYTVDiyB
saoAMeMDAeKGpvuSKvOesSsrAZKLyVr3McIhskqtgggt9iuue862H6Fxomq6p8Ro
84u/u9JRHvN1pXLMx6ows8U9iwuD/eSChlP5viB3daNq2tsm4+xbVim4WhfTR+Km
Ze3sSr/y7N3nwcM7uqZ2jfuVaWrEJT7Kh/iXPo3AAXx+h2TYvjzLv1jV6sgHItp1
YWg56uXOQMhSs29XNH4ir+SmcjMnP9we6BtZSU4dVucB4qBUmPUIKQL8CEJsb+0y
/X8g+AX0EDqEoTZB3mzBCIUb5vsBhHlk9XXtKMzWwJZnjDeaT7C8Pt5KbLWmP21F
iBIT0roatjzyrPeJXrk7Ah2vDQNPNDFagga/ZcvWnAr12qJ+QULoVVziJPqrqKBn
m1oJFqPqRlqXJ5LbtiHbRzJt4IW3566DNkTBDt/gxyHfpkKBSExw8HcrjlEdFG+H
L9Txcczi/iVguOxAigkyjQ0u14ZPjEMLV0yN/VBtXvj/oCo6OwzKdDvNEOWuD6+Z
RD9y8n2VxnosNhzB9FNFMxqi9kNtjTEr8XFdL8AsgWGOiG6auCLTpPWg7xJfu43B
J5ehAtmmFp0cNyZaMso8YfftHQzjE+iLJtl+dKqTsPX68QsItDb1QANnCzAyccJj
vr9vmiRs36QqA2gdqy+vbKsETbkotvnBxY3H9HvDPwopdxSYATDDzfBNPmiS2yIU
/CtxBtUhH2Fwn72R6W18ANAdP/qv2w2Pa/CKF7KBtjHBGV0jMPqz52xw6EZJpdcG
2AlW+8sPaW0I5FH8xfKWmRZI7BDndGen0z4LwYJ5DO/18LxfkTK3BieH9/0onB45
DjSwuc0j1wn7y9xGM4fVBDOkigsJpFIWvTlJchOujBqq39g9n6Lh2mz/rzBjuq1P
DgUD+PqjLdaTStfjKrfGfoowQSA73bnuZ04ddRWwqsOJgy+XkjSBBoXtdSsdYdey
2lCMuh1ADyF3TB+m9SCaYHLIeeHRxWtJLxybWKYvlUu5VXC5hk+sDVySqeQeNGWm
LUQwzSnxvw1THsx/G8WCGfkJnYkyEwN+INr8R1PpJKvRugvCLyGjUpXfgf0r6Kih
IASHM+vxv6ANh4Ih/RHT3aStk/YVA2Kz1JUGS6512eMoVUSedGSsyhPEHFAxmtb0
wGMWCdPeHxhrAcUch4wJpyH/6Fd+xXD4/F4VSoKbDF/9uJGNzF8rG+W+c0sgTuhc
nv7pIl5lTug6oIVgNNxkIsqiLEu0vHX7ye66MenLd1796nWo5I6EtYeW04e2l+xb
Rorstc+HlQwbbD5ZEwNOwZzdowgeGRGRBu3n2qSOXG81oFHk16C4rEZ/kKLXWmG3
J+qE+FUYk7YfbNFHsxcHYuPaKGEBORm2PSI2VzSDJRefC3YavR27ZjXX4KPlr2oU
tc+2q7XcLgh/e1Ai8ULj3KGZFJxz76ECWIF7lC5cU+K1H5HDfMhuvBvncvhGOyz8
BUEkZ2GYkbAfpa2rbsWPh+SewGXSQyMROljLrF43ORHUTFmCXynigCu2IftNqBd+
wiPYi11D+j9nYTVyOcDs4t4qITOG4HKjqEXs4j6fBrl4ggFP5khZitQ+J1P49gEK
fiStsdpLq2pXaD/Rckt8lFYhLuxE4kDbLNR6sYbPdpn0jfPfGEWnbyoiG114C7NB
oKDyTj4YmAFghwXZXoP8lzHDHRcxgcE9jrkYRj38Uthf1FHf13loXjy14i9v0hJL
SvyWPmU5YjaBzBhOKNgFGczYeVxvuP3qZUn4RVU1dyVBZiWTK6vlUUNGTCFdnLm4
mxp87jVlRR+OB+P0rMZHCxd1ujLnb09svHWNd3nrWUbsDX6o9VBK62g/Cs/9iZFr
i6/uik6nxX9a4zRQqZJ7ctjn2Vy8HrstbA/5bcKPwL2G7Ccr5XyQAEwEOQkce1JS
Jtnqf7ud8XEdK8/LZv9mkF+7FDN2uJl8Y+cv2O1KsatjgTDIyf96TZrufv1RLkBp
zeBDelKoFqDA3ei6ca3vG/B1J8qLjNedWcFZ5tJd9nNBJo2pymAKfs5GBPEXphtc
yuWdVoTwFBKW01lWL7yrR9B20VBE/lckrz9sj7ThoaB1u4GXdLUAc0c0+YlV0XYa
tg3opdWW4c4szBQ5fhnNH7WcyII0q7YwbvTnxjCyrsCPUWIaesFyBVlryxtarPWk
BebSvY9+R/DqFxgex6piRRtLokJu8GFjGqqJ7yqhTHIqxUAIeyCichI41BGtAVUI
JjHtVAZAUuXGX8Tkici9Gg3V06xSSVXOUlk/1BTC/exXNh2ukRY7UNHiea3mqXqS
2oxz/WMuZJhDemenVoIDDSPrNvLz00OpPRIWq2UtpxaqOxOFCcPsIFJrPhzKQL2V
rRYsVUra3n2ICG4AZOcDxjF0riKikNUEAFoRvLcXqsMCd0IWBIOVbNB8kjVcENW3
oN6J9ZXx9ySqws4NRjYewoxYwPfrkUtiP3d7uGC6zhH7T/2nzyfwrNfqdnlIwwhb
soGGT+iC+Nyl3tZPTY1I6jEFd0655xef5Sw/08IydmBtGFH822ROhz2HOoYMJP6Z
G/i5/ksLnbnoM5J13m1efZWX2z1GSX43uqN6tJARbyqLFWdBSuoLYewZ+YBg/XOv
Fi7XAi9E35/dYrr7QEmjZcloAKKWdHoSHubba0+PeKaLrEKHxmVsOfPMTsFi44nT
KpOEgxgFN7lot/lnDLqso/jCv3Di1NRCmyfnwjHOOtaMZ76oStWEBs9F4PSBpKpv
o05l4eLAlOTbz7UpM1ks13nrLvg7PVSQsgcn1Z/z6c+SKMZM9tOCY8hK5GaDDTOu
fFPvyKH1UCyBUen3BppGKqz55OdQb+lcfdiaIBoYVpwvIVbXkIIOquKPw5lPhz4n
hYA8LC+Ko1MptVKz3tHT9QOy10r3+1Jjf+aZPreyNmKSow4Lx9kgZbENFu5sAVfi
78C07cFPJMQ72L3HcwUjQhLTGjZEgB4KWTHICjerk4qojQ1wPEgqh1E5T1ss9jOh
Rq20oo11QO+H4NKMhjJKvRiCQglmDkTVKg83HWWAtPRX3t2A38tRMfpNEGHvW9kG
PlxqAmcAGv4quc+xQbOGVjLHy0KJsSodBafqqCZARIgE1Og4bgmdETwU+MXAxLOp
IHBsH0be7Wq5zE2AfXH114YESnsvLFUoxxOrp2cL7atpTbCHVdyErSH418PKniC7
SuWKn3Xz1SsS4I5YaUTbs/8JIXpHqBLaViBvjoia91skt/+4pu3mAg0ZqbSj0yrw
5KGoJ0grXrmN7cRFLYO6c7uYkIZM/A7n4W9yhNxvl0oaTNOPVvp5rkbiM1JNPbMO
9W40OV6Y3kw5HhAsicC8cqLGHAXpjkGJkUnNwFAwpSeE8qzZYt3YepSgS0jicqXU
kp9Ctsym/Fs7OmTw0CgByyu1qg/vhCnYEvrjAF8231Zn4Vw1NKRb/Znh+vqEGyrl
737NrN618oKRr00di1FrAq4NoLkglHF+YTwIA0O/oCkUdyGuQ3YHngpLHP8SZAoy
Nep+wu4E5801f3sl1e8rb5toEuihhVW12SBEHPxfarD+7j0MeXx2s9In7t4ShycA
5rFfyLvqBoAzvtO8V1RalTEy16vqIgeRUqgsbc3z4rBdY3RHxquLGUHyx2UtZui+
Y7fsGkrkoSBPR7K/iKbG95HjxZfHSRtL52f57nBqv0KmwgcvXnQLAL6hmflxUsP0
UJ5AJgxuyA4lUQq2Mj11AoQpovqvgaSEAOQ5zZ1gFC2/WZb+W6X0KCjLls76pOYH
U23cv9blu4ln3/yo2LKv1uHFWUTXxsONcqbEW7Rd4jsIsL/CWApy72P2cJFMAlcB
Ji1kSYU3yAGYJNVZvjRjkFdja+iMP0++fDFtNjoU7epS6vOJiZ3F7RDC0l+7llzO
rGoL7y6yck6yJDBk4bdAfvPqU3ah466oOVoQfxjg+8kb8XqicmF2dlZfeSGnx0O/
oiv/h5tWqEDlmUsMMwpa3yiOrKACLPBlO6X9nCMii4zycIV7e22P2A+XQz02fuHp
4s4R3As+iQM+bvs51txhgtGpPfHR4md8l4gt9BVAuTPkp+M/ixwsKvF2DWri1+n0
SLfUBEGhspkiWvhr8VwVo5/9A/u/UYCUeGkQZJ/utRZxr+v9T3apVQf7srI/eVew
bjR82W0EYlFOY7rpfPoyT2cft2dWDD8rayqqwN+WxT9DPBnznTqMekI80jp0Xp9h
7B8ZbF8Cg20mDEQqgU+G3UCkjXON2i3OEhJ3pFVovIZ3j1Y45fbli98XpLdTPcRV
A2dYTGgvDscd99+Iom0ISUZa/maraEubl1L1QSVRm8qoY4W+X1gXYkX4+qKlesVA
lCwTl2a0wybysrAZoppSWrReD8PYn/MGAgTru5IxcoAR9sa+IyIoPlt/I9vB/kAk
EXMddZyX5OGvvnuP8NrxXEIJL/aEfVeZeXiL1o+0o1EJD5rjgSyYGhtg/PtGN+gx
8WF0YAfCmPe/XAXYwIOjVb/wf0Nbf37MmgrgqqK7ndHBdQrybecvDwi+45Ta0+pz
fCvLNKJZTrSC00kVRi6+PMswY+KxCurfLxdLD47m98YEO6s8gk7TqPXqq7GMYLq0
tSpPkUJiGkE9GCI8lotc9Lbz0vLmgLEEBDIPAQxMig4niu2DHLkSegnuAah5q3l3
mVcrrHb3TjNGzd+h1AU91sWoPotcTkIQ2tWSXalZwHH4ROkNPGFy4q6nLf0zZQ6W
N38uPUrPxD6ugkOU+cuUW25QqW6Sb76NuuPyIN14DQQUpUgAk+J1xGii0EQkaodH
KiK34V7vEZxa6AljQQ2YsTjSF5RMiGvGCc+han3vNaJmsuxH871GVklUCmx9njAA
WPtrPoWSrzOIT/ahURirdOWCqBsxHdH9nWdp6fnsWUqqCjscpG5LubDuzuctPS0S
0bsi0HDCuJHOBHiClD4fKOcbGuAzbljpP+RM8k583kh/mgGd0lvKyVa95KDeIjih
WzC4ep7/xAxV+dxZ+Bu2GdGbNfViQhZQDMSA1iSTfgNI1I7+OMjEl71cZV4LJJZv
H4zrfxeMR1eCUKFdZwb5rDpKblwYGf5PQZ+/O1nd4TN3JhEkBlvBHl79MTVIyqcS
VF0sl8/8jR+KMtTJjOtZA0CW4YL43hpyOvxEseTcSA5h/MuWCHoVcS/RYaa8dPcL
TI4HUxQaPIJAJ4DSCAFWd4sZthwha86hnZJVeakeDc5avXh5ERvppek6/eEB1o9H
0kHd4y0cwZqk3K19vKfidZM8QXJbSEoutiMyaZsMJM6XpWPH4C6BxIIbI3oG1G7h
QpfvJlXflNwo9/YySlvm6Yg9hNyJix6m0w6nhYCt7jLYtunlNnO2cO5wrDmy+A9+
p7NC6j/8bKxzIoxzb3L3szC/NEDYhhGhZPyKcsXZABlwuraOePb5/D2gF1W7X97H
bu13GBp05Ja1YQpZ2JaMab246NgvY9vcpWohLR2ZMI1F2MYQYguLKvCyY3fhG3U3
sPD/eb+AqGZihvVJpCI2v70JT6v7Olz1eaepV87YaMiDlSv9WPYavGKoQcLgjq27
2N7wVvxw3x3ChMYqxhrBzpLf3W1ApxnxO3fC3axdcN9/6GIOmGMPkb7kKwCfphLH
pRU4J6rqPGn8cRaqlvJ4Xxs/mvCodYBLX1ZNrKEdyV9WxPIf8sbTRYYAaxYa/0jT
unGPhjLxLQwGJENZF3fVO5UuTJDNxieAZjxZiWxcu/ExJM+7SAU25iAL7qhCwE4k
x8Mr3WZB91j/Dd/HPV/B7TohIdTJtF8YoUJ7lgSRGkouyhUf6EDRbtmaK3jjS3pG
fEvTFrmlBFvlbjILMTPRf5S6aOMTDU72HfkBn7EivGx0admXUt/P5+R/hoM9s8EN
zOUA1duSBvgxZwsODSQdNMXuSdu1UoBF3Yqkbz8fv4J3hz856oCkXzm2cAqukhX8
41VerBbXoO7jgbEtFPCBmNs2D+uEx1hO8OoIVAI8uzQcg80llQwa0P6CEe2/l0p4
G8z59DVocD0IxsYKRwZGD/kJZgOX0IvT7TDk48zfh3HpIDFyiNYys3n3J44In0T5
5xLoPrhBlSq9EhLA2rIuLzZXAKSMijRRiMWDb1g9Q7lkuHagM8hYVL7k8qaehQhg
kflnn2hkmtNEOb08Rh4OStIw4QLYCsDuYL0geR8jqBMqxfDZRGcqWLAwYZdULUzP
H8V0au2+FtBtr6jRFWFCNoANXoIKgxkHqt5DM3GkxATENzntA0h4gGKjttQ38scG
NxbFqOsC/eknzFpnmlMjdyIDlTzzf00c6/pBGOkTdnmeNPXQnwH7weZmk6xUxuej
49Cb8e3nPdt69stTpwgmX7cHX/UqvaI+eZQyFoSauYIPMNfLnIR0aJoKiXu003XZ
xx9f2Qhw64ozREf6bjqqqqjADIb5W4OsxBdbMTzF0ldXnUnQ7galFxRCg04RuR/o
OSNUJ7ezw+dzuvbmrGjmuPw1KIxUrw4HBdsKAb9en/DSleG9jEa6+oeGGNKbo1cI
JOF4zMLgwicmxr8rfUZDafeeOiKEfGfIfgIFNcYnE+DyDQiDiby+aZGqit9Fvwn9
1sjCdqWma+8BUJ7tWgbWPjDXtSM0CfQdubUK13uE0NpE9UQtd26CSz0cu7xXasq4
avwujJr6vfluf536Xn8qA7QIoxm4f93fhmm5MvUukSQ+QFAgl7xLlEF6v8XsMGFP
hDfStAj4Z5vKwvOFm//V7XEP5vYa64Mkitk6yCI5Cieee7v3txtzBTumrzISe6gK
WsWqyGa1SaLbOC2bOmusbwaAPbLO3JWWGDeA0Rn0ffPMNkqtm0J9prtDyJJmYEgv
VOg7nC96NsaaO7oCJ952yVDqOqwBABqXn6Limtwsnf+by4RXY9efLygnZsDOXIk4
P20KaLrl2IaQoR6F7pbSFszYXttwZIwx8E44RPs1bl2WDPYwQrwrdE6a9kAcIKCc
/QLtfCkKp9xKyUAp3yWXJlWI7nwoDhQeop9Q/2o5XyHceZrcjka4hYFThbriUF8a
XMvDUkWG1gixpgwawEtsZX65zgdZ7/uYPTboXXdW3/XjkaHMZZCgrrCdt6Jt3ViX
W/7N/V6/3RaZUlHZNHuDUpGPaGAG+yfRE+OX/DwD9oJSisEDUTX5s/IYgXMM3i7D
xuYGAiWG4U/YiIYX6nfMXVMPS7Rf8g4jl06H0/P+2TUqN8o6n6M+dCWHn4uhd/dj
IF0THQAyc93ZqkixhSi0NwuaJowCOsgU+DNgJURNrDQJLw8dC22Z93ESHtuDq1SK
sN9tj6GdtKacM2RG9SGXbvc/VPM7WTQmFlHyqjDJ2oyFqls3daMoqaPOioAYWXK8
pkQD09Xj0MNOh3cspS2e9JvKy+taIYXXjvr2JC/72+5jQ2o+zG5NaczWwG6/bMwE
JUtAIoRZD7aFNXstU/Qu03/lZdsuRvwi9RsrWcNzjKB8CSQpw99i3ecrCNzM6y6T
hgFHc8Z/AIEdE8mFB9n1uQRwVf8fLLJZrz4uYhuiYMIo8zLaTomECFwaSketi6FT
RdRYf/1F7V0+4een/1/vXBfWQRPskD1joIevEuPaiG+3rSAku7cgkNczmXw6JJE6
MYYSj9iiZ0uz1EDFaszshg==
>>>>>>> main
`protect end_protected