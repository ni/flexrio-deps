`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
JVp6A46tRdjg/Tc2e7jmDNv05OKzjRlw3XTH09qUJ7NV+HotD/UihAeyzbnezroP
euB1j3xbXzr8ckGaEw9iDdA6jjZQN4VbS33jydVZHQo22+mWms7Bf2wxQgHsftUP
AhG/xvLdg5LVax7xsXXZtnrj85N24MewGXzInLhtb7pL3oFitaQ7/xZWoQzMb+6k
Z3tIdF5ITE7UG1YP/qoUv7kZxqojx3qDxfyjwW+LUKzoEX3KOAUM71ymOez3WWdW
oql/it/qO4h6VpKxBJCrBh/CCwn9HbFRKCX8or4BsG1wpk7JxvQzn3F7VWZ1rLGy
vOvCJpanmMGd/IYfv3k9g08AuMQ3VfKMc8PuLdf+2fByFk6KWj92Eu4Udj8cicSW
m2GpjXn1M4btMt/7yOny4OgmOGw/4CcfEpPEwY0oJikDlh0JRhJ3l7MwQvq2eAIH
V9ayQaO1msYbaexiG57T9+bvYwVt/iM5VSXRNUgifGR9+Z60SyczcGwWu3IvhqWP
D2HAimz6TnYXbHctKFOPGDLCZezLAomD3ZyhW9oCG6jGSSxLRFDK0tcv08JBAYKq
ll/hx+zROoxBMR4gK/wUmKHB29MEkItTQRC8Rzayzvbios7cofrT5XkGDY9eyNmr
7ULfjitW0gdQ59+sGF88IVyXXFoLjRNxAjAzh0GYNFYjWOBVHHl+JN7gaHbqqwun
w1LYUgqcDFeMwqbLZlmXZV3SNmwHIRKX019O75XY/oPbqjc3uPBHjpiDrozRZGBs
PkPTdC8lHarZy0/N7h+meEgfJZ6TTQNNRWIVR2UIAq5xvum+YTN9D4e70kuMll3M
u7bCe+QEKOQ2WEZqzLQTHEXMml6XnFITsFsC9LFrITWg+eQyWa2Z22o6KBEaVKzr
v1jt8WaHsjFMyjkirXJfGzBgKG20dOX1JlF2zCWt3PUmpTI/PQrtwwtkmbyhZxJF
vfOZQ91vBfZO7O9Dt9NYjc5lMvYxISNbw6f78KoBxsZ7TLCR3ANfnLTghbKv9ZSL
G/0Xy30fcx2pClCtCcmQZPbBPIpI/rbvk6tPqgespneY2ODr/RxyBzoidsXIuAYc
0ski84vsoI+kV//I28gnmdHyKcEMhPWv6uImYcwFui2WoLllYekDSnPsG+zn1QG6
x0EURr+b2bhyPmMRgIEINJ7gz2US7yIBZ8YPsJhvzvte1QqpoBttSQGOvoBsBTV2
I4tgQj1FrUjOsnFc2xy3PQudN4HDg1yhweOBk3xzkIXkX21px6G+c/7o+JNS5lUR
dy30eBxaLR7JmYrHwfVFpBCSkMPqHKHZelqhLw3WrNs2Jv8G1mp4xTvXibV/IkHT
Syq/MouamzOzEooNeAewrif4XZxE4+6doYgCKfJ6NonFQRIgZv74OYkUbugoiABL
Qu5HzdRX0RiG9YPxI8Mf+WAHWcbKHDzhpgCZUURcxcqe2Os7Q/G7Qv681LwRBOkm
kuvWajiqxcUt0fx9oaDe+egmreDgSy1WKlNOgkEWu8JmtZ8WH1Yn+KajhbHubENy
sKnC1hGi+nxaDbGxcZPhByiY6vcrx+8RAcyVyIL3OxonlRLIkYfGZgFwZrL/2yKZ
zcefNuBjpMyDfzUck7yHf+KsMGme6GDdJCEivb486QsPYXRK+36NLf1hgCxpGiDr
O9YCOJ8ryEkFkGi/w8u/LezZ9NVOoYT+zOBA6Ze/ZV2JNnPmo8Hhn9QVPkVXdtV2
spV+FNF1ngUPPYsHpzLnmnqpqyEgMdIChlNuvxQW/JeQ91Ga4IwrRPy2ZFbnxYOL
tj2WoP6HnqMgrkz+sV1Cm3yCJTbMW04NFEWV6FTRr7n0i/mzKXhTNS41f+SeYPif
xFEWV62eY9rmXlnUhrPxPT0jtXP9NlDTenwCZFMepgiuwVTLnkTRQ6RvlEl0YUmm
QBATlWzrLCen6pGsNwF3DKGKJcuJKjbPz8xZmdzciXjbC1lhGQx/ksiaZ0snTgjP
IO53c2fa46T7meca2koYrXi1m+deqBLeojgd96NtzPJethEKINiDKc0mLmP83KFB
VccJXw3+iKvN0E1cgsi13XLAYs4sm6Z8fnNgSKS/4AECmZnQIbEkmziTKd1bp2Rr
GA0mzVh1inpFQA5Ee3A4UAwteHwC66mfw/DyY6IkAtTDr2EenppRPuRbOIo6uQ81
ZrWK7Zodpq7vJmQKPEQPW3V5F83pqS1a7cRbMnVA3N6b3sSqHAMCeS+r1v86JjPw
SEIloNSqNZaYtc2z4lbEi4exAcMJDrb/fE7WzcUxBsUBijo8FML4QZA1LAiRf66r
6326jTYi/E+KgP/X7XGiyZPBpn5IaoWeIKX1EO8Ruo+sBPk88slaooraUd3++kk+
MsZSuOxghlUSiy6wOwmdpxRA0YiSAtB+HbBrJrhIBYFfjnJSajal/BXdWAXueI3P
lWJfZxETxY9zLFsgw76XBmccfOF+aCcPzSqpGyRmz8SsNOkAIQBxDgDmXOnNJ7UQ
Gm/qz7LOgrD2VXccPD3IF1/sVQTnT9hzW0MtW6dr/T4xvOe8wiW1v+WXfhOo0mmz
s1hHZaFvHzN+AvADlZm8SXumam+3HbkruTJWtYgYMvKo0uH0RiZRra3Oq+39orfC
c+Zm7HLGooCrCKwp/ftkQkeQ9YVDpMJ2KaeFHRRU0h3WI1RshQ9XTB5vCqRFIRme
IrPHA1c0k9dzdQICLWOH3K16/yf9BFZlkuZ4CpUvDXKDUH6w4Q/j8lYEqrxF1Cfo
clmSRnSUSLEFrlN8G1oKOzR9LPfo8VSsVgfNyWhM9X8b2/6RGckHXZv/upPY/b1/
lccs7vOHdJpYKTeM+ZpbKPnl6CruRoUdmPuyH7J6wJhM2QykMZ7LGwdmJ4cYXfME
SuWkvI6sgYe7Yo0MlbAt0iGrHw1gIiR77+5klySbP9xVxDumuxsUxBCWye4skbmP
XdIRSvSpuDuPW4O4vVue6Xaou6cosYGr/CotYIJVH1TLDUro+prD5HThMfaGnfUB
DHRZn/NFV2IJ+5DB2MI+NEEwPjYSGp/MH+XSyw+sCqKaE7R3ieCMk9Ur2DWuKLmH
VrkMrwbMQ2YNNQSt5kbjmFxn4eoIPnHdtfsL9L3ncGdjrez3PA5zXpjVfSD3Wizu
GYFahFU8FzdqY0UFTI9NdoiI+eim+2mduKzc7TVzdWzAdpMipUxdqeazSR5o1u/Z
eb10pHDeEz3XLzrlPuAAsIReHFZN7aJMPWeWUachDl+pTkD/yH6OmsuXJlf5TFjz
DxpwaGP/YVEIic8QldgjkCRaaq0W2H5g2mX3bHYfNVbIOYk+GGTAwa/xMUll/2Gv
6BgKAXtCeJfupz1sBV4vrLfZ2GotNbTs1X4CdDLDHCJholYvKcTAt03sALPQKcg8
l5CMNQ3VQZ8CRDHSkGZfTNxJExs75+YJ9BVS4UO6dtlnd+CYfCeBNcozRtWP6ZD/
`protect end_protected