`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCxJP2IrjSeGTG1/XKiQfrCRWpLtKouCgr61lojmUIZJ
m/jKacvkQnOifMy5zgBBYS1y2XKa1TGJ6JuHJ+RS098+l8Q05h8B6bQqN1PLkTJp
1bpvtmYvm9ds2sHHd2pMmiZ04kkiJZISeBo8ITlOk2Trgvxgs7xPBcNFmV9zC07u
xTv+Q8xSECrFnFGoHi/oBTlJ3Z4NDbbAasxC4ZSFXItcGI+NEBh644mQFSQR8whP
5u2UGQRwQtSPO2eZUdrgaFdJJpxB4oi+hPDZE8w+/tW7TmP2b4cbBVhUgDEkpALn
jZXSOJ8lEqPPHIIvbEGLVGfjDg1qpcSzbA4L3bURTqrr0a16ysDkYTACmYMXXEhX
g9qIf+MYrGzMhx43/ZCrxC3BJ+L1cALezzx6u7sfZMP6B0f2CDzqtFScZ/HlazK9
lU9bOG+vNB0e6phxiq3ihhFaJKsA8i2FSw8GJEh1+Y/tXsZRq9rOByXt/+GN8Q4Y
nptfQmQkYqwyXQx05WG/5vWuP032SRVYgROaCJwfUiYvslI5s63cDuUGIzQgVPCb
5xDOC8EJNSqsgyDBEY1Ex5JMeDpYbV24I9nGydKaipXRqjnf4rgmMZHRyAZMVjt/
BVPJFzPNHtntkqf2unc1mrTKfsg3DjQy7ln0MJniomawOgqHjj4atnm9rq6Lo7bZ
FKEcuIyhvxZbG+66LSITfrljpu5VeU71eXRqD1A++nj5CZzmFokFJkJYvY6l5ntw
CBEc9mkRCNkSerutz+3IkuTWkzgDwykgJgVVqJ7u4uNCSUtPpREXHYZjIRQKT60t
UiYwCVf67KcczP+OfCUbdVrfq2MWdT+BzKXq9wZRNpv8pAkKWcdZ0SpNKGnflZMs
QbM1VjyL0KPc8EC/QavLUXJlYq3Z5LnTMY1QUL2IMsc+bXLmChPD+z+EXJa4o26G
jDAszGPfq3sdoK2VNJGQLKKPDnQp+MNqMuckYz1xTvUk0BevZxMNY/kIAybaETLr
gIoctve+rrM0cB6HSteNTNloGQ4Ilf5FjlF5yesOKRQWovHRhT0+uYhUSwiUgftw
KsUcBh1bLLPk58AAqloNNtN8CYAi8hlFK/fCL3ZZtUd//3sFl1Lrf7kk9gQtYgQu
C+Wp+vUY3P+tFYJ+hGggsxPjCzkn10h2s2Nz+80nt/kJ787JXokzG5kNQfOVmfTl
kTY5kamKTqIlK0tA1sKyEabRBfLLBkf/vcdANrzS6MuNkJ6BKyDMvICbKAfuOvIS
r3PvaEkSXimYoHx9mPJB1u5bybzBItWqBTBPyHDqkvDmCcepZznGQWgV1S6htqNL
YfrbIVNGKHq5EFl9mncdSjSL6OejZ4fBnQ5MKNKTd4fmvXM8aINrmXEn32AAPUdM
scwUJPnt5iXKkCNa+AswSmGP9JGQBjkuU6fFr6xzmV9iWi3qzuG44bFVT/ECzArk
mr2xppdsPuraNKTn59LWjb8sTym2Tu6vzsCGkLSWGZW4Hdd9xstxpyDMgk9Sf2R6
wTFbJBreMq2tqHKiiFuFqWroMKnYCp0O1LPBGtj7+yWEgr7qp3XxKyuth2uK2U9r
Lrg0hojwAXrNbPLSb4UUa3JPE744FVuMqCECiNbue+4R2rbMNAS2OA4HqJZ63n0i
EyJzgM1bdPXkRMQJ3ECiEHAVsvtdUoxzLcmRwIA/S9bPnelDGKrwATvp0f+8SX1X
6iOcqbKgiYRMRNX44LQ6bBb47nqZlqk8yQlW0IlUWgNjKdEpMT5D1FA3VxmKrOUa
eJkUSIMvb9HJOhu7ZgE519/h5ROWq8jD5KwHkxZkNqSWmFktuP0zY6D9MoOtKRb9
FHm7grQy6spuy6Ggc37qwmqnsbpXKb1RRk4IfhKNRPTou0Jrb7zyrWYdSSzEZIHB
xlELv7pRuz8nzrmB3o8zxoKeXf2J0XKit1OEtxBnRAzyP99f2hm1nFNJI0DXnigr
0lLYu+oAEBx9EFTqv2ZZ8DVfCv0Te7Pj3A4Log5BUUQPYAEJimXkyxsClNdNd6v8
IKWQCpWfK+2lcZiKpBI6cq8Yp8rxFi+V6cjyuNBCfjb+LAxf1/j1gvoHRY/Hzydv
di59KKkdnA2NVhy0TJRz/1CwsNnzRGZx+SENdAjUIvCx/xI4NAMgzBqyIa+jKoT9
iek9FgrvRbxyhuHMpTK2G9fKjVOc9M5gmAi1YnmXiJHldHfTKiopNvlkf+bsdzmW
iVXx+9oCtFWz8qPzLb11r24w3j863Q721k+8prwkJJd5jmdqpYeJzmJQ5jWKM1YD
mYoIjzs3YkLH9j46Wq4nJFLeUfFl42qOf4KOhk/A3RchfEvyyw9UOZo26X3GFdby
gtPyIhTtj/fmo7mDReqaYnRyj/tgXMm1m5uNPAQn1lVtyz4y/OFW43aEJz9mkHZw
JDsz/xVpSKjy6qrqfejngAReAmNrD/w39VnPjr0wXlOo3yenJaHH9fmlqdDpn7/v
N2k1phMH6A4hQm1C+pxbKWhU3PqsNAiccJzY4VGr3hDxXXDrR1svspD9Uk7ZHti+
HJNiVJapcE9g9TPqhzZdq8eL1C3qaXJwiy8hTv3OZfhUqVyxzrNc1crElUMFV6dy
u+kFdgu2Mq9GJIpq4ieBD/AgLjAZraUWziSpHGzAvUFdUKA0t6hRrTvwzxNc4/bo
AqVfuU8fENenbTBTlxER+QEgYEmS4p6V2VOLJrSEgpzAXF9m9Ah6u0KX6DVBZ81Q
IlusNe4dhKmmVUGw7upVb59ps19PRJOP5nsq4kCQzUy+gnq3ui8Caxe0/mXuXfdj
WI8eAMYErM96L4ihhT7J4FYXE+J84xtRHEeg8O8Osu4leUp7aqg/gfu7DNAC/VE0
N4tIljZcGpxhV2DVPzmb/J3WjukzPZga5Yz6HA1lSsf7jdRNKnEMCj7EmFu1WI19
FghZuUVNXXt+4VzhIa4pAtKfwJEH4ZXTpoQjsnNgnna6Wg3ZimhWk8+KjmFHYcP4
wbYSTQqFRqRgFIIkWQVVVjXQmU9VqzLXTH9EUwTaYu/5iq8N2MdH+2DLWFaMah89
DACOWDecbjVhlc3yNbHVX83mamIIGIARJOnM1Oz1axA/szfFFTRWUyibkrUojhB2
t4sKrdQELuOBlcrXakPlt7a3VtymchZi+id3OnURXVTKE/EWBpedEf8rEVQs1Bqx
1N5ShtrKXcgIUBl8JVd6NQrIdWBBbG1LvWO+J858dX6Tv4UAWJo5ZCbysKcuVqlN
0YItphdB9tydY3ezYCN5GqyJNwquxyblNjiLH06wDWeZTCGZnvCBlqXyVxTQgntF
fEBSHEXAlazksXEGxRJ6OUPj2fTgWlOuMP8Vdsjz4maumL9KXcd2c6binD9/9+iu
9U6inS3nXkMjdrDQAsAzO7BpyLLa1g2YAygNlIoCeAQoKd3wGvxEhJ84Tt20bbmM
YPWAMAQ+4dvj0pZq3byLohemrMsJH4IVkMQadz3n5APQfYKZIKHB9pXb7xevVCkA
J4b/j4j+F/0YYAkRcqQfJeLsdQKFR7BeGOW6wy5DK5FDTdmkhlGq8e3ElMt5Z+lf
HG81kmNzOsRbulRAtl/PRwsi4oKMLo+rfRukJ7EEARiKrL8jV12toKbZ3V05yY6Q
LjZhjYnRkhbLRSMXnIU7hP2cOccS4EUzRUb9VqvHqJLPAR0GfNnzuDNlmUWO1oib
6xFDFkLpi+STCchtbxYxoKTPwyT8gIT8BxpgMih27N+i2IlKTzC2dHK5zPjBb+Ea
nhQJ66TrpxtzHkuZy9Y+pjGw8o1P6SxBk8IRxRAdUeefaTr/nnoQ8wXa8BIoAMA/
bIQ46tzalfy2ugkHcn8z2IIxu9AtCbYeiQLamXKlXtLSxSLXM9UIYjzhcnK6G5DQ
VEuLEHrMZFA6g7Hibof58Jrqn95gnhwTUehJa4rgmTZcKzOXNDa2RO6W9XqXXpFF
s/qgzMBKaVmizSR2GEPsqgcJB7MxQN/8+geJwhk3JTgfctiHuMOEAMBtfsDZKuBu
p190vT/0COTKTpC2BE+Qxoc40zH+plYZRpfpY6Gq4JlBaupum6+17Fj3Gqb8ZZVU
S/ffFCMq7DvWKtUeOSuADmT0TJ+YnmtLLTKrzQZvCoTCgJxXbGbCWeFlK//mqsUF
isYcivpBObz1LFptD4BV8lt2+85Dx9SHUcYaldugcvPWENsu4MaLS6FXuhvQ/IOK
pH0fcdO80fvqZS5AFyJi9NgO6MzeNkPDEsclWOkXKrnREim+Y8s/Fyp+tuqcxBDC
5zmEcmoTyVG5cMehxr0dsmHeEtNjVk/TfoN/rJZSi50TVjQO92giZfdNfSm5K9kT
SH1wZlqIzo+0He1T/n8xa7Aw/ULDT4e9ryIwxqNPBCn1xgqRuepVUvt/3YliEL6C
xT4+h0KKrmfD7XN6aRnQEy3Lon7ElA97RKH7rQserNh8x0PbFZ69NXIwEPf4682G
u43CyPhqBNQ2X7iDSGVqLukA6uigSaC0Qhp0Exkjgp15+PG68EOVsOMJm1nVhXa3
RiMyqoRwQVtUJsygvXHpe0Y1dKbJ6FLSmLAel+NpIveccojO8ByvSX4wDsy4ug4+
GtdQivGCS3fNOJ8tPZsnpT2KEhoMP4IoONFIrozAUQ3FiAZLvirrQcFGWCuXSf3B
YZ114OwPVwaMZ8vkSHhsr8vj6eAKv4E4veJzLz4vUh3O7/BQezVXQ5+Mvia6r5fS
LQ3jEv61M++HmB5spdUAbVkQdMeGkMdBgABzlOq9UbqcvHRVOXxGtP/7xQhQ7+Mh
OCCQMcRv6nMFsuI2gl17DnxLkFSgzKyvWMWCD0gqTrTdwNYYYUyb41Lon0lyqwER
3gWZZ7/zKH3klgnuwvtI7VJnf9obIEZEHTgHeq0N+TUt0iVile9IW+8K6lNflzc3
Ctx0E2gazRkM0h89cWd4uMbUQAGz/gVWQC0HloEeT9svuxyiB8Z+CyoNxEIWhLlO
Xyg2rwk/R4kLzfEvJQ9IF/1dWXOQ9p+kn5ppxxJhIByYCSXyElYo5Hj0v4j1PMNc
m5kl68vd60KfreYT1MMxDHPZK/l08KHAH58UyGRHGt46xUahYfC2n2wPxGHRsgTK
0XRA/tu7dbKtR+3hgTlX/A==
`protect end_protected